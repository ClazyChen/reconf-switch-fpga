module Hash(
  input          clock,
  input  [7:0]   io_pipe_phv_in_data_0,
  input  [7:0]   io_pipe_phv_in_data_1,
  input  [7:0]   io_pipe_phv_in_data_2,
  input  [7:0]   io_pipe_phv_in_data_3,
  input  [7:0]   io_pipe_phv_in_data_4,
  input  [7:0]   io_pipe_phv_in_data_5,
  input  [7:0]   io_pipe_phv_in_data_6,
  input  [7:0]   io_pipe_phv_in_data_7,
  input  [7:0]   io_pipe_phv_in_data_8,
  input  [7:0]   io_pipe_phv_in_data_9,
  input  [7:0]   io_pipe_phv_in_data_10,
  input  [7:0]   io_pipe_phv_in_data_11,
  input  [7:0]   io_pipe_phv_in_data_12,
  input  [7:0]   io_pipe_phv_in_data_13,
  input  [7:0]   io_pipe_phv_in_data_14,
  input  [7:0]   io_pipe_phv_in_data_15,
  input  [7:0]   io_pipe_phv_in_data_16,
  input  [7:0]   io_pipe_phv_in_data_17,
  input  [7:0]   io_pipe_phv_in_data_18,
  input  [7:0]   io_pipe_phv_in_data_19,
  input  [7:0]   io_pipe_phv_in_data_20,
  input  [7:0]   io_pipe_phv_in_data_21,
  input  [7:0]   io_pipe_phv_in_data_22,
  input  [7:0]   io_pipe_phv_in_data_23,
  input  [7:0]   io_pipe_phv_in_data_24,
  input  [7:0]   io_pipe_phv_in_data_25,
  input  [7:0]   io_pipe_phv_in_data_26,
  input  [7:0]   io_pipe_phv_in_data_27,
  input  [7:0]   io_pipe_phv_in_data_28,
  input  [7:0]   io_pipe_phv_in_data_29,
  input  [7:0]   io_pipe_phv_in_data_30,
  input  [7:0]   io_pipe_phv_in_data_31,
  input  [7:0]   io_pipe_phv_in_data_32,
  input  [7:0]   io_pipe_phv_in_data_33,
  input  [7:0]   io_pipe_phv_in_data_34,
  input  [7:0]   io_pipe_phv_in_data_35,
  input  [7:0]   io_pipe_phv_in_data_36,
  input  [7:0]   io_pipe_phv_in_data_37,
  input  [7:0]   io_pipe_phv_in_data_38,
  input  [7:0]   io_pipe_phv_in_data_39,
  input  [7:0]   io_pipe_phv_in_data_40,
  input  [7:0]   io_pipe_phv_in_data_41,
  input  [7:0]   io_pipe_phv_in_data_42,
  input  [7:0]   io_pipe_phv_in_data_43,
  input  [7:0]   io_pipe_phv_in_data_44,
  input  [7:0]   io_pipe_phv_in_data_45,
  input  [7:0]   io_pipe_phv_in_data_46,
  input  [7:0]   io_pipe_phv_in_data_47,
  input  [7:0]   io_pipe_phv_in_data_48,
  input  [7:0]   io_pipe_phv_in_data_49,
  input  [7:0]   io_pipe_phv_in_data_50,
  input  [7:0]   io_pipe_phv_in_data_51,
  input  [7:0]   io_pipe_phv_in_data_52,
  input  [7:0]   io_pipe_phv_in_data_53,
  input  [7:0]   io_pipe_phv_in_data_54,
  input  [7:0]   io_pipe_phv_in_data_55,
  input  [7:0]   io_pipe_phv_in_data_56,
  input  [7:0]   io_pipe_phv_in_data_57,
  input  [7:0]   io_pipe_phv_in_data_58,
  input  [7:0]   io_pipe_phv_in_data_59,
  input  [7:0]   io_pipe_phv_in_data_60,
  input  [7:0]   io_pipe_phv_in_data_61,
  input  [7:0]   io_pipe_phv_in_data_62,
  input  [7:0]   io_pipe_phv_in_data_63,
  input  [7:0]   io_pipe_phv_in_data_64,
  input  [7:0]   io_pipe_phv_in_data_65,
  input  [7:0]   io_pipe_phv_in_data_66,
  input  [7:0]   io_pipe_phv_in_data_67,
  input  [7:0]   io_pipe_phv_in_data_68,
  input  [7:0]   io_pipe_phv_in_data_69,
  input  [7:0]   io_pipe_phv_in_data_70,
  input  [7:0]   io_pipe_phv_in_data_71,
  input  [7:0]   io_pipe_phv_in_data_72,
  input  [7:0]   io_pipe_phv_in_data_73,
  input  [7:0]   io_pipe_phv_in_data_74,
  input  [7:0]   io_pipe_phv_in_data_75,
  input  [7:0]   io_pipe_phv_in_data_76,
  input  [7:0]   io_pipe_phv_in_data_77,
  input  [7:0]   io_pipe_phv_in_data_78,
  input  [7:0]   io_pipe_phv_in_data_79,
  input  [7:0]   io_pipe_phv_in_data_80,
  input  [7:0]   io_pipe_phv_in_data_81,
  input  [7:0]   io_pipe_phv_in_data_82,
  input  [7:0]   io_pipe_phv_in_data_83,
  input  [7:0]   io_pipe_phv_in_data_84,
  input  [7:0]   io_pipe_phv_in_data_85,
  input  [7:0]   io_pipe_phv_in_data_86,
  input  [7:0]   io_pipe_phv_in_data_87,
  input  [7:0]   io_pipe_phv_in_data_88,
  input  [7:0]   io_pipe_phv_in_data_89,
  input  [7:0]   io_pipe_phv_in_data_90,
  input  [7:0]   io_pipe_phv_in_data_91,
  input  [7:0]   io_pipe_phv_in_data_92,
  input  [7:0]   io_pipe_phv_in_data_93,
  input  [7:0]   io_pipe_phv_in_data_94,
  input  [7:0]   io_pipe_phv_in_data_95,
  input  [7:0]   io_pipe_phv_in_data_96,
  input  [7:0]   io_pipe_phv_in_data_97,
  input  [7:0]   io_pipe_phv_in_data_98,
  input  [7:0]   io_pipe_phv_in_data_99,
  input  [7:0]   io_pipe_phv_in_data_100,
  input  [7:0]   io_pipe_phv_in_data_101,
  input  [7:0]   io_pipe_phv_in_data_102,
  input  [7:0]   io_pipe_phv_in_data_103,
  input  [7:0]   io_pipe_phv_in_data_104,
  input  [7:0]   io_pipe_phv_in_data_105,
  input  [7:0]   io_pipe_phv_in_data_106,
  input  [7:0]   io_pipe_phv_in_data_107,
  input  [7:0]   io_pipe_phv_in_data_108,
  input  [7:0]   io_pipe_phv_in_data_109,
  input  [7:0]   io_pipe_phv_in_data_110,
  input  [7:0]   io_pipe_phv_in_data_111,
  input  [7:0]   io_pipe_phv_in_data_112,
  input  [7:0]   io_pipe_phv_in_data_113,
  input  [7:0]   io_pipe_phv_in_data_114,
  input  [7:0]   io_pipe_phv_in_data_115,
  input  [7:0]   io_pipe_phv_in_data_116,
  input  [7:0]   io_pipe_phv_in_data_117,
  input  [7:0]   io_pipe_phv_in_data_118,
  input  [7:0]   io_pipe_phv_in_data_119,
  input  [7:0]   io_pipe_phv_in_data_120,
  input  [7:0]   io_pipe_phv_in_data_121,
  input  [7:0]   io_pipe_phv_in_data_122,
  input  [7:0]   io_pipe_phv_in_data_123,
  input  [7:0]   io_pipe_phv_in_data_124,
  input  [7:0]   io_pipe_phv_in_data_125,
  input  [7:0]   io_pipe_phv_in_data_126,
  input  [7:0]   io_pipe_phv_in_data_127,
  input  [7:0]   io_pipe_phv_in_data_128,
  input  [7:0]   io_pipe_phv_in_data_129,
  input  [7:0]   io_pipe_phv_in_data_130,
  input  [7:0]   io_pipe_phv_in_data_131,
  input  [7:0]   io_pipe_phv_in_data_132,
  input  [7:0]   io_pipe_phv_in_data_133,
  input  [7:0]   io_pipe_phv_in_data_134,
  input  [7:0]   io_pipe_phv_in_data_135,
  input  [7:0]   io_pipe_phv_in_data_136,
  input  [7:0]   io_pipe_phv_in_data_137,
  input  [7:0]   io_pipe_phv_in_data_138,
  input  [7:0]   io_pipe_phv_in_data_139,
  input  [7:0]   io_pipe_phv_in_data_140,
  input  [7:0]   io_pipe_phv_in_data_141,
  input  [7:0]   io_pipe_phv_in_data_142,
  input  [7:0]   io_pipe_phv_in_data_143,
  input  [7:0]   io_pipe_phv_in_data_144,
  input  [7:0]   io_pipe_phv_in_data_145,
  input  [7:0]   io_pipe_phv_in_data_146,
  input  [7:0]   io_pipe_phv_in_data_147,
  input  [7:0]   io_pipe_phv_in_data_148,
  input  [7:0]   io_pipe_phv_in_data_149,
  input  [7:0]   io_pipe_phv_in_data_150,
  input  [7:0]   io_pipe_phv_in_data_151,
  input  [7:0]   io_pipe_phv_in_data_152,
  input  [7:0]   io_pipe_phv_in_data_153,
  input  [7:0]   io_pipe_phv_in_data_154,
  input  [7:0]   io_pipe_phv_in_data_155,
  input  [7:0]   io_pipe_phv_in_data_156,
  input  [7:0]   io_pipe_phv_in_data_157,
  input  [7:0]   io_pipe_phv_in_data_158,
  input  [7:0]   io_pipe_phv_in_data_159,
  input  [7:0]   io_pipe_phv_in_data_160,
  input  [7:0]   io_pipe_phv_in_data_161,
  input  [7:0]   io_pipe_phv_in_data_162,
  input  [7:0]   io_pipe_phv_in_data_163,
  input  [7:0]   io_pipe_phv_in_data_164,
  input  [7:0]   io_pipe_phv_in_data_165,
  input  [7:0]   io_pipe_phv_in_data_166,
  input  [7:0]   io_pipe_phv_in_data_167,
  input  [7:0]   io_pipe_phv_in_data_168,
  input  [7:0]   io_pipe_phv_in_data_169,
  input  [7:0]   io_pipe_phv_in_data_170,
  input  [7:0]   io_pipe_phv_in_data_171,
  input  [7:0]   io_pipe_phv_in_data_172,
  input  [7:0]   io_pipe_phv_in_data_173,
  input  [7:0]   io_pipe_phv_in_data_174,
  input  [7:0]   io_pipe_phv_in_data_175,
  input  [7:0]   io_pipe_phv_in_data_176,
  input  [7:0]   io_pipe_phv_in_data_177,
  input  [7:0]   io_pipe_phv_in_data_178,
  input  [7:0]   io_pipe_phv_in_data_179,
  input  [7:0]   io_pipe_phv_in_data_180,
  input  [7:0]   io_pipe_phv_in_data_181,
  input  [7:0]   io_pipe_phv_in_data_182,
  input  [7:0]   io_pipe_phv_in_data_183,
  input  [7:0]   io_pipe_phv_in_data_184,
  input  [7:0]   io_pipe_phv_in_data_185,
  input  [7:0]   io_pipe_phv_in_data_186,
  input  [7:0]   io_pipe_phv_in_data_187,
  input  [7:0]   io_pipe_phv_in_data_188,
  input  [7:0]   io_pipe_phv_in_data_189,
  input  [7:0]   io_pipe_phv_in_data_190,
  input  [7:0]   io_pipe_phv_in_data_191,
  input  [7:0]   io_pipe_phv_in_data_192,
  input  [7:0]   io_pipe_phv_in_data_193,
  input  [7:0]   io_pipe_phv_in_data_194,
  input  [7:0]   io_pipe_phv_in_data_195,
  input  [7:0]   io_pipe_phv_in_data_196,
  input  [7:0]   io_pipe_phv_in_data_197,
  input  [7:0]   io_pipe_phv_in_data_198,
  input  [7:0]   io_pipe_phv_in_data_199,
  input  [7:0]   io_pipe_phv_in_data_200,
  input  [7:0]   io_pipe_phv_in_data_201,
  input  [7:0]   io_pipe_phv_in_data_202,
  input  [7:0]   io_pipe_phv_in_data_203,
  input  [7:0]   io_pipe_phv_in_data_204,
  input  [7:0]   io_pipe_phv_in_data_205,
  input  [7:0]   io_pipe_phv_in_data_206,
  input  [7:0]   io_pipe_phv_in_data_207,
  input  [7:0]   io_pipe_phv_in_data_208,
  input  [7:0]   io_pipe_phv_in_data_209,
  input  [7:0]   io_pipe_phv_in_data_210,
  input  [7:0]   io_pipe_phv_in_data_211,
  input  [7:0]   io_pipe_phv_in_data_212,
  input  [7:0]   io_pipe_phv_in_data_213,
  input  [7:0]   io_pipe_phv_in_data_214,
  input  [7:0]   io_pipe_phv_in_data_215,
  input  [7:0]   io_pipe_phv_in_data_216,
  input  [7:0]   io_pipe_phv_in_data_217,
  input  [7:0]   io_pipe_phv_in_data_218,
  input  [7:0]   io_pipe_phv_in_data_219,
  input  [7:0]   io_pipe_phv_in_data_220,
  input  [7:0]   io_pipe_phv_in_data_221,
  input  [7:0]   io_pipe_phv_in_data_222,
  input  [7:0]   io_pipe_phv_in_data_223,
  input  [7:0]   io_pipe_phv_in_data_224,
  input  [7:0]   io_pipe_phv_in_data_225,
  input  [7:0]   io_pipe_phv_in_data_226,
  input  [7:0]   io_pipe_phv_in_data_227,
  input  [7:0]   io_pipe_phv_in_data_228,
  input  [7:0]   io_pipe_phv_in_data_229,
  input  [7:0]   io_pipe_phv_in_data_230,
  input  [7:0]   io_pipe_phv_in_data_231,
  input  [7:0]   io_pipe_phv_in_data_232,
  input  [7:0]   io_pipe_phv_in_data_233,
  input  [7:0]   io_pipe_phv_in_data_234,
  input  [7:0]   io_pipe_phv_in_data_235,
  input  [7:0]   io_pipe_phv_in_data_236,
  input  [7:0]   io_pipe_phv_in_data_237,
  input  [7:0]   io_pipe_phv_in_data_238,
  input  [7:0]   io_pipe_phv_in_data_239,
  input  [7:0]   io_pipe_phv_in_data_240,
  input  [7:0]   io_pipe_phv_in_data_241,
  input  [7:0]   io_pipe_phv_in_data_242,
  input  [7:0]   io_pipe_phv_in_data_243,
  input  [7:0]   io_pipe_phv_in_data_244,
  input  [7:0]   io_pipe_phv_in_data_245,
  input  [7:0]   io_pipe_phv_in_data_246,
  input  [7:0]   io_pipe_phv_in_data_247,
  input  [7:0]   io_pipe_phv_in_data_248,
  input  [7:0]   io_pipe_phv_in_data_249,
  input  [7:0]   io_pipe_phv_in_data_250,
  input  [7:0]   io_pipe_phv_in_data_251,
  input  [7:0]   io_pipe_phv_in_data_252,
  input  [7:0]   io_pipe_phv_in_data_253,
  input  [7:0]   io_pipe_phv_in_data_254,
  input  [7:0]   io_pipe_phv_in_data_255,
  input  [15:0]  io_pipe_phv_in_header_0,
  input  [15:0]  io_pipe_phv_in_header_1,
  input  [15:0]  io_pipe_phv_in_header_2,
  input  [15:0]  io_pipe_phv_in_header_3,
  input  [15:0]  io_pipe_phv_in_header_4,
  input  [15:0]  io_pipe_phv_in_header_5,
  input  [15:0]  io_pipe_phv_in_header_6,
  input  [15:0]  io_pipe_phv_in_header_7,
  input  [15:0]  io_pipe_phv_in_header_8,
  input  [15:0]  io_pipe_phv_in_header_9,
  input  [15:0]  io_pipe_phv_in_header_10,
  input  [15:0]  io_pipe_phv_in_header_11,
  input  [15:0]  io_pipe_phv_in_header_12,
  input  [15:0]  io_pipe_phv_in_header_13,
  input  [15:0]  io_pipe_phv_in_header_14,
  input  [15:0]  io_pipe_phv_in_header_15,
  input  [7:0]   io_pipe_phv_in_parse_current_state,
  input  [7:0]   io_pipe_phv_in_parse_current_offset,
  input  [15:0]  io_pipe_phv_in_parse_transition_field,
  input  [3:0]   io_pipe_phv_in_next_processor_id,
  input          io_pipe_phv_in_next_config_id,
  input          io_pipe_phv_in_is_valid_processor,
  output [7:0]   io_pipe_phv_out_data_0,
  output [7:0]   io_pipe_phv_out_data_1,
  output [7:0]   io_pipe_phv_out_data_2,
  output [7:0]   io_pipe_phv_out_data_3,
  output [7:0]   io_pipe_phv_out_data_4,
  output [7:0]   io_pipe_phv_out_data_5,
  output [7:0]   io_pipe_phv_out_data_6,
  output [7:0]   io_pipe_phv_out_data_7,
  output [7:0]   io_pipe_phv_out_data_8,
  output [7:0]   io_pipe_phv_out_data_9,
  output [7:0]   io_pipe_phv_out_data_10,
  output [7:0]   io_pipe_phv_out_data_11,
  output [7:0]   io_pipe_phv_out_data_12,
  output [7:0]   io_pipe_phv_out_data_13,
  output [7:0]   io_pipe_phv_out_data_14,
  output [7:0]   io_pipe_phv_out_data_15,
  output [7:0]   io_pipe_phv_out_data_16,
  output [7:0]   io_pipe_phv_out_data_17,
  output [7:0]   io_pipe_phv_out_data_18,
  output [7:0]   io_pipe_phv_out_data_19,
  output [7:0]   io_pipe_phv_out_data_20,
  output [7:0]   io_pipe_phv_out_data_21,
  output [7:0]   io_pipe_phv_out_data_22,
  output [7:0]   io_pipe_phv_out_data_23,
  output [7:0]   io_pipe_phv_out_data_24,
  output [7:0]   io_pipe_phv_out_data_25,
  output [7:0]   io_pipe_phv_out_data_26,
  output [7:0]   io_pipe_phv_out_data_27,
  output [7:0]   io_pipe_phv_out_data_28,
  output [7:0]   io_pipe_phv_out_data_29,
  output [7:0]   io_pipe_phv_out_data_30,
  output [7:0]   io_pipe_phv_out_data_31,
  output [7:0]   io_pipe_phv_out_data_32,
  output [7:0]   io_pipe_phv_out_data_33,
  output [7:0]   io_pipe_phv_out_data_34,
  output [7:0]   io_pipe_phv_out_data_35,
  output [7:0]   io_pipe_phv_out_data_36,
  output [7:0]   io_pipe_phv_out_data_37,
  output [7:0]   io_pipe_phv_out_data_38,
  output [7:0]   io_pipe_phv_out_data_39,
  output [7:0]   io_pipe_phv_out_data_40,
  output [7:0]   io_pipe_phv_out_data_41,
  output [7:0]   io_pipe_phv_out_data_42,
  output [7:0]   io_pipe_phv_out_data_43,
  output [7:0]   io_pipe_phv_out_data_44,
  output [7:0]   io_pipe_phv_out_data_45,
  output [7:0]   io_pipe_phv_out_data_46,
  output [7:0]   io_pipe_phv_out_data_47,
  output [7:0]   io_pipe_phv_out_data_48,
  output [7:0]   io_pipe_phv_out_data_49,
  output [7:0]   io_pipe_phv_out_data_50,
  output [7:0]   io_pipe_phv_out_data_51,
  output [7:0]   io_pipe_phv_out_data_52,
  output [7:0]   io_pipe_phv_out_data_53,
  output [7:0]   io_pipe_phv_out_data_54,
  output [7:0]   io_pipe_phv_out_data_55,
  output [7:0]   io_pipe_phv_out_data_56,
  output [7:0]   io_pipe_phv_out_data_57,
  output [7:0]   io_pipe_phv_out_data_58,
  output [7:0]   io_pipe_phv_out_data_59,
  output [7:0]   io_pipe_phv_out_data_60,
  output [7:0]   io_pipe_phv_out_data_61,
  output [7:0]   io_pipe_phv_out_data_62,
  output [7:0]   io_pipe_phv_out_data_63,
  output [7:0]   io_pipe_phv_out_data_64,
  output [7:0]   io_pipe_phv_out_data_65,
  output [7:0]   io_pipe_phv_out_data_66,
  output [7:0]   io_pipe_phv_out_data_67,
  output [7:0]   io_pipe_phv_out_data_68,
  output [7:0]   io_pipe_phv_out_data_69,
  output [7:0]   io_pipe_phv_out_data_70,
  output [7:0]   io_pipe_phv_out_data_71,
  output [7:0]   io_pipe_phv_out_data_72,
  output [7:0]   io_pipe_phv_out_data_73,
  output [7:0]   io_pipe_phv_out_data_74,
  output [7:0]   io_pipe_phv_out_data_75,
  output [7:0]   io_pipe_phv_out_data_76,
  output [7:0]   io_pipe_phv_out_data_77,
  output [7:0]   io_pipe_phv_out_data_78,
  output [7:0]   io_pipe_phv_out_data_79,
  output [7:0]   io_pipe_phv_out_data_80,
  output [7:0]   io_pipe_phv_out_data_81,
  output [7:0]   io_pipe_phv_out_data_82,
  output [7:0]   io_pipe_phv_out_data_83,
  output [7:0]   io_pipe_phv_out_data_84,
  output [7:0]   io_pipe_phv_out_data_85,
  output [7:0]   io_pipe_phv_out_data_86,
  output [7:0]   io_pipe_phv_out_data_87,
  output [7:0]   io_pipe_phv_out_data_88,
  output [7:0]   io_pipe_phv_out_data_89,
  output [7:0]   io_pipe_phv_out_data_90,
  output [7:0]   io_pipe_phv_out_data_91,
  output [7:0]   io_pipe_phv_out_data_92,
  output [7:0]   io_pipe_phv_out_data_93,
  output [7:0]   io_pipe_phv_out_data_94,
  output [7:0]   io_pipe_phv_out_data_95,
  output [7:0]   io_pipe_phv_out_data_96,
  output [7:0]   io_pipe_phv_out_data_97,
  output [7:0]   io_pipe_phv_out_data_98,
  output [7:0]   io_pipe_phv_out_data_99,
  output [7:0]   io_pipe_phv_out_data_100,
  output [7:0]   io_pipe_phv_out_data_101,
  output [7:0]   io_pipe_phv_out_data_102,
  output [7:0]   io_pipe_phv_out_data_103,
  output [7:0]   io_pipe_phv_out_data_104,
  output [7:0]   io_pipe_phv_out_data_105,
  output [7:0]   io_pipe_phv_out_data_106,
  output [7:0]   io_pipe_phv_out_data_107,
  output [7:0]   io_pipe_phv_out_data_108,
  output [7:0]   io_pipe_phv_out_data_109,
  output [7:0]   io_pipe_phv_out_data_110,
  output [7:0]   io_pipe_phv_out_data_111,
  output [7:0]   io_pipe_phv_out_data_112,
  output [7:0]   io_pipe_phv_out_data_113,
  output [7:0]   io_pipe_phv_out_data_114,
  output [7:0]   io_pipe_phv_out_data_115,
  output [7:0]   io_pipe_phv_out_data_116,
  output [7:0]   io_pipe_phv_out_data_117,
  output [7:0]   io_pipe_phv_out_data_118,
  output [7:0]   io_pipe_phv_out_data_119,
  output [7:0]   io_pipe_phv_out_data_120,
  output [7:0]   io_pipe_phv_out_data_121,
  output [7:0]   io_pipe_phv_out_data_122,
  output [7:0]   io_pipe_phv_out_data_123,
  output [7:0]   io_pipe_phv_out_data_124,
  output [7:0]   io_pipe_phv_out_data_125,
  output [7:0]   io_pipe_phv_out_data_126,
  output [7:0]   io_pipe_phv_out_data_127,
  output [7:0]   io_pipe_phv_out_data_128,
  output [7:0]   io_pipe_phv_out_data_129,
  output [7:0]   io_pipe_phv_out_data_130,
  output [7:0]   io_pipe_phv_out_data_131,
  output [7:0]   io_pipe_phv_out_data_132,
  output [7:0]   io_pipe_phv_out_data_133,
  output [7:0]   io_pipe_phv_out_data_134,
  output [7:0]   io_pipe_phv_out_data_135,
  output [7:0]   io_pipe_phv_out_data_136,
  output [7:0]   io_pipe_phv_out_data_137,
  output [7:0]   io_pipe_phv_out_data_138,
  output [7:0]   io_pipe_phv_out_data_139,
  output [7:0]   io_pipe_phv_out_data_140,
  output [7:0]   io_pipe_phv_out_data_141,
  output [7:0]   io_pipe_phv_out_data_142,
  output [7:0]   io_pipe_phv_out_data_143,
  output [7:0]   io_pipe_phv_out_data_144,
  output [7:0]   io_pipe_phv_out_data_145,
  output [7:0]   io_pipe_phv_out_data_146,
  output [7:0]   io_pipe_phv_out_data_147,
  output [7:0]   io_pipe_phv_out_data_148,
  output [7:0]   io_pipe_phv_out_data_149,
  output [7:0]   io_pipe_phv_out_data_150,
  output [7:0]   io_pipe_phv_out_data_151,
  output [7:0]   io_pipe_phv_out_data_152,
  output [7:0]   io_pipe_phv_out_data_153,
  output [7:0]   io_pipe_phv_out_data_154,
  output [7:0]   io_pipe_phv_out_data_155,
  output [7:0]   io_pipe_phv_out_data_156,
  output [7:0]   io_pipe_phv_out_data_157,
  output [7:0]   io_pipe_phv_out_data_158,
  output [7:0]   io_pipe_phv_out_data_159,
  output [7:0]   io_pipe_phv_out_data_160,
  output [7:0]   io_pipe_phv_out_data_161,
  output [7:0]   io_pipe_phv_out_data_162,
  output [7:0]   io_pipe_phv_out_data_163,
  output [7:0]   io_pipe_phv_out_data_164,
  output [7:0]   io_pipe_phv_out_data_165,
  output [7:0]   io_pipe_phv_out_data_166,
  output [7:0]   io_pipe_phv_out_data_167,
  output [7:0]   io_pipe_phv_out_data_168,
  output [7:0]   io_pipe_phv_out_data_169,
  output [7:0]   io_pipe_phv_out_data_170,
  output [7:0]   io_pipe_phv_out_data_171,
  output [7:0]   io_pipe_phv_out_data_172,
  output [7:0]   io_pipe_phv_out_data_173,
  output [7:0]   io_pipe_phv_out_data_174,
  output [7:0]   io_pipe_phv_out_data_175,
  output [7:0]   io_pipe_phv_out_data_176,
  output [7:0]   io_pipe_phv_out_data_177,
  output [7:0]   io_pipe_phv_out_data_178,
  output [7:0]   io_pipe_phv_out_data_179,
  output [7:0]   io_pipe_phv_out_data_180,
  output [7:0]   io_pipe_phv_out_data_181,
  output [7:0]   io_pipe_phv_out_data_182,
  output [7:0]   io_pipe_phv_out_data_183,
  output [7:0]   io_pipe_phv_out_data_184,
  output [7:0]   io_pipe_phv_out_data_185,
  output [7:0]   io_pipe_phv_out_data_186,
  output [7:0]   io_pipe_phv_out_data_187,
  output [7:0]   io_pipe_phv_out_data_188,
  output [7:0]   io_pipe_phv_out_data_189,
  output [7:0]   io_pipe_phv_out_data_190,
  output [7:0]   io_pipe_phv_out_data_191,
  output [7:0]   io_pipe_phv_out_data_192,
  output [7:0]   io_pipe_phv_out_data_193,
  output [7:0]   io_pipe_phv_out_data_194,
  output [7:0]   io_pipe_phv_out_data_195,
  output [7:0]   io_pipe_phv_out_data_196,
  output [7:0]   io_pipe_phv_out_data_197,
  output [7:0]   io_pipe_phv_out_data_198,
  output [7:0]   io_pipe_phv_out_data_199,
  output [7:0]   io_pipe_phv_out_data_200,
  output [7:0]   io_pipe_phv_out_data_201,
  output [7:0]   io_pipe_phv_out_data_202,
  output [7:0]   io_pipe_phv_out_data_203,
  output [7:0]   io_pipe_phv_out_data_204,
  output [7:0]   io_pipe_phv_out_data_205,
  output [7:0]   io_pipe_phv_out_data_206,
  output [7:0]   io_pipe_phv_out_data_207,
  output [7:0]   io_pipe_phv_out_data_208,
  output [7:0]   io_pipe_phv_out_data_209,
  output [7:0]   io_pipe_phv_out_data_210,
  output [7:0]   io_pipe_phv_out_data_211,
  output [7:0]   io_pipe_phv_out_data_212,
  output [7:0]   io_pipe_phv_out_data_213,
  output [7:0]   io_pipe_phv_out_data_214,
  output [7:0]   io_pipe_phv_out_data_215,
  output [7:0]   io_pipe_phv_out_data_216,
  output [7:0]   io_pipe_phv_out_data_217,
  output [7:0]   io_pipe_phv_out_data_218,
  output [7:0]   io_pipe_phv_out_data_219,
  output [7:0]   io_pipe_phv_out_data_220,
  output [7:0]   io_pipe_phv_out_data_221,
  output [7:0]   io_pipe_phv_out_data_222,
  output [7:0]   io_pipe_phv_out_data_223,
  output [7:0]   io_pipe_phv_out_data_224,
  output [7:0]   io_pipe_phv_out_data_225,
  output [7:0]   io_pipe_phv_out_data_226,
  output [7:0]   io_pipe_phv_out_data_227,
  output [7:0]   io_pipe_phv_out_data_228,
  output [7:0]   io_pipe_phv_out_data_229,
  output [7:0]   io_pipe_phv_out_data_230,
  output [7:0]   io_pipe_phv_out_data_231,
  output [7:0]   io_pipe_phv_out_data_232,
  output [7:0]   io_pipe_phv_out_data_233,
  output [7:0]   io_pipe_phv_out_data_234,
  output [7:0]   io_pipe_phv_out_data_235,
  output [7:0]   io_pipe_phv_out_data_236,
  output [7:0]   io_pipe_phv_out_data_237,
  output [7:0]   io_pipe_phv_out_data_238,
  output [7:0]   io_pipe_phv_out_data_239,
  output [7:0]   io_pipe_phv_out_data_240,
  output [7:0]   io_pipe_phv_out_data_241,
  output [7:0]   io_pipe_phv_out_data_242,
  output [7:0]   io_pipe_phv_out_data_243,
  output [7:0]   io_pipe_phv_out_data_244,
  output [7:0]   io_pipe_phv_out_data_245,
  output [7:0]   io_pipe_phv_out_data_246,
  output [7:0]   io_pipe_phv_out_data_247,
  output [7:0]   io_pipe_phv_out_data_248,
  output [7:0]   io_pipe_phv_out_data_249,
  output [7:0]   io_pipe_phv_out_data_250,
  output [7:0]   io_pipe_phv_out_data_251,
  output [7:0]   io_pipe_phv_out_data_252,
  output [7:0]   io_pipe_phv_out_data_253,
  output [7:0]   io_pipe_phv_out_data_254,
  output [7:0]   io_pipe_phv_out_data_255,
  output [15:0]  io_pipe_phv_out_header_0,
  output [15:0]  io_pipe_phv_out_header_1,
  output [15:0]  io_pipe_phv_out_header_2,
  output [15:0]  io_pipe_phv_out_header_3,
  output [15:0]  io_pipe_phv_out_header_4,
  output [15:0]  io_pipe_phv_out_header_5,
  output [15:0]  io_pipe_phv_out_header_6,
  output [15:0]  io_pipe_phv_out_header_7,
  output [15:0]  io_pipe_phv_out_header_8,
  output [15:0]  io_pipe_phv_out_header_9,
  output [15:0]  io_pipe_phv_out_header_10,
  output [15:0]  io_pipe_phv_out_header_11,
  output [15:0]  io_pipe_phv_out_header_12,
  output [15:0]  io_pipe_phv_out_header_13,
  output [15:0]  io_pipe_phv_out_header_14,
  output [15:0]  io_pipe_phv_out_header_15,
  output [7:0]   io_pipe_phv_out_parse_current_state,
  output [7:0]   io_pipe_phv_out_parse_current_offset,
  output [15:0]  io_pipe_phv_out_parse_transition_field,
  output [3:0]   io_pipe_phv_out_next_processor_id,
  output         io_pipe_phv_out_next_config_id,
  output         io_pipe_phv_out_is_valid_processor,
  input          io_mod_hash_depth_mod,
  input          io_mod_config_id,
  input  [3:0]   io_mod_hash_depth,
  input  [191:0] io_key_in,
  output [191:0] io_key_out,
  output [7:0]   io_hash_val,
  output [3:0]   io_hash_val_cs
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  pipe1_clock; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_0; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_1; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_2; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_3; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_4; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_5; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_6; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_7; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_8; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_9; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_10; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_11; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_12; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_13; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_14; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_15; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_16; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_17; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_18; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_19; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_20; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_21; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_22; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_23; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_24; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_25; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_26; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_27; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_28; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_29; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_30; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_31; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_32; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_33; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_34; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_35; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_36; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_37; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_38; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_39; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_40; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_41; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_42; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_43; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_44; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_45; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_46; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_47; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_48; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_49; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_50; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_51; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_52; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_53; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_54; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_55; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_56; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_57; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_58; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_59; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_60; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_61; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_62; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_63; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_64; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_65; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_66; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_67; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_68; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_69; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_70; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_71; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_72; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_73; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_74; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_75; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_76; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_77; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_78; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_79; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_80; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_81; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_82; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_83; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_84; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_85; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_86; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_87; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_88; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_89; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_90; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_91; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_92; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_93; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_94; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_95; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_96; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_97; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_98; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_99; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_100; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_101; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_102; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_103; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_104; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_105; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_106; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_107; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_108; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_109; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_110; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_111; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_112; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_113; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_114; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_115; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_116; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_117; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_118; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_119; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_120; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_121; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_122; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_123; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_124; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_125; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_126; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_127; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_128; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_129; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_130; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_131; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_132; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_133; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_134; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_135; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_136; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_137; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_138; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_139; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_140; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_141; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_142; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_143; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_144; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_145; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_146; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_147; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_148; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_149; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_150; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_151; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_152; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_153; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_154; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_155; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_156; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_157; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_158; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_159; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_160; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_161; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_162; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_163; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_164; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_165; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_166; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_167; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_168; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_169; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_170; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_171; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_172; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_173; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_174; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_175; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_176; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_177; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_178; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_179; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_180; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_181; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_182; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_183; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_184; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_185; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_186; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_187; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_188; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_189; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_190; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_191; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_192; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_193; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_194; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_195; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_196; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_197; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_198; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_199; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_200; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_201; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_202; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_203; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_204; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_205; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_206; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_207; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_208; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_209; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_210; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_211; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_212; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_213; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_214; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_215; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_216; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_217; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_218; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_219; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_220; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_221; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_222; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_223; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_224; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_225; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_226; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_227; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_228; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_229; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_230; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_231; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_232; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_233; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_234; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_235; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_236; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_237; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_238; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_239; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_240; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_241; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_242; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_243; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_244; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_245; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_246; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_247; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_248; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_249; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_250; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_251; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_252; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_253; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_254; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_255; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_0; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_1; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_2; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_3; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_4; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_5; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_6; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_7; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_8; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_9; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_10; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_11; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_12; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_13; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_14; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_15; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_state; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_offset; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_parse_transition_field; // @[hash.scala 127:23]
  wire [3:0] pipe1_io_pipe_phv_in_next_processor_id; // @[hash.scala 127:23]
  wire  pipe1_io_pipe_phv_in_next_config_id; // @[hash.scala 127:23]
  wire  pipe1_io_pipe_phv_in_is_valid_processor; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_0; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_1; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_2; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_3; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_4; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_5; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_6; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_7; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_8; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_9; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_10; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_11; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_12; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_13; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_14; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_15; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_16; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_17; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_18; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_19; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_20; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_21; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_22; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_23; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_24; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_25; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_26; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_27; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_28; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_29; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_30; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_31; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_32; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_33; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_34; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_35; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_36; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_37; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_38; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_39; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_40; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_41; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_42; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_43; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_44; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_45; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_46; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_47; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_48; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_49; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_50; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_51; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_52; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_53; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_54; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_55; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_56; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_57; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_58; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_59; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_60; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_61; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_62; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_63; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_64; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_65; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_66; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_67; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_68; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_69; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_70; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_71; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_72; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_73; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_74; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_75; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_76; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_77; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_78; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_79; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_80; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_81; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_82; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_83; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_84; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_85; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_86; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_87; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_88; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_89; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_90; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_91; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_92; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_93; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_94; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_95; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_96; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_97; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_98; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_99; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_100; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_101; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_102; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_103; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_104; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_105; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_106; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_107; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_108; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_109; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_110; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_111; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_112; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_113; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_114; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_115; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_116; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_117; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_118; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_119; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_120; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_121; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_122; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_123; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_124; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_125; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_126; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_127; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_128; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_129; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_130; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_131; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_132; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_133; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_134; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_135; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_136; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_137; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_138; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_139; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_140; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_141; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_142; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_143; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_144; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_145; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_146; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_147; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_148; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_149; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_150; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_151; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_152; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_153; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_154; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_155; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_156; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_157; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_158; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_159; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_160; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_161; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_162; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_163; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_164; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_165; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_166; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_167; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_168; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_169; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_170; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_171; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_172; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_173; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_174; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_175; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_176; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_177; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_178; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_179; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_180; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_181; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_182; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_183; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_184; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_185; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_186; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_187; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_188; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_189; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_190; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_191; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_192; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_193; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_194; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_195; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_196; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_197; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_198; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_199; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_200; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_201; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_202; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_203; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_204; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_205; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_206; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_207; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_208; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_209; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_210; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_211; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_212; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_213; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_214; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_215; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_216; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_217; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_218; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_219; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_220; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_221; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_222; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_223; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_224; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_225; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_226; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_227; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_228; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_229; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_230; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_231; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_232; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_233; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_234; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_235; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_236; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_237; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_238; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_239; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_240; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_241; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_242; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_243; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_244; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_245; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_246; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_247; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_248; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_249; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_250; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_251; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_252; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_253; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_254; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_255; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_0; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_1; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_2; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_3; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_4; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_5; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_6; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_7; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_8; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_9; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_10; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_11; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_12; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_13; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_14; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_15; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_state; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_offset; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_parse_transition_field; // @[hash.scala 127:23]
  wire [3:0] pipe1_io_pipe_phv_out_next_processor_id; // @[hash.scala 127:23]
  wire  pipe1_io_pipe_phv_out_next_config_id; // @[hash.scala 127:23]
  wire  pipe1_io_pipe_phv_out_is_valid_processor; // @[hash.scala 127:23]
  wire [191:0] pipe1_io_key_in; // @[hash.scala 127:23]
  wire [191:0] pipe1_io_key_out; // @[hash.scala 127:23]
  wire [191:0] pipe1_io_sum_in; // @[hash.scala 127:23]
  wire [191:0] pipe1_io_sum_out; // @[hash.scala 127:23]
  wire  pipe2_clock; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_0; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_1; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_2; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_3; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_4; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_5; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_6; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_7; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_8; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_9; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_10; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_11; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_12; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_13; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_14; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_15; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_16; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_17; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_18; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_19; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_20; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_21; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_22; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_23; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_24; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_25; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_26; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_27; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_28; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_29; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_30; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_31; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_32; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_33; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_34; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_35; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_36; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_37; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_38; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_39; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_40; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_41; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_42; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_43; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_44; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_45; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_46; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_47; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_48; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_49; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_50; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_51; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_52; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_53; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_54; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_55; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_56; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_57; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_58; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_59; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_60; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_61; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_62; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_63; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_64; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_65; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_66; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_67; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_68; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_69; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_70; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_71; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_72; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_73; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_74; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_75; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_76; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_77; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_78; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_79; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_80; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_81; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_82; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_83; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_84; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_85; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_86; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_87; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_88; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_89; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_90; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_91; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_92; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_93; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_94; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_95; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_96; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_97; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_98; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_99; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_100; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_101; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_102; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_103; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_104; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_105; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_106; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_107; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_108; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_109; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_110; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_111; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_112; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_113; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_114; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_115; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_116; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_117; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_118; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_119; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_120; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_121; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_122; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_123; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_124; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_125; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_126; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_127; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_128; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_129; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_130; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_131; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_132; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_133; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_134; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_135; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_136; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_137; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_138; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_139; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_140; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_141; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_142; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_143; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_144; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_145; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_146; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_147; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_148; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_149; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_150; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_151; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_152; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_153; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_154; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_155; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_156; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_157; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_158; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_159; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_160; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_161; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_162; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_163; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_164; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_165; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_166; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_167; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_168; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_169; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_170; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_171; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_172; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_173; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_174; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_175; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_176; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_177; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_178; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_179; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_180; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_181; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_182; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_183; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_184; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_185; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_186; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_187; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_188; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_189; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_190; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_191; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_192; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_193; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_194; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_195; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_196; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_197; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_198; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_199; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_200; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_201; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_202; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_203; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_204; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_205; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_206; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_207; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_208; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_209; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_210; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_211; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_212; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_213; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_214; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_215; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_216; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_217; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_218; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_219; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_220; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_221; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_222; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_223; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_224; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_225; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_226; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_227; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_228; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_229; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_230; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_231; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_232; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_233; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_234; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_235; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_236; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_237; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_238; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_239; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_240; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_241; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_242; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_243; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_244; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_245; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_246; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_247; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_248; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_249; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_250; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_251; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_252; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_253; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_254; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_255; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_0; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_1; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_2; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_3; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_4; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_5; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_6; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_7; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_8; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_9; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_10; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_11; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_12; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_13; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_14; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_15; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_state; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_offset; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_parse_transition_field; // @[hash.scala 128:23]
  wire [3:0] pipe2_io_pipe_phv_in_next_processor_id; // @[hash.scala 128:23]
  wire  pipe2_io_pipe_phv_in_next_config_id; // @[hash.scala 128:23]
  wire  pipe2_io_pipe_phv_in_is_valid_processor; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_0; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_1; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_2; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_3; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_4; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_5; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_6; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_7; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_8; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_9; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_10; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_11; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_12; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_13; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_14; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_15; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_16; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_17; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_18; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_19; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_20; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_21; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_22; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_23; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_24; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_25; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_26; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_27; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_28; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_29; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_30; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_31; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_32; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_33; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_34; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_35; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_36; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_37; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_38; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_39; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_40; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_41; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_42; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_43; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_44; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_45; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_46; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_47; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_48; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_49; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_50; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_51; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_52; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_53; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_54; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_55; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_56; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_57; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_58; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_59; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_60; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_61; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_62; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_63; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_64; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_65; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_66; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_67; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_68; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_69; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_70; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_71; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_72; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_73; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_74; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_75; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_76; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_77; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_78; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_79; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_80; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_81; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_82; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_83; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_84; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_85; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_86; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_87; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_88; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_89; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_90; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_91; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_92; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_93; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_94; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_95; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_96; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_97; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_98; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_99; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_100; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_101; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_102; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_103; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_104; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_105; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_106; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_107; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_108; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_109; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_110; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_111; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_112; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_113; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_114; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_115; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_116; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_117; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_118; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_119; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_120; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_121; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_122; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_123; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_124; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_125; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_126; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_127; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_128; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_129; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_130; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_131; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_132; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_133; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_134; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_135; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_136; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_137; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_138; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_139; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_140; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_141; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_142; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_143; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_144; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_145; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_146; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_147; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_148; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_149; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_150; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_151; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_152; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_153; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_154; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_155; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_156; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_157; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_158; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_159; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_160; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_161; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_162; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_163; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_164; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_165; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_166; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_167; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_168; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_169; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_170; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_171; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_172; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_173; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_174; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_175; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_176; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_177; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_178; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_179; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_180; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_181; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_182; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_183; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_184; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_185; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_186; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_187; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_188; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_189; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_190; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_191; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_192; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_193; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_194; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_195; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_196; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_197; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_198; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_199; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_200; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_201; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_202; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_203; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_204; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_205; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_206; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_207; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_208; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_209; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_210; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_211; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_212; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_213; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_214; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_215; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_216; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_217; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_218; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_219; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_220; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_221; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_222; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_223; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_224; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_225; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_226; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_227; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_228; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_229; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_230; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_231; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_232; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_233; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_234; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_235; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_236; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_237; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_238; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_239; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_240; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_241; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_242; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_243; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_244; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_245; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_246; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_247; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_248; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_249; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_250; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_251; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_252; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_253; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_254; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_255; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_0; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_1; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_2; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_3; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_4; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_5; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_6; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_7; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_8; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_9; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_10; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_11; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_12; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_13; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_14; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_15; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_state; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_offset; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_parse_transition_field; // @[hash.scala 128:23]
  wire [3:0] pipe2_io_pipe_phv_out_next_processor_id; // @[hash.scala 128:23]
  wire  pipe2_io_pipe_phv_out_next_config_id; // @[hash.scala 128:23]
  wire  pipe2_io_pipe_phv_out_is_valid_processor; // @[hash.scala 128:23]
  wire [191:0] pipe2_io_key_in; // @[hash.scala 128:23]
  wire [191:0] pipe2_io_key_out; // @[hash.scala 128:23]
  wire [191:0] pipe2_io_sum_in; // @[hash.scala 128:23]
  wire [191:0] pipe2_io_sum_out; // @[hash.scala 128:23]
  wire  pipe3_clock; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_0; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_1; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_2; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_3; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_4; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_5; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_6; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_7; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_8; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_9; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_10; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_11; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_12; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_13; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_14; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_15; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_16; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_17; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_18; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_19; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_20; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_21; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_22; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_23; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_24; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_25; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_26; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_27; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_28; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_29; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_30; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_31; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_32; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_33; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_34; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_35; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_36; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_37; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_38; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_39; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_40; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_41; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_42; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_43; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_44; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_45; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_46; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_47; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_48; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_49; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_50; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_51; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_52; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_53; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_54; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_55; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_56; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_57; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_58; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_59; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_60; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_61; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_62; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_63; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_64; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_65; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_66; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_67; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_68; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_69; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_70; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_71; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_72; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_73; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_74; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_75; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_76; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_77; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_78; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_79; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_80; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_81; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_82; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_83; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_84; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_85; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_86; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_87; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_88; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_89; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_90; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_91; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_92; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_93; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_94; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_95; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_96; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_97; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_98; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_99; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_100; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_101; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_102; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_103; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_104; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_105; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_106; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_107; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_108; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_109; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_110; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_111; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_112; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_113; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_114; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_115; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_116; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_117; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_118; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_119; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_120; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_121; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_122; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_123; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_124; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_125; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_126; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_127; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_128; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_129; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_130; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_131; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_132; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_133; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_134; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_135; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_136; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_137; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_138; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_139; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_140; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_141; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_142; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_143; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_144; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_145; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_146; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_147; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_148; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_149; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_150; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_151; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_152; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_153; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_154; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_155; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_156; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_157; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_158; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_159; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_160; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_161; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_162; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_163; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_164; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_165; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_166; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_167; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_168; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_169; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_170; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_171; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_172; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_173; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_174; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_175; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_176; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_177; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_178; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_179; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_180; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_181; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_182; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_183; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_184; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_185; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_186; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_187; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_188; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_189; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_190; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_191; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_192; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_193; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_194; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_195; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_196; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_197; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_198; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_199; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_200; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_201; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_202; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_203; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_204; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_205; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_206; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_207; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_208; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_209; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_210; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_211; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_212; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_213; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_214; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_215; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_216; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_217; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_218; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_219; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_220; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_221; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_222; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_223; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_224; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_225; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_226; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_227; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_228; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_229; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_230; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_231; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_232; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_233; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_234; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_235; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_236; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_237; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_238; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_239; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_240; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_241; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_242; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_243; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_244; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_245; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_246; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_247; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_248; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_249; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_250; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_251; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_252; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_253; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_254; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_255; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_0; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_1; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_2; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_3; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_4; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_5; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_6; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_7; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_8; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_9; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_10; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_11; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_12; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_13; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_14; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_15; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_parse_current_state; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_parse_current_offset; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_parse_transition_field; // @[hash.scala 129:23]
  wire [3:0] pipe3_io_pipe_phv_in_next_processor_id; // @[hash.scala 129:23]
  wire  pipe3_io_pipe_phv_in_next_config_id; // @[hash.scala 129:23]
  wire  pipe3_io_pipe_phv_in_is_valid_processor; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_0; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_1; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_2; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_3; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_4; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_5; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_6; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_7; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_8; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_9; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_10; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_11; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_12; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_13; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_14; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_15; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_16; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_17; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_18; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_19; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_20; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_21; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_22; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_23; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_24; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_25; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_26; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_27; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_28; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_29; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_30; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_31; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_32; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_33; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_34; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_35; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_36; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_37; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_38; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_39; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_40; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_41; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_42; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_43; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_44; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_45; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_46; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_47; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_48; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_49; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_50; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_51; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_52; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_53; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_54; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_55; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_56; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_57; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_58; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_59; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_60; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_61; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_62; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_63; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_64; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_65; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_66; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_67; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_68; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_69; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_70; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_71; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_72; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_73; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_74; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_75; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_76; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_77; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_78; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_79; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_80; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_81; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_82; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_83; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_84; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_85; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_86; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_87; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_88; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_89; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_90; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_91; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_92; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_93; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_94; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_95; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_96; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_97; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_98; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_99; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_100; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_101; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_102; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_103; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_104; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_105; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_106; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_107; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_108; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_109; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_110; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_111; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_112; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_113; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_114; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_115; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_116; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_117; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_118; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_119; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_120; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_121; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_122; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_123; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_124; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_125; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_126; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_127; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_128; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_129; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_130; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_131; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_132; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_133; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_134; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_135; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_136; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_137; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_138; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_139; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_140; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_141; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_142; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_143; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_144; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_145; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_146; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_147; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_148; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_149; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_150; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_151; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_152; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_153; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_154; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_155; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_156; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_157; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_158; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_159; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_160; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_161; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_162; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_163; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_164; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_165; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_166; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_167; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_168; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_169; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_170; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_171; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_172; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_173; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_174; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_175; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_176; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_177; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_178; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_179; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_180; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_181; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_182; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_183; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_184; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_185; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_186; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_187; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_188; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_189; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_190; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_191; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_192; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_193; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_194; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_195; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_196; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_197; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_198; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_199; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_200; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_201; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_202; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_203; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_204; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_205; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_206; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_207; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_208; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_209; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_210; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_211; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_212; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_213; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_214; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_215; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_216; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_217; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_218; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_219; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_220; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_221; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_222; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_223; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_224; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_225; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_226; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_227; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_228; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_229; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_230; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_231; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_232; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_233; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_234; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_235; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_236; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_237; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_238; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_239; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_240; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_241; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_242; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_243; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_244; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_245; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_246; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_247; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_248; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_249; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_250; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_251; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_252; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_253; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_254; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_255; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_0; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_1; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_2; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_3; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_4; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_5; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_6; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_7; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_8; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_9; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_10; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_11; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_12; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_13; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_14; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_15; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_parse_current_state; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_parse_current_offset; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_parse_transition_field; // @[hash.scala 129:23]
  wire [3:0] pipe3_io_pipe_phv_out_next_processor_id; // @[hash.scala 129:23]
  wire  pipe3_io_pipe_phv_out_next_config_id; // @[hash.scala 129:23]
  wire  pipe3_io_pipe_phv_out_is_valid_processor; // @[hash.scala 129:23]
  wire [191:0] pipe3_io_key_in; // @[hash.scala 129:23]
  wire [191:0] pipe3_io_key_out; // @[hash.scala 129:23]
  wire [191:0] pipe3_io_sum_in; // @[hash.scala 129:23]
  wire [191:0] pipe3_io_sum_out; // @[hash.scala 129:23]
  wire  pipe4_clock; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_0; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_1; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_2; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_3; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_4; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_5; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_6; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_7; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_8; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_9; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_10; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_11; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_12; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_13; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_14; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_15; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_16; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_17; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_18; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_19; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_20; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_21; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_22; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_23; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_24; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_25; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_26; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_27; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_28; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_29; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_30; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_31; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_32; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_33; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_34; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_35; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_36; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_37; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_38; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_39; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_40; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_41; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_42; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_43; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_44; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_45; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_46; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_47; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_48; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_49; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_50; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_51; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_52; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_53; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_54; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_55; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_56; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_57; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_58; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_59; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_60; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_61; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_62; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_63; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_64; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_65; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_66; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_67; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_68; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_69; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_70; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_71; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_72; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_73; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_74; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_75; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_76; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_77; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_78; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_79; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_80; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_81; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_82; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_83; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_84; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_85; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_86; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_87; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_88; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_89; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_90; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_91; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_92; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_93; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_94; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_95; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_96; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_97; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_98; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_99; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_100; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_101; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_102; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_103; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_104; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_105; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_106; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_107; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_108; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_109; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_110; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_111; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_112; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_113; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_114; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_115; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_116; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_117; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_118; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_119; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_120; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_121; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_122; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_123; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_124; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_125; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_126; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_127; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_128; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_129; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_130; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_131; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_132; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_133; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_134; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_135; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_136; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_137; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_138; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_139; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_140; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_141; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_142; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_143; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_144; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_145; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_146; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_147; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_148; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_149; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_150; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_151; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_152; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_153; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_154; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_155; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_156; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_157; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_158; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_159; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_160; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_161; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_162; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_163; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_164; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_165; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_166; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_167; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_168; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_169; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_170; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_171; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_172; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_173; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_174; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_175; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_176; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_177; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_178; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_179; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_180; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_181; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_182; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_183; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_184; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_185; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_186; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_187; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_188; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_189; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_190; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_191; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_192; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_193; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_194; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_195; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_196; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_197; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_198; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_199; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_200; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_201; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_202; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_203; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_204; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_205; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_206; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_207; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_208; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_209; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_210; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_211; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_212; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_213; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_214; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_215; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_216; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_217; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_218; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_219; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_220; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_221; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_222; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_223; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_224; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_225; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_226; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_227; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_228; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_229; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_230; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_231; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_232; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_233; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_234; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_235; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_236; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_237; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_238; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_239; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_240; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_241; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_242; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_243; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_244; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_245; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_246; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_247; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_248; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_249; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_250; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_251; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_252; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_253; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_254; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_255; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_0; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_1; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_2; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_3; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_4; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_5; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_6; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_7; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_8; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_9; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_10; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_11; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_12; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_13; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_14; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_15; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_parse_current_state; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_parse_current_offset; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_parse_transition_field; // @[hash.scala 130:23]
  wire [3:0] pipe4_io_pipe_phv_in_next_processor_id; // @[hash.scala 130:23]
  wire  pipe4_io_pipe_phv_in_next_config_id; // @[hash.scala 130:23]
  wire  pipe4_io_pipe_phv_in_is_valid_processor; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_0; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_1; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_2; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_3; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_4; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_5; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_6; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_7; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_8; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_9; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_10; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_11; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_12; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_13; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_14; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_15; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_16; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_17; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_18; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_19; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_20; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_21; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_22; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_23; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_24; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_25; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_26; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_27; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_28; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_29; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_30; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_31; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_32; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_33; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_34; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_35; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_36; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_37; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_38; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_39; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_40; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_41; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_42; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_43; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_44; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_45; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_46; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_47; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_48; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_49; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_50; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_51; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_52; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_53; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_54; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_55; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_56; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_57; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_58; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_59; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_60; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_61; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_62; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_63; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_64; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_65; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_66; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_67; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_68; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_69; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_70; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_71; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_72; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_73; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_74; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_75; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_76; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_77; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_78; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_79; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_80; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_81; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_82; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_83; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_84; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_85; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_86; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_87; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_88; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_89; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_90; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_91; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_92; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_93; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_94; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_95; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_96; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_97; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_98; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_99; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_100; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_101; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_102; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_103; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_104; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_105; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_106; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_107; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_108; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_109; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_110; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_111; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_112; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_113; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_114; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_115; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_116; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_117; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_118; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_119; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_120; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_121; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_122; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_123; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_124; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_125; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_126; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_127; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_128; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_129; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_130; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_131; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_132; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_133; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_134; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_135; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_136; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_137; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_138; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_139; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_140; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_141; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_142; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_143; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_144; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_145; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_146; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_147; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_148; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_149; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_150; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_151; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_152; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_153; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_154; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_155; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_156; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_157; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_158; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_159; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_160; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_161; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_162; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_163; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_164; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_165; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_166; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_167; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_168; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_169; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_170; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_171; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_172; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_173; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_174; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_175; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_176; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_177; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_178; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_179; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_180; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_181; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_182; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_183; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_184; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_185; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_186; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_187; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_188; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_189; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_190; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_191; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_192; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_193; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_194; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_195; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_196; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_197; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_198; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_199; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_200; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_201; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_202; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_203; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_204; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_205; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_206; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_207; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_208; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_209; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_210; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_211; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_212; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_213; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_214; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_215; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_216; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_217; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_218; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_219; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_220; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_221; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_222; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_223; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_224; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_225; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_226; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_227; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_228; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_229; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_230; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_231; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_232; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_233; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_234; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_235; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_236; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_237; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_238; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_239; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_240; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_241; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_242; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_243; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_244; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_245; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_246; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_247; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_248; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_249; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_250; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_251; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_252; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_253; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_254; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_255; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_0; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_1; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_2; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_3; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_4; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_5; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_6; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_7; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_8; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_9; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_10; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_11; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_12; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_13; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_14; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_15; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_parse_current_state; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_parse_current_offset; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_parse_transition_field; // @[hash.scala 130:23]
  wire [3:0] pipe4_io_pipe_phv_out_next_processor_id; // @[hash.scala 130:23]
  wire  pipe4_io_pipe_phv_out_next_config_id; // @[hash.scala 130:23]
  wire  pipe4_io_pipe_phv_out_is_valid_processor; // @[hash.scala 130:23]
  wire [191:0] pipe4_io_key_in; // @[hash.scala 130:23]
  wire [191:0] pipe4_io_key_out; // @[hash.scala 130:23]
  wire [191:0] pipe4_io_sum_in; // @[hash.scala 130:23]
  wire [191:0] pipe4_io_sum_out; // @[hash.scala 130:23]
  wire  pipe5_clock; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_0; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_1; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_2; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_3; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_4; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_5; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_6; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_7; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_8; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_9; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_10; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_11; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_12; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_13; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_14; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_15; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_16; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_17; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_18; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_19; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_20; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_21; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_22; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_23; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_24; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_25; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_26; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_27; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_28; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_29; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_30; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_31; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_32; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_33; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_34; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_35; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_36; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_37; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_38; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_39; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_40; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_41; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_42; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_43; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_44; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_45; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_46; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_47; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_48; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_49; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_50; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_51; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_52; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_53; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_54; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_55; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_56; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_57; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_58; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_59; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_60; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_61; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_62; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_63; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_64; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_65; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_66; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_67; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_68; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_69; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_70; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_71; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_72; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_73; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_74; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_75; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_76; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_77; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_78; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_79; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_80; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_81; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_82; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_83; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_84; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_85; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_86; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_87; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_88; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_89; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_90; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_91; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_92; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_93; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_94; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_95; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_96; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_97; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_98; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_99; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_100; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_101; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_102; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_103; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_104; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_105; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_106; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_107; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_108; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_109; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_110; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_111; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_112; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_113; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_114; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_115; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_116; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_117; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_118; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_119; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_120; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_121; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_122; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_123; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_124; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_125; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_126; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_127; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_128; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_129; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_130; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_131; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_132; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_133; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_134; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_135; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_136; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_137; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_138; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_139; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_140; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_141; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_142; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_143; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_144; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_145; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_146; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_147; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_148; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_149; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_150; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_151; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_152; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_153; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_154; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_155; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_156; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_157; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_158; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_159; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_160; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_161; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_162; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_163; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_164; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_165; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_166; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_167; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_168; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_169; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_170; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_171; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_172; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_173; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_174; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_175; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_176; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_177; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_178; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_179; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_180; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_181; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_182; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_183; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_184; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_185; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_186; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_187; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_188; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_189; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_190; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_191; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_192; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_193; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_194; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_195; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_196; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_197; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_198; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_199; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_200; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_201; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_202; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_203; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_204; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_205; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_206; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_207; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_208; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_209; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_210; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_211; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_212; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_213; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_214; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_215; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_216; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_217; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_218; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_219; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_220; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_221; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_222; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_223; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_224; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_225; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_226; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_227; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_228; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_229; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_230; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_231; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_232; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_233; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_234; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_235; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_236; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_237; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_238; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_239; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_240; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_241; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_242; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_243; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_244; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_245; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_246; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_247; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_248; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_249; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_250; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_251; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_252; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_253; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_254; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_255; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_0; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_1; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_2; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_3; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_4; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_5; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_6; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_7; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_8; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_9; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_10; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_11; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_12; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_13; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_14; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_15; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_parse_current_state; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_parse_current_offset; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_parse_transition_field; // @[hash.scala 131:23]
  wire [3:0] pipe5_io_pipe_phv_in_next_processor_id; // @[hash.scala 131:23]
  wire  pipe5_io_pipe_phv_in_next_config_id; // @[hash.scala 131:23]
  wire  pipe5_io_pipe_phv_in_is_valid_processor; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_0; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_1; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_2; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_3; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_4; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_5; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_6; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_7; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_8; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_9; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_10; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_11; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_12; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_13; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_14; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_15; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_16; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_17; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_18; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_19; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_20; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_21; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_22; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_23; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_24; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_25; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_26; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_27; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_28; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_29; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_30; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_31; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_32; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_33; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_34; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_35; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_36; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_37; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_38; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_39; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_40; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_41; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_42; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_43; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_44; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_45; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_46; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_47; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_48; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_49; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_50; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_51; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_52; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_53; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_54; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_55; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_56; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_57; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_58; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_59; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_60; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_61; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_62; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_63; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_64; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_65; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_66; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_67; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_68; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_69; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_70; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_71; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_72; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_73; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_74; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_75; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_76; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_77; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_78; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_79; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_80; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_81; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_82; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_83; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_84; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_85; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_86; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_87; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_88; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_89; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_90; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_91; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_92; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_93; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_94; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_95; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_96; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_97; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_98; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_99; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_100; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_101; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_102; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_103; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_104; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_105; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_106; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_107; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_108; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_109; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_110; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_111; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_112; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_113; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_114; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_115; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_116; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_117; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_118; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_119; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_120; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_121; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_122; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_123; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_124; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_125; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_126; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_127; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_128; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_129; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_130; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_131; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_132; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_133; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_134; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_135; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_136; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_137; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_138; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_139; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_140; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_141; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_142; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_143; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_144; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_145; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_146; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_147; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_148; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_149; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_150; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_151; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_152; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_153; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_154; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_155; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_156; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_157; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_158; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_159; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_160; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_161; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_162; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_163; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_164; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_165; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_166; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_167; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_168; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_169; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_170; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_171; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_172; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_173; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_174; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_175; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_176; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_177; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_178; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_179; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_180; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_181; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_182; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_183; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_184; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_185; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_186; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_187; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_188; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_189; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_190; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_191; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_192; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_193; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_194; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_195; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_196; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_197; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_198; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_199; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_200; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_201; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_202; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_203; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_204; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_205; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_206; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_207; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_208; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_209; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_210; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_211; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_212; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_213; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_214; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_215; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_216; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_217; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_218; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_219; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_220; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_221; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_222; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_223; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_224; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_225; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_226; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_227; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_228; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_229; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_230; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_231; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_232; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_233; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_234; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_235; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_236; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_237; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_238; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_239; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_240; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_241; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_242; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_243; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_244; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_245; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_246; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_247; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_248; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_249; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_250; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_251; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_252; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_253; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_254; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_255; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_0; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_1; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_2; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_3; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_4; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_5; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_6; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_7; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_8; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_9; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_10; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_11; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_12; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_13; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_14; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_15; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_parse_current_state; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_parse_current_offset; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_parse_transition_field; // @[hash.scala 131:23]
  wire [3:0] pipe5_io_pipe_phv_out_next_processor_id; // @[hash.scala 131:23]
  wire  pipe5_io_pipe_phv_out_next_config_id; // @[hash.scala 131:23]
  wire  pipe5_io_pipe_phv_out_is_valid_processor; // @[hash.scala 131:23]
  wire [3:0] pipe5_io_hash_depth_0; // @[hash.scala 131:23]
  wire [3:0] pipe5_io_hash_depth_1; // @[hash.scala 131:23]
  wire [191:0] pipe5_io_key_in; // @[hash.scala 131:23]
  wire [191:0] pipe5_io_key_out; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_sum_in; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_sum_out; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_val_out; // @[hash.scala 131:23]
  wire  pipe6_clock; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_0; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_1; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_2; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_3; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_4; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_5; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_6; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_7; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_8; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_9; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_10; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_11; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_12; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_13; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_14; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_15; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_16; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_17; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_18; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_19; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_20; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_21; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_22; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_23; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_24; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_25; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_26; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_27; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_28; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_29; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_30; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_31; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_32; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_33; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_34; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_35; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_36; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_37; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_38; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_39; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_40; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_41; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_42; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_43; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_44; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_45; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_46; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_47; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_48; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_49; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_50; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_51; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_52; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_53; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_54; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_55; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_56; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_57; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_58; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_59; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_60; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_61; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_62; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_63; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_64; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_65; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_66; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_67; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_68; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_69; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_70; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_71; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_72; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_73; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_74; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_75; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_76; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_77; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_78; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_79; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_80; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_81; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_82; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_83; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_84; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_85; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_86; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_87; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_88; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_89; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_90; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_91; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_92; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_93; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_94; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_95; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_96; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_97; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_98; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_99; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_100; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_101; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_102; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_103; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_104; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_105; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_106; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_107; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_108; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_109; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_110; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_111; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_112; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_113; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_114; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_115; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_116; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_117; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_118; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_119; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_120; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_121; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_122; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_123; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_124; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_125; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_126; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_127; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_128; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_129; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_130; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_131; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_132; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_133; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_134; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_135; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_136; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_137; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_138; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_139; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_140; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_141; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_142; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_143; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_144; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_145; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_146; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_147; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_148; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_149; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_150; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_151; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_152; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_153; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_154; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_155; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_156; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_157; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_158; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_159; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_160; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_161; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_162; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_163; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_164; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_165; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_166; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_167; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_168; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_169; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_170; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_171; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_172; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_173; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_174; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_175; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_176; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_177; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_178; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_179; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_180; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_181; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_182; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_183; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_184; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_185; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_186; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_187; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_188; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_189; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_190; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_191; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_192; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_193; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_194; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_195; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_196; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_197; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_198; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_199; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_200; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_201; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_202; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_203; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_204; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_205; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_206; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_207; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_208; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_209; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_210; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_211; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_212; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_213; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_214; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_215; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_216; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_217; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_218; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_219; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_220; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_221; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_222; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_223; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_224; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_225; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_226; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_227; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_228; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_229; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_230; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_231; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_232; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_233; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_234; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_235; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_236; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_237; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_238; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_239; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_240; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_241; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_242; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_243; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_244; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_245; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_246; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_247; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_248; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_249; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_250; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_251; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_252; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_253; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_254; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_255; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_0; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_1; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_2; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_3; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_4; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_5; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_6; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_7; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_8; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_9; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_10; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_11; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_12; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_13; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_14; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_15; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_parse_current_state; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_parse_current_offset; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_parse_transition_field; // @[hash.scala 132:23]
  wire [3:0] pipe6_io_pipe_phv_in_next_processor_id; // @[hash.scala 132:23]
  wire  pipe6_io_pipe_phv_in_next_config_id; // @[hash.scala 132:23]
  wire  pipe6_io_pipe_phv_in_is_valid_processor; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_0; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_1; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_2; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_3; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_4; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_5; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_6; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_7; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_8; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_9; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_10; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_11; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_12; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_13; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_14; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_15; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_16; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_17; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_18; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_19; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_20; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_21; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_22; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_23; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_24; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_25; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_26; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_27; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_28; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_29; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_30; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_31; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_32; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_33; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_34; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_35; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_36; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_37; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_38; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_39; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_40; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_41; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_42; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_43; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_44; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_45; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_46; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_47; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_48; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_49; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_50; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_51; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_52; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_53; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_54; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_55; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_56; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_57; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_58; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_59; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_60; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_61; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_62; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_63; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_64; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_65; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_66; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_67; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_68; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_69; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_70; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_71; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_72; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_73; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_74; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_75; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_76; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_77; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_78; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_79; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_80; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_81; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_82; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_83; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_84; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_85; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_86; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_87; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_88; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_89; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_90; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_91; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_92; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_93; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_94; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_95; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_96; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_97; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_98; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_99; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_100; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_101; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_102; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_103; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_104; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_105; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_106; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_107; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_108; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_109; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_110; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_111; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_112; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_113; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_114; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_115; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_116; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_117; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_118; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_119; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_120; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_121; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_122; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_123; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_124; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_125; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_126; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_127; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_128; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_129; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_130; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_131; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_132; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_133; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_134; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_135; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_136; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_137; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_138; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_139; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_140; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_141; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_142; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_143; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_144; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_145; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_146; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_147; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_148; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_149; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_150; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_151; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_152; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_153; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_154; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_155; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_156; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_157; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_158; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_159; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_160; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_161; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_162; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_163; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_164; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_165; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_166; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_167; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_168; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_169; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_170; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_171; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_172; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_173; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_174; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_175; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_176; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_177; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_178; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_179; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_180; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_181; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_182; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_183; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_184; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_185; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_186; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_187; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_188; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_189; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_190; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_191; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_192; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_193; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_194; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_195; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_196; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_197; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_198; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_199; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_200; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_201; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_202; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_203; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_204; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_205; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_206; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_207; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_208; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_209; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_210; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_211; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_212; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_213; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_214; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_215; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_216; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_217; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_218; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_219; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_220; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_221; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_222; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_223; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_224; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_225; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_226; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_227; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_228; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_229; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_230; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_231; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_232; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_233; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_234; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_235; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_236; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_237; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_238; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_239; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_240; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_241; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_242; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_243; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_244; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_245; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_246; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_247; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_248; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_249; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_250; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_251; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_252; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_253; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_254; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_255; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_0; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_1; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_2; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_3; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_4; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_5; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_6; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_7; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_8; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_9; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_10; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_11; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_12; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_13; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_14; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_15; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_parse_current_state; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_parse_current_offset; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_parse_transition_field; // @[hash.scala 132:23]
  wire [3:0] pipe6_io_pipe_phv_out_next_processor_id; // @[hash.scala 132:23]
  wire  pipe6_io_pipe_phv_out_next_config_id; // @[hash.scala 132:23]
  wire  pipe6_io_pipe_phv_out_is_valid_processor; // @[hash.scala 132:23]
  wire [3:0] pipe6_io_hash_depth_0; // @[hash.scala 132:23]
  wire [3:0] pipe6_io_hash_depth_1; // @[hash.scala 132:23]
  wire [191:0] pipe6_io_key_in; // @[hash.scala 132:23]
  wire [191:0] pipe6_io_key_out; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_sum_in; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_sum_out; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_val_in; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_val_out; // @[hash.scala 132:23]
  wire  pipe7_clock; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_0; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_1; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_2; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_3; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_4; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_5; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_6; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_7; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_8; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_9; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_10; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_11; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_12; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_13; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_14; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_15; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_16; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_17; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_18; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_19; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_20; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_21; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_22; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_23; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_24; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_25; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_26; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_27; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_28; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_29; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_30; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_31; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_32; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_33; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_34; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_35; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_36; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_37; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_38; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_39; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_40; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_41; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_42; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_43; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_44; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_45; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_46; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_47; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_48; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_49; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_50; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_51; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_52; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_53; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_54; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_55; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_56; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_57; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_58; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_59; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_60; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_61; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_62; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_63; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_64; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_65; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_66; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_67; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_68; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_69; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_70; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_71; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_72; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_73; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_74; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_75; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_76; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_77; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_78; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_79; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_80; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_81; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_82; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_83; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_84; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_85; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_86; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_87; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_88; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_89; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_90; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_91; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_92; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_93; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_94; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_95; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_96; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_97; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_98; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_99; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_100; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_101; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_102; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_103; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_104; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_105; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_106; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_107; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_108; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_109; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_110; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_111; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_112; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_113; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_114; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_115; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_116; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_117; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_118; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_119; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_120; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_121; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_122; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_123; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_124; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_125; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_126; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_127; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_128; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_129; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_130; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_131; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_132; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_133; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_134; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_135; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_136; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_137; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_138; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_139; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_140; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_141; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_142; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_143; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_144; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_145; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_146; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_147; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_148; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_149; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_150; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_151; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_152; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_153; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_154; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_155; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_156; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_157; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_158; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_159; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_160; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_161; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_162; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_163; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_164; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_165; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_166; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_167; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_168; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_169; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_170; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_171; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_172; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_173; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_174; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_175; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_176; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_177; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_178; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_179; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_180; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_181; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_182; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_183; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_184; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_185; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_186; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_187; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_188; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_189; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_190; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_191; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_192; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_193; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_194; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_195; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_196; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_197; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_198; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_199; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_200; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_201; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_202; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_203; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_204; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_205; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_206; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_207; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_208; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_209; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_210; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_211; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_212; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_213; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_214; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_215; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_216; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_217; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_218; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_219; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_220; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_221; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_222; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_223; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_224; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_225; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_226; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_227; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_228; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_229; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_230; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_231; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_232; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_233; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_234; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_235; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_236; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_237; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_238; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_239; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_240; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_241; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_242; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_243; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_244; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_245; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_246; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_247; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_248; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_249; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_250; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_251; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_252; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_253; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_254; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_255; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_0; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_1; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_2; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_3; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_4; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_5; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_6; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_7; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_8; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_9; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_10; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_11; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_12; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_13; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_14; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_15; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_parse_current_state; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_parse_current_offset; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_parse_transition_field; // @[hash.scala 133:23]
  wire [3:0] pipe7_io_pipe_phv_in_next_processor_id; // @[hash.scala 133:23]
  wire  pipe7_io_pipe_phv_in_next_config_id; // @[hash.scala 133:23]
  wire  pipe7_io_pipe_phv_in_is_valid_processor; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_0; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_1; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_2; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_3; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_4; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_5; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_6; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_7; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_8; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_9; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_10; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_11; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_12; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_13; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_14; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_15; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_16; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_17; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_18; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_19; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_20; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_21; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_22; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_23; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_24; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_25; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_26; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_27; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_28; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_29; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_30; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_31; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_32; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_33; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_34; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_35; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_36; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_37; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_38; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_39; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_40; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_41; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_42; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_43; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_44; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_45; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_46; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_47; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_48; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_49; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_50; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_51; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_52; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_53; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_54; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_55; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_56; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_57; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_58; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_59; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_60; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_61; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_62; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_63; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_64; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_65; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_66; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_67; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_68; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_69; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_70; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_71; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_72; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_73; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_74; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_75; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_76; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_77; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_78; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_79; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_80; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_81; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_82; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_83; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_84; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_85; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_86; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_87; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_88; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_89; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_90; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_91; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_92; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_93; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_94; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_95; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_96; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_97; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_98; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_99; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_100; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_101; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_102; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_103; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_104; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_105; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_106; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_107; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_108; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_109; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_110; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_111; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_112; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_113; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_114; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_115; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_116; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_117; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_118; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_119; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_120; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_121; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_122; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_123; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_124; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_125; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_126; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_127; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_128; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_129; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_130; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_131; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_132; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_133; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_134; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_135; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_136; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_137; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_138; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_139; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_140; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_141; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_142; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_143; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_144; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_145; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_146; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_147; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_148; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_149; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_150; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_151; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_152; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_153; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_154; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_155; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_156; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_157; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_158; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_159; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_160; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_161; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_162; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_163; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_164; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_165; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_166; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_167; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_168; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_169; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_170; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_171; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_172; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_173; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_174; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_175; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_176; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_177; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_178; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_179; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_180; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_181; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_182; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_183; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_184; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_185; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_186; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_187; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_188; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_189; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_190; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_191; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_192; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_193; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_194; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_195; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_196; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_197; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_198; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_199; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_200; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_201; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_202; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_203; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_204; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_205; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_206; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_207; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_208; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_209; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_210; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_211; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_212; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_213; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_214; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_215; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_216; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_217; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_218; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_219; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_220; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_221; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_222; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_223; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_224; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_225; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_226; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_227; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_228; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_229; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_230; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_231; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_232; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_233; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_234; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_235; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_236; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_237; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_238; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_239; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_240; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_241; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_242; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_243; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_244; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_245; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_246; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_247; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_248; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_249; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_250; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_251; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_252; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_253; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_254; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_255; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_0; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_1; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_2; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_3; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_4; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_5; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_6; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_7; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_8; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_9; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_10; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_11; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_12; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_13; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_14; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_15; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_parse_current_state; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_parse_current_offset; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_parse_transition_field; // @[hash.scala 133:23]
  wire [3:0] pipe7_io_pipe_phv_out_next_processor_id; // @[hash.scala 133:23]
  wire  pipe7_io_pipe_phv_out_next_config_id; // @[hash.scala 133:23]
  wire  pipe7_io_pipe_phv_out_is_valid_processor; // @[hash.scala 133:23]
  wire [3:0] pipe7_io_hash_depth_0; // @[hash.scala 133:23]
  wire [3:0] pipe7_io_hash_depth_1; // @[hash.scala 133:23]
  wire [191:0] pipe7_io_key_in; // @[hash.scala 133:23]
  wire [191:0] pipe7_io_key_out; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_sum_in; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_sum_out; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_val_in; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_val_out; // @[hash.scala 133:23]
  wire  pipe8_clock; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_0; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_1; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_2; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_3; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_4; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_5; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_6; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_7; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_8; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_9; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_10; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_11; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_12; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_13; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_14; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_15; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_16; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_17; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_18; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_19; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_20; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_21; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_22; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_23; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_24; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_25; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_26; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_27; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_28; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_29; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_30; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_31; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_32; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_33; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_34; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_35; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_36; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_37; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_38; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_39; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_40; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_41; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_42; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_43; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_44; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_45; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_46; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_47; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_48; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_49; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_50; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_51; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_52; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_53; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_54; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_55; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_56; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_57; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_58; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_59; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_60; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_61; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_62; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_63; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_64; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_65; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_66; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_67; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_68; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_69; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_70; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_71; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_72; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_73; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_74; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_75; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_76; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_77; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_78; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_79; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_80; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_81; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_82; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_83; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_84; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_85; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_86; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_87; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_88; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_89; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_90; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_91; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_92; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_93; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_94; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_95; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_96; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_97; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_98; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_99; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_100; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_101; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_102; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_103; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_104; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_105; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_106; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_107; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_108; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_109; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_110; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_111; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_112; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_113; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_114; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_115; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_116; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_117; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_118; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_119; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_120; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_121; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_122; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_123; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_124; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_125; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_126; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_127; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_128; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_129; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_130; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_131; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_132; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_133; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_134; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_135; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_136; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_137; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_138; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_139; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_140; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_141; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_142; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_143; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_144; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_145; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_146; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_147; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_148; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_149; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_150; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_151; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_152; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_153; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_154; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_155; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_156; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_157; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_158; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_159; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_160; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_161; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_162; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_163; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_164; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_165; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_166; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_167; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_168; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_169; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_170; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_171; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_172; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_173; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_174; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_175; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_176; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_177; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_178; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_179; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_180; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_181; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_182; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_183; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_184; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_185; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_186; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_187; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_188; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_189; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_190; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_191; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_192; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_193; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_194; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_195; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_196; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_197; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_198; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_199; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_200; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_201; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_202; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_203; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_204; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_205; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_206; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_207; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_208; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_209; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_210; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_211; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_212; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_213; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_214; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_215; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_216; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_217; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_218; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_219; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_220; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_221; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_222; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_223; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_224; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_225; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_226; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_227; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_228; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_229; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_230; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_231; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_232; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_233; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_234; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_235; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_236; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_237; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_238; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_239; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_240; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_241; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_242; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_243; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_244; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_245; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_246; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_247; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_248; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_249; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_250; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_251; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_252; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_253; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_254; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_255; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_0; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_1; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_2; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_3; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_4; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_5; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_6; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_7; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_8; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_9; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_10; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_11; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_12; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_13; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_14; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_15; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_parse_current_state; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_parse_current_offset; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_parse_transition_field; // @[hash.scala 134:23]
  wire [3:0] pipe8_io_pipe_phv_in_next_processor_id; // @[hash.scala 134:23]
  wire  pipe8_io_pipe_phv_in_next_config_id; // @[hash.scala 134:23]
  wire  pipe8_io_pipe_phv_in_is_valid_processor; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_0; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_1; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_2; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_3; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_4; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_5; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_6; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_7; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_8; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_9; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_10; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_11; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_12; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_13; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_14; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_15; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_16; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_17; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_18; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_19; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_20; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_21; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_22; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_23; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_24; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_25; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_26; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_27; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_28; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_29; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_30; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_31; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_32; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_33; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_34; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_35; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_36; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_37; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_38; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_39; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_40; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_41; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_42; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_43; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_44; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_45; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_46; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_47; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_48; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_49; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_50; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_51; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_52; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_53; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_54; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_55; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_56; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_57; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_58; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_59; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_60; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_61; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_62; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_63; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_64; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_65; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_66; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_67; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_68; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_69; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_70; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_71; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_72; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_73; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_74; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_75; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_76; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_77; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_78; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_79; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_80; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_81; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_82; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_83; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_84; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_85; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_86; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_87; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_88; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_89; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_90; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_91; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_92; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_93; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_94; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_95; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_96; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_97; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_98; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_99; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_100; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_101; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_102; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_103; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_104; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_105; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_106; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_107; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_108; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_109; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_110; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_111; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_112; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_113; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_114; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_115; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_116; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_117; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_118; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_119; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_120; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_121; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_122; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_123; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_124; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_125; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_126; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_127; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_128; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_129; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_130; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_131; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_132; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_133; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_134; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_135; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_136; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_137; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_138; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_139; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_140; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_141; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_142; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_143; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_144; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_145; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_146; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_147; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_148; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_149; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_150; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_151; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_152; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_153; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_154; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_155; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_156; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_157; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_158; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_159; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_160; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_161; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_162; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_163; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_164; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_165; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_166; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_167; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_168; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_169; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_170; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_171; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_172; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_173; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_174; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_175; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_176; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_177; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_178; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_179; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_180; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_181; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_182; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_183; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_184; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_185; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_186; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_187; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_188; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_189; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_190; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_191; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_192; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_193; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_194; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_195; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_196; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_197; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_198; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_199; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_200; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_201; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_202; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_203; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_204; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_205; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_206; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_207; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_208; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_209; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_210; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_211; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_212; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_213; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_214; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_215; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_216; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_217; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_218; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_219; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_220; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_221; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_222; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_223; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_224; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_225; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_226; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_227; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_228; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_229; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_230; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_231; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_232; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_233; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_234; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_235; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_236; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_237; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_238; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_239; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_240; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_241; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_242; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_243; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_244; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_245; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_246; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_247; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_248; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_249; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_250; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_251; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_252; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_253; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_254; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_255; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_0; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_1; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_2; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_3; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_4; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_5; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_6; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_7; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_8; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_9; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_10; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_11; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_12; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_13; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_14; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_15; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_parse_current_state; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_parse_current_offset; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_parse_transition_field; // @[hash.scala 134:23]
  wire [3:0] pipe8_io_pipe_phv_out_next_processor_id; // @[hash.scala 134:23]
  wire  pipe8_io_pipe_phv_out_next_config_id; // @[hash.scala 134:23]
  wire  pipe8_io_pipe_phv_out_is_valid_processor; // @[hash.scala 134:23]
  wire [3:0] pipe8_io_hash_depth_0; // @[hash.scala 134:23]
  wire [3:0] pipe8_io_hash_depth_1; // @[hash.scala 134:23]
  wire [191:0] pipe8_io_key_in; // @[hash.scala 134:23]
  wire [191:0] pipe8_io_key_out; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_sum_in; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_sum_out; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_val_in; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_val_out; // @[hash.scala 134:23]
  reg [3:0] hash_depth_0; // @[hash.scala 18:26]
  reg [3:0] hash_depth_1; // @[hash.scala 18:26]
  HashSumLevel pipe1 ( // @[hash.scala 127:23]
    .clock(pipe1_clock),
    .io_pipe_phv_in_data_0(pipe1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe1_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe1_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe1_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe1_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe1_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe1_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe1_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe1_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe1_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe1_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe1_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe1_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe1_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe1_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe1_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe1_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe1_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe1_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe1_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe1_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe1_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe1_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe1_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe1_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe1_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe1_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe1_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe1_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe1_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe1_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe1_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe1_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe1_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe1_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe1_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe1_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe1_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe1_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe1_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe1_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe1_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe1_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe1_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe1_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe1_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe1_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe1_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe1_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe1_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe1_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe1_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe1_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe1_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe1_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe1_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe1_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe1_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe1_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe1_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe1_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe1_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe1_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe1_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe1_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe1_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe1_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe1_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe1_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe1_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe1_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe1_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe1_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe1_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe1_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe1_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe1_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe1_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe1_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe1_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe1_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe1_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe1_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe1_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe1_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe1_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe1_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe1_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe1_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe1_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe1_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe1_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe1_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe1_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe1_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe1_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe1_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe1_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe1_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe1_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe1_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe1_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe1_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe1_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe1_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe1_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe1_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe1_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe1_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe1_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe1_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe1_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe1_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe1_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe1_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe1_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe1_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe1_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe1_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe1_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe1_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe1_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe1_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe1_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe1_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe1_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe1_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe1_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe1_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe1_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe1_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe1_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe1_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe1_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe1_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe1_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe1_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe1_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe1_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe1_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe1_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe1_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe1_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe1_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe1_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe1_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe1_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe1_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe1_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe1_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe1_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe1_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe1_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe1_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe1_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe1_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe1_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe1_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe1_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe1_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe1_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe1_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe1_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe1_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe1_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe1_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe1_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe1_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe1_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe1_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe1_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe1_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe1_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe1_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe1_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe1_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe1_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe1_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe1_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe1_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe1_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe1_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe1_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe1_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe1_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe1_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe1_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe1_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe1_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe1_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe1_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe1_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe1_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe1_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe1_io_key_in),
    .io_key_out(pipe1_io_key_out),
    .io_sum_in(pipe1_io_sum_in),
    .io_sum_out(pipe1_io_sum_out)
  );
  HashSumLevel_1 pipe2 ( // @[hash.scala 128:23]
    .clock(pipe2_clock),
    .io_pipe_phv_in_data_0(pipe2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe2_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe2_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe2_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe2_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe2_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe2_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe2_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe2_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe2_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe2_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe2_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe2_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe2_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe2_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe2_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe2_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe2_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe2_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe2_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe2_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe2_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe2_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe2_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe2_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe2_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe2_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe2_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe2_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe2_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe2_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe2_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe2_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe2_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe2_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe2_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe2_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe2_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe2_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe2_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe2_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe2_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe2_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe2_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe2_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe2_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe2_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe2_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe2_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe2_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe2_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe2_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe2_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe2_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe2_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe2_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe2_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe2_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe2_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe2_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe2_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe2_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe2_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe2_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe2_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe2_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe2_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe2_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe2_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe2_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe2_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe2_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe2_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe2_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe2_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe2_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe2_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe2_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe2_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe2_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe2_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe2_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe2_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe2_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe2_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe2_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe2_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe2_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe2_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe2_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe2_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe2_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe2_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe2_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe2_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe2_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe2_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe2_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe2_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe2_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe2_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe2_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe2_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe2_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe2_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe2_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe2_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe2_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe2_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe2_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe2_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe2_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe2_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe2_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe2_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe2_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe2_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe2_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe2_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe2_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe2_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe2_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe2_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe2_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe2_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe2_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe2_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe2_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe2_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe2_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe2_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe2_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe2_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe2_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe2_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe2_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe2_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe2_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe2_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe2_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe2_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe2_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe2_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe2_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe2_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe2_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe2_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe2_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe2_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe2_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe2_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe2_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe2_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe2_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe2_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe2_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe2_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe2_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe2_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe2_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe2_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe2_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe2_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe2_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe2_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe2_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe2_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe2_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe2_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe2_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe2_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe2_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe2_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe2_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe2_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe2_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe2_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe2_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe2_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe2_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe2_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe2_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe2_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe2_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe2_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe2_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe2_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe2_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe2_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe2_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe2_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe2_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe2_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe2_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe2_io_key_in),
    .io_key_out(pipe2_io_key_out),
    .io_sum_in(pipe2_io_sum_in),
    .io_sum_out(pipe2_io_sum_out)
  );
  HashSumLevel_2 pipe3 ( // @[hash.scala 129:23]
    .clock(pipe3_clock),
    .io_pipe_phv_in_data_0(pipe3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe3_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe3_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe3_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe3_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe3_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe3_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe3_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe3_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe3_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe3_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe3_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe3_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe3_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe3_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe3_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe3_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe3_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe3_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe3_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe3_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe3_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe3_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe3_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe3_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe3_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe3_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe3_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe3_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe3_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe3_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe3_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe3_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe3_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe3_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe3_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe3_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe3_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe3_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe3_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe3_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe3_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe3_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe3_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe3_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe3_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe3_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe3_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe3_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe3_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe3_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe3_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe3_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe3_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe3_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe3_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe3_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe3_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe3_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe3_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe3_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe3_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe3_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe3_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe3_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe3_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe3_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe3_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe3_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe3_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe3_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe3_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe3_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe3_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe3_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe3_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe3_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe3_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe3_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe3_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe3_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe3_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe3_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe3_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe3_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe3_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe3_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe3_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe3_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe3_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe3_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe3_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe3_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe3_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe3_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe3_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe3_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe3_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe3_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe3_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe3_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe3_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe3_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe3_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe3_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe3_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe3_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe3_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe3_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe3_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe3_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe3_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe3_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe3_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe3_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe3_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe3_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe3_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe3_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe3_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe3_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe3_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe3_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe3_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe3_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe3_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe3_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe3_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe3_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe3_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe3_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe3_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe3_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe3_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe3_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe3_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe3_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe3_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe3_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe3_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe3_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe3_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe3_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe3_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe3_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe3_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe3_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe3_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe3_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe3_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe3_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe3_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe3_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe3_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe3_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe3_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe3_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe3_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe3_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe3_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe3_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe3_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe3_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe3_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe3_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe3_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe3_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe3_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe3_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe3_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe3_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe3_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe3_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe3_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe3_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe3_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe3_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe3_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe3_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe3_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe3_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe3_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe3_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe3_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe3_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe3_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe3_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe3_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe3_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe3_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe3_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe3_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe3_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe3_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe3_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe3_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe3_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe3_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe3_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe3_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe3_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe3_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe3_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe3_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe3_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe3_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe3_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe3_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe3_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe3_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe3_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe3_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe3_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe3_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe3_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe3_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe3_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe3_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe3_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe3_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe3_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe3_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe3_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe3_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe3_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe3_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe3_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe3_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe3_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe3_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe3_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe3_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe3_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe3_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe3_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe3_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe3_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe3_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe3_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe3_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe3_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe3_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe3_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe3_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe3_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe3_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe3_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe3_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe3_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe3_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe3_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe3_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe3_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe3_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe3_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe3_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe3_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe3_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe3_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe3_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe3_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe3_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe3_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe3_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe3_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe3_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe3_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe3_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe3_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe3_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe3_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe3_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe3_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe3_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe3_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe3_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe3_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe3_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe3_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe3_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe3_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe3_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe3_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe3_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe3_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe3_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe3_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe3_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe3_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe3_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe3_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe3_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe3_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe3_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe3_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe3_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe3_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe3_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe3_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe3_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe3_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe3_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe3_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe3_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe3_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe3_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe3_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe3_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe3_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe3_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe3_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe3_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe3_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe3_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe3_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe3_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe3_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe3_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe3_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe3_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe3_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe3_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe3_io_key_in),
    .io_key_out(pipe3_io_key_out),
    .io_sum_in(pipe3_io_sum_in),
    .io_sum_out(pipe3_io_sum_out)
  );
  HashSumLevel_3 pipe4 ( // @[hash.scala 130:23]
    .clock(pipe4_clock),
    .io_pipe_phv_in_data_0(pipe4_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe4_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe4_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe4_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe4_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe4_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe4_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe4_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe4_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe4_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe4_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe4_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe4_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe4_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe4_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe4_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe4_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe4_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe4_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe4_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe4_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe4_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe4_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe4_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe4_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe4_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe4_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe4_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe4_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe4_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe4_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe4_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe4_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe4_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe4_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe4_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe4_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe4_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe4_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe4_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe4_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe4_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe4_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe4_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe4_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe4_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe4_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe4_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe4_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe4_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe4_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe4_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe4_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe4_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe4_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe4_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe4_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe4_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe4_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe4_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe4_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe4_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe4_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe4_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe4_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe4_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe4_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe4_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe4_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe4_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe4_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe4_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe4_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe4_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe4_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe4_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe4_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe4_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe4_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe4_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe4_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe4_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe4_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe4_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe4_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe4_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe4_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe4_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe4_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe4_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe4_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe4_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe4_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe4_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe4_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe4_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe4_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe4_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe4_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe4_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe4_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe4_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe4_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe4_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe4_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe4_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe4_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe4_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe4_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe4_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe4_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe4_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe4_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe4_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe4_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe4_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe4_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe4_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe4_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe4_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe4_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe4_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe4_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe4_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe4_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe4_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe4_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe4_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe4_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe4_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe4_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe4_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe4_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe4_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe4_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe4_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe4_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe4_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe4_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe4_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe4_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe4_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe4_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe4_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe4_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe4_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe4_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe4_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe4_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe4_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe4_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe4_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe4_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe4_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe4_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe4_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe4_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe4_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe4_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe4_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe4_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe4_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe4_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe4_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe4_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe4_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe4_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe4_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe4_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe4_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe4_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe4_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe4_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe4_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe4_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe4_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe4_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe4_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe4_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe4_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe4_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe4_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe4_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe4_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe4_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe4_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe4_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe4_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe4_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe4_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe4_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe4_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe4_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe4_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe4_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe4_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe4_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe4_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe4_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe4_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe4_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe4_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe4_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe4_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe4_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe4_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe4_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe4_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe4_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe4_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe4_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe4_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe4_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe4_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe4_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe4_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe4_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe4_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe4_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe4_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe4_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe4_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe4_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe4_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe4_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe4_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe4_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe4_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe4_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe4_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe4_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe4_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe4_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe4_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe4_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe4_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe4_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe4_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe4_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe4_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe4_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe4_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe4_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe4_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe4_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe4_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe4_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe4_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe4_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe4_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe4_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe4_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe4_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe4_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe4_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe4_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe4_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe4_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe4_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe4_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe4_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe4_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe4_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe4_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe4_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe4_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe4_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe4_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe4_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe4_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe4_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe4_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe4_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe4_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe4_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe4_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe4_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe4_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe4_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe4_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe4_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe4_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe4_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe4_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe4_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe4_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe4_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe4_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe4_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe4_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe4_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe4_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe4_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe4_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe4_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe4_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe4_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe4_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe4_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe4_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe4_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe4_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe4_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe4_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe4_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe4_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe4_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe4_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe4_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe4_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe4_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe4_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe4_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe4_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe4_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe4_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe4_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe4_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe4_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe4_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe4_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe4_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe4_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe4_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe4_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe4_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe4_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe4_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe4_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe4_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe4_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe4_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe4_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe4_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe4_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe4_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe4_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe4_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe4_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe4_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe4_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe4_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe4_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe4_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe4_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe4_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe4_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe4_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe4_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe4_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe4_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe4_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe4_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe4_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe4_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe4_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe4_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe4_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe4_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe4_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe4_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe4_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe4_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe4_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe4_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe4_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe4_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe4_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe4_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe4_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe4_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe4_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe4_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe4_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe4_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe4_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe4_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe4_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe4_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe4_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe4_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe4_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe4_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe4_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe4_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe4_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe4_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe4_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe4_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe4_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe4_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe4_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe4_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe4_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe4_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe4_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe4_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe4_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe4_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe4_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe4_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe4_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe4_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe4_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe4_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe4_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe4_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe4_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe4_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe4_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe4_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe4_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe4_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe4_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe4_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe4_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe4_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe4_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe4_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe4_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe4_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe4_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe4_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe4_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe4_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe4_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe4_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe4_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe4_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe4_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe4_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe4_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe4_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe4_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe4_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe4_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe4_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe4_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe4_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe4_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe4_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe4_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe4_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe4_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe4_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe4_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe4_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe4_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe4_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe4_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe4_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe4_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe4_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe4_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe4_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe4_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe4_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe4_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe4_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe4_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe4_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe4_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe4_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe4_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe4_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe4_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe4_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe4_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe4_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe4_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe4_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe4_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe4_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe4_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe4_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe4_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe4_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe4_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe4_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe4_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe4_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe4_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe4_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe4_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe4_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe4_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe4_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe4_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe4_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe4_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe4_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe4_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe4_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe4_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe4_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe4_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe4_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe4_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe4_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe4_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe4_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe4_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe4_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe4_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe4_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe4_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe4_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe4_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe4_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe4_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe4_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe4_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe4_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe4_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe4_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe4_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe4_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe4_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe4_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe4_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe4_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe4_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe4_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe4_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe4_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe4_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe4_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe4_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe4_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe4_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe4_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe4_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe4_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe4_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe4_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe4_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe4_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe4_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe4_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe4_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe4_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe4_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe4_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe4_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe4_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe4_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe4_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe4_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe4_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe4_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe4_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe4_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe4_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe4_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe4_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe4_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe4_io_key_in),
    .io_key_out(pipe4_io_key_out),
    .io_sum_in(pipe4_io_sum_in),
    .io_sum_out(pipe4_io_sum_out)
  );
  HashReshapeLevel pipe5 ( // @[hash.scala 131:23]
    .clock(pipe5_clock),
    .io_pipe_phv_in_data_0(pipe5_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe5_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe5_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe5_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe5_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe5_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe5_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe5_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe5_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe5_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe5_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe5_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe5_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe5_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe5_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe5_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe5_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe5_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe5_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe5_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe5_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe5_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe5_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe5_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe5_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe5_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe5_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe5_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe5_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe5_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe5_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe5_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe5_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe5_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe5_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe5_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe5_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe5_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe5_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe5_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe5_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe5_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe5_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe5_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe5_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe5_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe5_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe5_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe5_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe5_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe5_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe5_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe5_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe5_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe5_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe5_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe5_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe5_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe5_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe5_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe5_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe5_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe5_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe5_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe5_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe5_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe5_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe5_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe5_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe5_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe5_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe5_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe5_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe5_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe5_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe5_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe5_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe5_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe5_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe5_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe5_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe5_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe5_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe5_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe5_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe5_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe5_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe5_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe5_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe5_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe5_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe5_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe5_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe5_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe5_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe5_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe5_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe5_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe5_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe5_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe5_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe5_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe5_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe5_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe5_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe5_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe5_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe5_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe5_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe5_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe5_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe5_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe5_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe5_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe5_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe5_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe5_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe5_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe5_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe5_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe5_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe5_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe5_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe5_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe5_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe5_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe5_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe5_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe5_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe5_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe5_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe5_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe5_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe5_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe5_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe5_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe5_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe5_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe5_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe5_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe5_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe5_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe5_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe5_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe5_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe5_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe5_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe5_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe5_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe5_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe5_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe5_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe5_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe5_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe5_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe5_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe5_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe5_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe5_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe5_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe5_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe5_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe5_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe5_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe5_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe5_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe5_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe5_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe5_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe5_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe5_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe5_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe5_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe5_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe5_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe5_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe5_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe5_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe5_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe5_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe5_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe5_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe5_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe5_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe5_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe5_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe5_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe5_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe5_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe5_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe5_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe5_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe5_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe5_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe5_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe5_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe5_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe5_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe5_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe5_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe5_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe5_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe5_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe5_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe5_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe5_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe5_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe5_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe5_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe5_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe5_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe5_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe5_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe5_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe5_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe5_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe5_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe5_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe5_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe5_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe5_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe5_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe5_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe5_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe5_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe5_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe5_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe5_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe5_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe5_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe5_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe5_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe5_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe5_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe5_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe5_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe5_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe5_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe5_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe5_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe5_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe5_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe5_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe5_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe5_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe5_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe5_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe5_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe5_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe5_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe5_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe5_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe5_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe5_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe5_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe5_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe5_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe5_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe5_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe5_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe5_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe5_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe5_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe5_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe5_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe5_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe5_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe5_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe5_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe5_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe5_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe5_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe5_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe5_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe5_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe5_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe5_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe5_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe5_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe5_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe5_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe5_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe5_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe5_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe5_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe5_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe5_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe5_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe5_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe5_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe5_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe5_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe5_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe5_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe5_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe5_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe5_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe5_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe5_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe5_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe5_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe5_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe5_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe5_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe5_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe5_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe5_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe5_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe5_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe5_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe5_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe5_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe5_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe5_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe5_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe5_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe5_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe5_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe5_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe5_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe5_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe5_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe5_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe5_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe5_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe5_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe5_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe5_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe5_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe5_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe5_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe5_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe5_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe5_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe5_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe5_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe5_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe5_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe5_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe5_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe5_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe5_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe5_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe5_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe5_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe5_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe5_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe5_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe5_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe5_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe5_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe5_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe5_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe5_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe5_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe5_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe5_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe5_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe5_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe5_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe5_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe5_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe5_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe5_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe5_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe5_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe5_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe5_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe5_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe5_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe5_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe5_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe5_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe5_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe5_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe5_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe5_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe5_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe5_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe5_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe5_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe5_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe5_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe5_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe5_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe5_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe5_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe5_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe5_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe5_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe5_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe5_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe5_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe5_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe5_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe5_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe5_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe5_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe5_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe5_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe5_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe5_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe5_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe5_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe5_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe5_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe5_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe5_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe5_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe5_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe5_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe5_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe5_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe5_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe5_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe5_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe5_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe5_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe5_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe5_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe5_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe5_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe5_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe5_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe5_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe5_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe5_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe5_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe5_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe5_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe5_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe5_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe5_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe5_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe5_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe5_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe5_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe5_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe5_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe5_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe5_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe5_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe5_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe5_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe5_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe5_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe5_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe5_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe5_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe5_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe5_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe5_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe5_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe5_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe5_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe5_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe5_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe5_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe5_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe5_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe5_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe5_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe5_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe5_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe5_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe5_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe5_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe5_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe5_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe5_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe5_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe5_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe5_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe5_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe5_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe5_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe5_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe5_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe5_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe5_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe5_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe5_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe5_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe5_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe5_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe5_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe5_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe5_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe5_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe5_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe5_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe5_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe5_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe5_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe5_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe5_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe5_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe5_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe5_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe5_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe5_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe5_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe5_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe5_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe5_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe5_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe5_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe5_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe5_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe5_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe5_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe5_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe5_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe5_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe5_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe5_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe5_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe5_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe5_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe5_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe5_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe5_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe5_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe5_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe5_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe5_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe5_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe5_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe5_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe5_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe5_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe5_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe5_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe5_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe5_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe5_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe5_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe5_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe5_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe5_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe5_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe5_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe5_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe5_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe5_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe5_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe5_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe5_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe5_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe5_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe5_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe5_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe5_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe5_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe5_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe5_io_pipe_phv_out_is_valid_processor),
    .io_hash_depth_0(pipe5_io_hash_depth_0),
    .io_hash_depth_1(pipe5_io_hash_depth_1),
    .io_key_in(pipe5_io_key_in),
    .io_key_out(pipe5_io_key_out),
    .io_sum_in(pipe5_io_sum_in),
    .io_sum_out(pipe5_io_sum_out),
    .io_val_out(pipe5_io_val_out)
  );
  HashReshapeLevel_1 pipe6 ( // @[hash.scala 132:23]
    .clock(pipe6_clock),
    .io_pipe_phv_in_data_0(pipe6_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe6_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe6_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe6_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe6_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe6_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe6_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe6_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe6_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe6_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe6_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe6_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe6_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe6_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe6_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe6_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe6_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe6_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe6_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe6_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe6_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe6_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe6_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe6_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe6_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe6_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe6_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe6_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe6_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe6_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe6_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe6_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe6_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe6_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe6_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe6_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe6_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe6_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe6_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe6_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe6_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe6_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe6_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe6_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe6_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe6_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe6_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe6_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe6_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe6_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe6_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe6_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe6_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe6_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe6_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe6_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe6_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe6_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe6_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe6_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe6_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe6_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe6_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe6_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe6_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe6_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe6_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe6_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe6_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe6_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe6_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe6_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe6_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe6_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe6_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe6_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe6_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe6_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe6_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe6_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe6_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe6_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe6_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe6_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe6_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe6_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe6_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe6_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe6_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe6_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe6_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe6_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe6_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe6_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe6_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe6_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe6_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe6_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe6_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe6_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe6_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe6_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe6_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe6_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe6_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe6_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe6_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe6_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe6_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe6_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe6_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe6_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe6_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe6_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe6_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe6_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe6_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe6_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe6_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe6_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe6_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe6_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe6_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe6_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe6_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe6_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe6_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe6_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe6_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe6_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe6_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe6_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe6_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe6_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe6_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe6_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe6_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe6_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe6_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe6_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe6_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe6_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe6_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe6_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe6_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe6_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe6_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe6_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe6_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe6_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe6_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe6_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe6_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe6_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe6_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe6_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe6_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe6_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe6_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe6_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe6_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe6_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe6_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe6_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe6_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe6_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe6_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe6_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe6_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe6_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe6_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe6_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe6_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe6_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe6_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe6_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe6_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe6_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe6_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe6_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe6_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe6_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe6_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe6_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe6_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe6_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe6_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe6_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe6_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe6_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe6_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe6_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe6_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe6_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe6_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe6_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe6_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe6_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe6_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe6_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe6_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe6_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe6_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe6_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe6_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe6_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe6_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe6_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe6_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe6_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe6_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe6_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe6_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe6_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe6_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe6_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe6_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe6_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe6_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe6_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe6_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe6_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe6_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe6_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe6_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe6_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe6_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe6_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe6_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe6_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe6_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe6_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe6_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe6_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe6_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe6_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe6_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe6_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe6_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe6_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe6_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe6_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe6_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe6_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe6_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe6_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe6_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe6_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe6_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe6_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe6_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe6_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe6_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe6_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe6_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe6_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe6_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe6_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe6_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe6_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe6_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe6_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe6_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe6_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe6_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe6_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe6_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe6_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe6_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe6_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe6_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe6_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe6_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe6_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe6_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe6_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe6_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe6_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe6_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe6_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe6_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe6_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe6_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe6_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe6_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe6_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe6_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe6_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe6_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe6_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe6_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe6_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe6_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe6_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe6_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe6_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe6_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe6_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe6_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe6_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe6_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe6_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe6_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe6_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe6_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe6_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe6_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe6_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe6_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe6_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe6_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe6_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe6_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe6_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe6_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe6_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe6_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe6_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe6_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe6_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe6_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe6_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe6_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe6_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe6_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe6_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe6_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe6_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe6_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe6_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe6_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe6_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe6_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe6_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe6_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe6_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe6_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe6_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe6_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe6_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe6_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe6_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe6_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe6_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe6_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe6_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe6_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe6_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe6_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe6_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe6_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe6_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe6_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe6_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe6_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe6_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe6_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe6_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe6_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe6_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe6_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe6_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe6_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe6_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe6_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe6_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe6_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe6_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe6_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe6_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe6_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe6_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe6_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe6_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe6_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe6_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe6_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe6_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe6_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe6_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe6_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe6_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe6_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe6_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe6_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe6_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe6_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe6_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe6_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe6_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe6_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe6_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe6_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe6_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe6_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe6_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe6_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe6_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe6_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe6_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe6_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe6_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe6_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe6_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe6_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe6_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe6_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe6_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe6_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe6_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe6_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe6_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe6_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe6_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe6_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe6_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe6_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe6_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe6_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe6_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe6_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe6_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe6_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe6_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe6_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe6_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe6_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe6_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe6_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe6_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe6_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe6_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe6_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe6_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe6_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe6_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe6_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe6_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe6_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe6_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe6_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe6_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe6_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe6_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe6_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe6_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe6_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe6_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe6_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe6_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe6_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe6_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe6_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe6_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe6_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe6_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe6_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe6_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe6_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe6_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe6_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe6_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe6_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe6_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe6_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe6_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe6_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe6_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe6_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe6_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe6_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe6_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe6_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe6_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe6_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe6_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe6_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe6_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe6_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe6_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe6_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe6_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe6_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe6_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe6_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe6_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe6_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe6_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe6_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe6_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe6_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe6_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe6_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe6_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe6_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe6_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe6_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe6_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe6_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe6_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe6_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe6_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe6_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe6_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe6_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe6_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe6_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe6_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe6_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe6_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe6_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe6_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe6_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe6_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe6_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe6_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe6_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe6_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe6_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe6_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe6_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe6_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe6_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe6_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe6_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe6_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe6_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe6_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe6_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe6_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe6_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe6_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe6_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe6_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe6_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe6_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe6_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe6_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe6_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe6_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe6_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe6_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe6_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe6_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe6_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe6_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe6_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe6_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe6_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe6_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe6_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe6_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe6_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe6_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe6_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe6_io_pipe_phv_out_is_valid_processor),
    .io_hash_depth_0(pipe6_io_hash_depth_0),
    .io_hash_depth_1(pipe6_io_hash_depth_1),
    .io_key_in(pipe6_io_key_in),
    .io_key_out(pipe6_io_key_out),
    .io_sum_in(pipe6_io_sum_in),
    .io_sum_out(pipe6_io_sum_out),
    .io_val_in(pipe6_io_val_in),
    .io_val_out(pipe6_io_val_out)
  );
  HashReshapeLevel_2 pipe7 ( // @[hash.scala 133:23]
    .clock(pipe7_clock),
    .io_pipe_phv_in_data_0(pipe7_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe7_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe7_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe7_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe7_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe7_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe7_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe7_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe7_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe7_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe7_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe7_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe7_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe7_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe7_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe7_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe7_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe7_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe7_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe7_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe7_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe7_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe7_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe7_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe7_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe7_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe7_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe7_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe7_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe7_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe7_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe7_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe7_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe7_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe7_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe7_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe7_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe7_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe7_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe7_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe7_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe7_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe7_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe7_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe7_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe7_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe7_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe7_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe7_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe7_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe7_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe7_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe7_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe7_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe7_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe7_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe7_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe7_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe7_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe7_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe7_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe7_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe7_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe7_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe7_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe7_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe7_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe7_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe7_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe7_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe7_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe7_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe7_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe7_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe7_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe7_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe7_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe7_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe7_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe7_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe7_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe7_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe7_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe7_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe7_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe7_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe7_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe7_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe7_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe7_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe7_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe7_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe7_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe7_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe7_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe7_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe7_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe7_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe7_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe7_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe7_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe7_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe7_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe7_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe7_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe7_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe7_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe7_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe7_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe7_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe7_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe7_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe7_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe7_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe7_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe7_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe7_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe7_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe7_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe7_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe7_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe7_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe7_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe7_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe7_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe7_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe7_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe7_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe7_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe7_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe7_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe7_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe7_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe7_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe7_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe7_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe7_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe7_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe7_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe7_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe7_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe7_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe7_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe7_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe7_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe7_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe7_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe7_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe7_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe7_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe7_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe7_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe7_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe7_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe7_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe7_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe7_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe7_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe7_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe7_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe7_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe7_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe7_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe7_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe7_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe7_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe7_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe7_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe7_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe7_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe7_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe7_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe7_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe7_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe7_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe7_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe7_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe7_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe7_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe7_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe7_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe7_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe7_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe7_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe7_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe7_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe7_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe7_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe7_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe7_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe7_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe7_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe7_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe7_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe7_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe7_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe7_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe7_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe7_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe7_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe7_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe7_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe7_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe7_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe7_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe7_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe7_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe7_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe7_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe7_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe7_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe7_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe7_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe7_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe7_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe7_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe7_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe7_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe7_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe7_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe7_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe7_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe7_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe7_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe7_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe7_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe7_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe7_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe7_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe7_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe7_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe7_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe7_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe7_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe7_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe7_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe7_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe7_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe7_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe7_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe7_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe7_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe7_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe7_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe7_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe7_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe7_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe7_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe7_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe7_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe7_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe7_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe7_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe7_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe7_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe7_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe7_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe7_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe7_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe7_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe7_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe7_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe7_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe7_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe7_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe7_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe7_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe7_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe7_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe7_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe7_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe7_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe7_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe7_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe7_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe7_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe7_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe7_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe7_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe7_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe7_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe7_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe7_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe7_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe7_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe7_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe7_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe7_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe7_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe7_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe7_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe7_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe7_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe7_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe7_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe7_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe7_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe7_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe7_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe7_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe7_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe7_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe7_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe7_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe7_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe7_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe7_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe7_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe7_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe7_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe7_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe7_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe7_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe7_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe7_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe7_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe7_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe7_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe7_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe7_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe7_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe7_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe7_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe7_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe7_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe7_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe7_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe7_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe7_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe7_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe7_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe7_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe7_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe7_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe7_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe7_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe7_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe7_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe7_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe7_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe7_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe7_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe7_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe7_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe7_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe7_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe7_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe7_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe7_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe7_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe7_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe7_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe7_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe7_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe7_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe7_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe7_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe7_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe7_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe7_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe7_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe7_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe7_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe7_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe7_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe7_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe7_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe7_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe7_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe7_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe7_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe7_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe7_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe7_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe7_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe7_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe7_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe7_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe7_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe7_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe7_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe7_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe7_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe7_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe7_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe7_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe7_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe7_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe7_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe7_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe7_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe7_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe7_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe7_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe7_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe7_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe7_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe7_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe7_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe7_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe7_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe7_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe7_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe7_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe7_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe7_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe7_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe7_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe7_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe7_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe7_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe7_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe7_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe7_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe7_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe7_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe7_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe7_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe7_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe7_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe7_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe7_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe7_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe7_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe7_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe7_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe7_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe7_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe7_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe7_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe7_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe7_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe7_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe7_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe7_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe7_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe7_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe7_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe7_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe7_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe7_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe7_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe7_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe7_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe7_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe7_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe7_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe7_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe7_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe7_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe7_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe7_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe7_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe7_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe7_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe7_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe7_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe7_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe7_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe7_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe7_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe7_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe7_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe7_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe7_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe7_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe7_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe7_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe7_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe7_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe7_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe7_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe7_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe7_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe7_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe7_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe7_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe7_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe7_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe7_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe7_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe7_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe7_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe7_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe7_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe7_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe7_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe7_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe7_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe7_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe7_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe7_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe7_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe7_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe7_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe7_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe7_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe7_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe7_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe7_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe7_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe7_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe7_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe7_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe7_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe7_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe7_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe7_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe7_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe7_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe7_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe7_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe7_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe7_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe7_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe7_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe7_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe7_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe7_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe7_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe7_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe7_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe7_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe7_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe7_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe7_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe7_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe7_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe7_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe7_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe7_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe7_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe7_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe7_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe7_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe7_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe7_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe7_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe7_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe7_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe7_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe7_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe7_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe7_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe7_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe7_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe7_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe7_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe7_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe7_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe7_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe7_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe7_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe7_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe7_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe7_io_pipe_phv_out_is_valid_processor),
    .io_hash_depth_0(pipe7_io_hash_depth_0),
    .io_hash_depth_1(pipe7_io_hash_depth_1),
    .io_key_in(pipe7_io_key_in),
    .io_key_out(pipe7_io_key_out),
    .io_sum_in(pipe7_io_sum_in),
    .io_sum_out(pipe7_io_sum_out),
    .io_val_in(pipe7_io_val_in),
    .io_val_out(pipe7_io_val_out)
  );
  HashReshapeLevel_3 pipe8 ( // @[hash.scala 134:23]
    .clock(pipe8_clock),
    .io_pipe_phv_in_data_0(pipe8_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe8_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe8_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe8_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe8_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe8_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe8_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe8_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe8_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe8_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe8_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe8_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe8_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe8_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe8_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe8_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe8_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe8_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe8_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe8_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe8_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe8_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe8_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe8_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe8_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe8_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe8_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe8_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe8_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe8_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe8_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe8_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe8_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe8_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe8_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe8_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe8_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe8_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe8_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe8_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe8_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe8_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe8_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe8_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe8_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe8_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe8_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe8_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe8_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe8_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe8_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe8_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe8_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe8_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe8_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe8_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe8_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe8_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe8_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe8_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe8_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe8_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe8_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe8_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe8_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe8_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe8_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe8_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe8_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe8_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe8_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe8_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe8_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe8_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe8_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe8_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe8_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe8_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe8_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe8_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe8_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe8_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe8_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe8_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe8_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe8_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe8_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe8_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe8_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe8_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe8_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe8_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe8_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe8_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe8_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe8_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe8_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe8_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe8_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe8_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe8_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe8_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe8_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe8_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe8_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe8_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe8_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe8_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe8_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe8_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe8_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe8_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe8_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe8_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe8_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe8_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe8_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe8_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe8_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe8_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe8_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe8_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe8_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe8_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe8_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe8_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe8_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe8_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe8_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe8_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe8_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe8_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe8_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe8_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe8_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe8_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe8_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe8_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe8_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe8_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe8_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe8_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe8_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe8_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe8_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe8_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe8_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe8_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe8_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe8_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe8_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe8_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe8_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe8_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe8_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe8_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe8_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe8_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe8_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe8_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe8_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe8_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe8_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe8_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe8_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe8_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe8_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe8_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe8_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe8_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe8_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe8_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe8_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe8_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe8_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe8_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe8_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe8_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe8_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe8_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe8_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe8_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe8_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe8_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe8_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe8_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe8_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe8_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe8_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe8_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe8_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe8_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe8_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe8_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe8_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe8_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe8_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe8_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe8_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe8_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe8_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe8_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe8_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe8_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe8_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe8_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe8_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe8_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe8_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe8_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe8_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe8_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe8_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe8_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe8_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe8_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe8_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe8_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe8_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe8_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe8_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe8_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe8_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe8_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe8_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe8_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe8_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe8_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe8_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe8_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe8_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe8_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe8_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe8_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe8_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe8_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe8_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe8_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe8_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe8_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe8_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe8_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe8_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe8_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe8_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe8_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe8_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe8_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe8_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe8_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe8_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe8_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe8_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe8_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe8_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe8_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe8_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe8_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe8_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe8_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe8_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe8_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe8_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe8_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe8_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe8_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe8_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe8_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe8_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe8_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe8_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe8_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe8_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe8_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe8_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe8_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe8_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe8_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe8_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe8_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe8_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe8_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe8_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe8_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe8_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe8_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe8_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe8_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe8_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe8_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe8_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe8_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe8_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe8_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe8_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe8_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe8_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe8_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe8_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe8_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe8_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe8_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe8_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe8_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe8_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe8_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe8_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe8_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe8_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe8_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe8_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe8_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe8_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe8_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe8_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe8_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe8_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe8_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe8_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe8_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe8_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe8_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe8_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe8_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe8_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe8_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe8_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe8_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe8_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe8_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe8_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe8_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe8_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe8_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe8_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe8_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe8_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe8_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe8_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe8_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe8_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe8_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe8_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe8_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe8_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe8_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe8_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe8_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe8_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe8_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe8_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe8_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe8_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe8_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe8_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe8_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe8_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe8_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe8_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe8_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe8_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe8_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe8_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe8_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe8_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe8_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe8_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe8_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe8_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe8_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe8_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe8_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe8_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe8_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe8_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe8_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe8_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe8_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe8_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe8_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe8_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe8_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe8_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe8_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe8_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe8_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe8_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe8_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe8_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe8_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe8_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe8_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe8_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe8_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe8_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe8_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe8_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe8_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe8_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe8_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe8_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe8_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe8_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe8_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe8_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe8_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe8_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe8_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe8_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe8_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe8_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe8_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe8_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe8_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe8_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe8_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe8_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe8_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe8_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe8_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe8_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe8_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe8_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe8_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe8_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe8_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe8_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe8_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe8_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe8_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe8_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe8_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe8_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe8_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe8_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe8_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe8_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe8_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe8_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe8_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe8_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe8_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe8_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe8_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe8_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe8_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe8_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe8_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe8_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe8_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe8_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe8_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe8_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe8_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe8_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe8_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe8_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe8_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe8_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe8_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe8_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe8_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe8_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe8_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe8_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe8_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe8_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe8_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe8_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe8_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe8_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe8_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe8_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe8_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe8_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe8_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe8_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe8_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe8_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe8_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe8_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe8_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe8_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe8_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe8_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe8_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe8_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe8_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe8_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe8_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe8_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe8_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe8_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe8_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe8_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe8_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe8_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe8_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe8_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe8_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe8_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe8_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe8_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe8_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe8_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe8_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe8_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe8_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe8_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe8_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe8_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe8_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe8_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe8_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe8_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe8_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe8_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe8_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe8_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe8_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe8_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe8_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe8_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe8_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe8_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe8_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe8_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe8_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe8_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe8_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe8_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe8_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe8_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe8_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe8_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe8_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe8_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe8_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe8_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe8_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe8_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe8_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe8_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe8_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe8_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe8_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe8_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe8_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe8_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe8_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe8_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe8_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe8_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe8_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe8_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe8_io_pipe_phv_out_is_valid_processor),
    .io_hash_depth_0(pipe8_io_hash_depth_0),
    .io_hash_depth_1(pipe8_io_hash_depth_1),
    .io_key_in(pipe8_io_key_in),
    .io_key_out(pipe8_io_key_out),
    .io_sum_in(pipe8_io_sum_in),
    .io_sum_out(pipe8_io_sum_out),
    .io_val_in(pipe8_io_val_in),
    .io_val_out(pipe8_io_val_out)
  );
  assign io_pipe_phv_out_data_0 = pipe8_io_pipe_phv_out_data_0; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_1 = pipe8_io_pipe_phv_out_data_1; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_2 = pipe8_io_pipe_phv_out_data_2; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_3 = pipe8_io_pipe_phv_out_data_3; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_4 = pipe8_io_pipe_phv_out_data_4; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_5 = pipe8_io_pipe_phv_out_data_5; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_6 = pipe8_io_pipe_phv_out_data_6; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_7 = pipe8_io_pipe_phv_out_data_7; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_8 = pipe8_io_pipe_phv_out_data_8; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_9 = pipe8_io_pipe_phv_out_data_9; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_10 = pipe8_io_pipe_phv_out_data_10; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_11 = pipe8_io_pipe_phv_out_data_11; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_12 = pipe8_io_pipe_phv_out_data_12; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_13 = pipe8_io_pipe_phv_out_data_13; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_14 = pipe8_io_pipe_phv_out_data_14; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_15 = pipe8_io_pipe_phv_out_data_15; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_16 = pipe8_io_pipe_phv_out_data_16; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_17 = pipe8_io_pipe_phv_out_data_17; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_18 = pipe8_io_pipe_phv_out_data_18; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_19 = pipe8_io_pipe_phv_out_data_19; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_20 = pipe8_io_pipe_phv_out_data_20; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_21 = pipe8_io_pipe_phv_out_data_21; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_22 = pipe8_io_pipe_phv_out_data_22; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_23 = pipe8_io_pipe_phv_out_data_23; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_24 = pipe8_io_pipe_phv_out_data_24; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_25 = pipe8_io_pipe_phv_out_data_25; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_26 = pipe8_io_pipe_phv_out_data_26; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_27 = pipe8_io_pipe_phv_out_data_27; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_28 = pipe8_io_pipe_phv_out_data_28; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_29 = pipe8_io_pipe_phv_out_data_29; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_30 = pipe8_io_pipe_phv_out_data_30; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_31 = pipe8_io_pipe_phv_out_data_31; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_32 = pipe8_io_pipe_phv_out_data_32; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_33 = pipe8_io_pipe_phv_out_data_33; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_34 = pipe8_io_pipe_phv_out_data_34; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_35 = pipe8_io_pipe_phv_out_data_35; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_36 = pipe8_io_pipe_phv_out_data_36; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_37 = pipe8_io_pipe_phv_out_data_37; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_38 = pipe8_io_pipe_phv_out_data_38; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_39 = pipe8_io_pipe_phv_out_data_39; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_40 = pipe8_io_pipe_phv_out_data_40; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_41 = pipe8_io_pipe_phv_out_data_41; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_42 = pipe8_io_pipe_phv_out_data_42; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_43 = pipe8_io_pipe_phv_out_data_43; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_44 = pipe8_io_pipe_phv_out_data_44; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_45 = pipe8_io_pipe_phv_out_data_45; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_46 = pipe8_io_pipe_phv_out_data_46; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_47 = pipe8_io_pipe_phv_out_data_47; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_48 = pipe8_io_pipe_phv_out_data_48; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_49 = pipe8_io_pipe_phv_out_data_49; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_50 = pipe8_io_pipe_phv_out_data_50; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_51 = pipe8_io_pipe_phv_out_data_51; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_52 = pipe8_io_pipe_phv_out_data_52; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_53 = pipe8_io_pipe_phv_out_data_53; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_54 = pipe8_io_pipe_phv_out_data_54; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_55 = pipe8_io_pipe_phv_out_data_55; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_56 = pipe8_io_pipe_phv_out_data_56; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_57 = pipe8_io_pipe_phv_out_data_57; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_58 = pipe8_io_pipe_phv_out_data_58; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_59 = pipe8_io_pipe_phv_out_data_59; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_60 = pipe8_io_pipe_phv_out_data_60; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_61 = pipe8_io_pipe_phv_out_data_61; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_62 = pipe8_io_pipe_phv_out_data_62; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_63 = pipe8_io_pipe_phv_out_data_63; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_64 = pipe8_io_pipe_phv_out_data_64; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_65 = pipe8_io_pipe_phv_out_data_65; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_66 = pipe8_io_pipe_phv_out_data_66; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_67 = pipe8_io_pipe_phv_out_data_67; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_68 = pipe8_io_pipe_phv_out_data_68; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_69 = pipe8_io_pipe_phv_out_data_69; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_70 = pipe8_io_pipe_phv_out_data_70; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_71 = pipe8_io_pipe_phv_out_data_71; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_72 = pipe8_io_pipe_phv_out_data_72; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_73 = pipe8_io_pipe_phv_out_data_73; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_74 = pipe8_io_pipe_phv_out_data_74; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_75 = pipe8_io_pipe_phv_out_data_75; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_76 = pipe8_io_pipe_phv_out_data_76; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_77 = pipe8_io_pipe_phv_out_data_77; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_78 = pipe8_io_pipe_phv_out_data_78; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_79 = pipe8_io_pipe_phv_out_data_79; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_80 = pipe8_io_pipe_phv_out_data_80; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_81 = pipe8_io_pipe_phv_out_data_81; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_82 = pipe8_io_pipe_phv_out_data_82; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_83 = pipe8_io_pipe_phv_out_data_83; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_84 = pipe8_io_pipe_phv_out_data_84; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_85 = pipe8_io_pipe_phv_out_data_85; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_86 = pipe8_io_pipe_phv_out_data_86; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_87 = pipe8_io_pipe_phv_out_data_87; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_88 = pipe8_io_pipe_phv_out_data_88; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_89 = pipe8_io_pipe_phv_out_data_89; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_90 = pipe8_io_pipe_phv_out_data_90; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_91 = pipe8_io_pipe_phv_out_data_91; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_92 = pipe8_io_pipe_phv_out_data_92; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_93 = pipe8_io_pipe_phv_out_data_93; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_94 = pipe8_io_pipe_phv_out_data_94; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_95 = pipe8_io_pipe_phv_out_data_95; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_96 = pipe8_io_pipe_phv_out_data_96; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_97 = pipe8_io_pipe_phv_out_data_97; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_98 = pipe8_io_pipe_phv_out_data_98; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_99 = pipe8_io_pipe_phv_out_data_99; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_100 = pipe8_io_pipe_phv_out_data_100; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_101 = pipe8_io_pipe_phv_out_data_101; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_102 = pipe8_io_pipe_phv_out_data_102; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_103 = pipe8_io_pipe_phv_out_data_103; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_104 = pipe8_io_pipe_phv_out_data_104; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_105 = pipe8_io_pipe_phv_out_data_105; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_106 = pipe8_io_pipe_phv_out_data_106; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_107 = pipe8_io_pipe_phv_out_data_107; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_108 = pipe8_io_pipe_phv_out_data_108; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_109 = pipe8_io_pipe_phv_out_data_109; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_110 = pipe8_io_pipe_phv_out_data_110; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_111 = pipe8_io_pipe_phv_out_data_111; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_112 = pipe8_io_pipe_phv_out_data_112; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_113 = pipe8_io_pipe_phv_out_data_113; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_114 = pipe8_io_pipe_phv_out_data_114; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_115 = pipe8_io_pipe_phv_out_data_115; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_116 = pipe8_io_pipe_phv_out_data_116; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_117 = pipe8_io_pipe_phv_out_data_117; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_118 = pipe8_io_pipe_phv_out_data_118; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_119 = pipe8_io_pipe_phv_out_data_119; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_120 = pipe8_io_pipe_phv_out_data_120; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_121 = pipe8_io_pipe_phv_out_data_121; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_122 = pipe8_io_pipe_phv_out_data_122; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_123 = pipe8_io_pipe_phv_out_data_123; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_124 = pipe8_io_pipe_phv_out_data_124; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_125 = pipe8_io_pipe_phv_out_data_125; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_126 = pipe8_io_pipe_phv_out_data_126; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_127 = pipe8_io_pipe_phv_out_data_127; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_128 = pipe8_io_pipe_phv_out_data_128; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_129 = pipe8_io_pipe_phv_out_data_129; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_130 = pipe8_io_pipe_phv_out_data_130; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_131 = pipe8_io_pipe_phv_out_data_131; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_132 = pipe8_io_pipe_phv_out_data_132; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_133 = pipe8_io_pipe_phv_out_data_133; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_134 = pipe8_io_pipe_phv_out_data_134; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_135 = pipe8_io_pipe_phv_out_data_135; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_136 = pipe8_io_pipe_phv_out_data_136; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_137 = pipe8_io_pipe_phv_out_data_137; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_138 = pipe8_io_pipe_phv_out_data_138; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_139 = pipe8_io_pipe_phv_out_data_139; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_140 = pipe8_io_pipe_phv_out_data_140; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_141 = pipe8_io_pipe_phv_out_data_141; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_142 = pipe8_io_pipe_phv_out_data_142; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_143 = pipe8_io_pipe_phv_out_data_143; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_144 = pipe8_io_pipe_phv_out_data_144; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_145 = pipe8_io_pipe_phv_out_data_145; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_146 = pipe8_io_pipe_phv_out_data_146; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_147 = pipe8_io_pipe_phv_out_data_147; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_148 = pipe8_io_pipe_phv_out_data_148; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_149 = pipe8_io_pipe_phv_out_data_149; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_150 = pipe8_io_pipe_phv_out_data_150; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_151 = pipe8_io_pipe_phv_out_data_151; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_152 = pipe8_io_pipe_phv_out_data_152; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_153 = pipe8_io_pipe_phv_out_data_153; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_154 = pipe8_io_pipe_phv_out_data_154; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_155 = pipe8_io_pipe_phv_out_data_155; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_156 = pipe8_io_pipe_phv_out_data_156; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_157 = pipe8_io_pipe_phv_out_data_157; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_158 = pipe8_io_pipe_phv_out_data_158; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_159 = pipe8_io_pipe_phv_out_data_159; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_160 = pipe8_io_pipe_phv_out_data_160; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_161 = pipe8_io_pipe_phv_out_data_161; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_162 = pipe8_io_pipe_phv_out_data_162; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_163 = pipe8_io_pipe_phv_out_data_163; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_164 = pipe8_io_pipe_phv_out_data_164; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_165 = pipe8_io_pipe_phv_out_data_165; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_166 = pipe8_io_pipe_phv_out_data_166; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_167 = pipe8_io_pipe_phv_out_data_167; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_168 = pipe8_io_pipe_phv_out_data_168; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_169 = pipe8_io_pipe_phv_out_data_169; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_170 = pipe8_io_pipe_phv_out_data_170; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_171 = pipe8_io_pipe_phv_out_data_171; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_172 = pipe8_io_pipe_phv_out_data_172; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_173 = pipe8_io_pipe_phv_out_data_173; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_174 = pipe8_io_pipe_phv_out_data_174; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_175 = pipe8_io_pipe_phv_out_data_175; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_176 = pipe8_io_pipe_phv_out_data_176; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_177 = pipe8_io_pipe_phv_out_data_177; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_178 = pipe8_io_pipe_phv_out_data_178; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_179 = pipe8_io_pipe_phv_out_data_179; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_180 = pipe8_io_pipe_phv_out_data_180; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_181 = pipe8_io_pipe_phv_out_data_181; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_182 = pipe8_io_pipe_phv_out_data_182; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_183 = pipe8_io_pipe_phv_out_data_183; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_184 = pipe8_io_pipe_phv_out_data_184; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_185 = pipe8_io_pipe_phv_out_data_185; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_186 = pipe8_io_pipe_phv_out_data_186; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_187 = pipe8_io_pipe_phv_out_data_187; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_188 = pipe8_io_pipe_phv_out_data_188; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_189 = pipe8_io_pipe_phv_out_data_189; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_190 = pipe8_io_pipe_phv_out_data_190; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_191 = pipe8_io_pipe_phv_out_data_191; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_192 = pipe8_io_pipe_phv_out_data_192; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_193 = pipe8_io_pipe_phv_out_data_193; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_194 = pipe8_io_pipe_phv_out_data_194; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_195 = pipe8_io_pipe_phv_out_data_195; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_196 = pipe8_io_pipe_phv_out_data_196; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_197 = pipe8_io_pipe_phv_out_data_197; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_198 = pipe8_io_pipe_phv_out_data_198; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_199 = pipe8_io_pipe_phv_out_data_199; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_200 = pipe8_io_pipe_phv_out_data_200; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_201 = pipe8_io_pipe_phv_out_data_201; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_202 = pipe8_io_pipe_phv_out_data_202; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_203 = pipe8_io_pipe_phv_out_data_203; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_204 = pipe8_io_pipe_phv_out_data_204; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_205 = pipe8_io_pipe_phv_out_data_205; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_206 = pipe8_io_pipe_phv_out_data_206; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_207 = pipe8_io_pipe_phv_out_data_207; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_208 = pipe8_io_pipe_phv_out_data_208; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_209 = pipe8_io_pipe_phv_out_data_209; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_210 = pipe8_io_pipe_phv_out_data_210; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_211 = pipe8_io_pipe_phv_out_data_211; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_212 = pipe8_io_pipe_phv_out_data_212; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_213 = pipe8_io_pipe_phv_out_data_213; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_214 = pipe8_io_pipe_phv_out_data_214; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_215 = pipe8_io_pipe_phv_out_data_215; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_216 = pipe8_io_pipe_phv_out_data_216; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_217 = pipe8_io_pipe_phv_out_data_217; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_218 = pipe8_io_pipe_phv_out_data_218; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_219 = pipe8_io_pipe_phv_out_data_219; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_220 = pipe8_io_pipe_phv_out_data_220; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_221 = pipe8_io_pipe_phv_out_data_221; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_222 = pipe8_io_pipe_phv_out_data_222; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_223 = pipe8_io_pipe_phv_out_data_223; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_224 = pipe8_io_pipe_phv_out_data_224; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_225 = pipe8_io_pipe_phv_out_data_225; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_226 = pipe8_io_pipe_phv_out_data_226; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_227 = pipe8_io_pipe_phv_out_data_227; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_228 = pipe8_io_pipe_phv_out_data_228; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_229 = pipe8_io_pipe_phv_out_data_229; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_230 = pipe8_io_pipe_phv_out_data_230; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_231 = pipe8_io_pipe_phv_out_data_231; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_232 = pipe8_io_pipe_phv_out_data_232; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_233 = pipe8_io_pipe_phv_out_data_233; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_234 = pipe8_io_pipe_phv_out_data_234; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_235 = pipe8_io_pipe_phv_out_data_235; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_236 = pipe8_io_pipe_phv_out_data_236; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_237 = pipe8_io_pipe_phv_out_data_237; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_238 = pipe8_io_pipe_phv_out_data_238; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_239 = pipe8_io_pipe_phv_out_data_239; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_240 = pipe8_io_pipe_phv_out_data_240; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_241 = pipe8_io_pipe_phv_out_data_241; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_242 = pipe8_io_pipe_phv_out_data_242; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_243 = pipe8_io_pipe_phv_out_data_243; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_244 = pipe8_io_pipe_phv_out_data_244; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_245 = pipe8_io_pipe_phv_out_data_245; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_246 = pipe8_io_pipe_phv_out_data_246; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_247 = pipe8_io_pipe_phv_out_data_247; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_248 = pipe8_io_pipe_phv_out_data_248; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_249 = pipe8_io_pipe_phv_out_data_249; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_250 = pipe8_io_pipe_phv_out_data_250; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_251 = pipe8_io_pipe_phv_out_data_251; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_252 = pipe8_io_pipe_phv_out_data_252; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_253 = pipe8_io_pipe_phv_out_data_253; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_254 = pipe8_io_pipe_phv_out_data_254; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_255 = pipe8_io_pipe_phv_out_data_255; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_0 = pipe8_io_pipe_phv_out_header_0; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_1 = pipe8_io_pipe_phv_out_header_1; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_2 = pipe8_io_pipe_phv_out_header_2; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_3 = pipe8_io_pipe_phv_out_header_3; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_4 = pipe8_io_pipe_phv_out_header_4; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_5 = pipe8_io_pipe_phv_out_header_5; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_6 = pipe8_io_pipe_phv_out_header_6; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_7 = pipe8_io_pipe_phv_out_header_7; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_8 = pipe8_io_pipe_phv_out_header_8; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_9 = pipe8_io_pipe_phv_out_header_9; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_10 = pipe8_io_pipe_phv_out_header_10; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_11 = pipe8_io_pipe_phv_out_header_11; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_12 = pipe8_io_pipe_phv_out_header_12; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_13 = pipe8_io_pipe_phv_out_header_13; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_14 = pipe8_io_pipe_phv_out_header_14; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_15 = pipe8_io_pipe_phv_out_header_15; // @[hash.scala 176:27]
  assign io_pipe_phv_out_parse_current_state = pipe8_io_pipe_phv_out_parse_current_state; // @[hash.scala 176:27]
  assign io_pipe_phv_out_parse_current_offset = pipe8_io_pipe_phv_out_parse_current_offset; // @[hash.scala 176:27]
  assign io_pipe_phv_out_parse_transition_field = pipe8_io_pipe_phv_out_parse_transition_field; // @[hash.scala 176:27]
  assign io_pipe_phv_out_next_processor_id = pipe8_io_pipe_phv_out_next_processor_id; // @[hash.scala 176:27]
  assign io_pipe_phv_out_next_config_id = pipe8_io_pipe_phv_out_next_config_id; // @[hash.scala 176:27]
  assign io_pipe_phv_out_is_valid_processor = pipe8_io_pipe_phv_out_is_valid_processor; // @[hash.scala 176:27]
  assign io_key_out = pipe8_io_key_out; // @[hash.scala 177:27]
  assign io_hash_val = pipe8_io_sum_out[7:0]; // @[hash.scala 178:46]
  assign io_hash_val_cs = pipe8_io_val_out[15:12]; // @[hash.scala 179:46]
  assign pipe1_clock = clock;
  assign pipe1_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_160 = io_pipe_phv_in_data_160; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_161 = io_pipe_phv_in_data_161; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_162 = io_pipe_phv_in_data_162; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_163 = io_pipe_phv_in_data_163; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_164 = io_pipe_phv_in_data_164; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_165 = io_pipe_phv_in_data_165; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_166 = io_pipe_phv_in_data_166; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_167 = io_pipe_phv_in_data_167; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_168 = io_pipe_phv_in_data_168; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_169 = io_pipe_phv_in_data_169; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_170 = io_pipe_phv_in_data_170; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_171 = io_pipe_phv_in_data_171; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_172 = io_pipe_phv_in_data_172; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_173 = io_pipe_phv_in_data_173; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_174 = io_pipe_phv_in_data_174; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_175 = io_pipe_phv_in_data_175; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_176 = io_pipe_phv_in_data_176; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_177 = io_pipe_phv_in_data_177; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_178 = io_pipe_phv_in_data_178; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_179 = io_pipe_phv_in_data_179; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_180 = io_pipe_phv_in_data_180; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_181 = io_pipe_phv_in_data_181; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_182 = io_pipe_phv_in_data_182; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_183 = io_pipe_phv_in_data_183; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_184 = io_pipe_phv_in_data_184; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_185 = io_pipe_phv_in_data_185; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_186 = io_pipe_phv_in_data_186; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_187 = io_pipe_phv_in_data_187; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_188 = io_pipe_phv_in_data_188; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_189 = io_pipe_phv_in_data_189; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_190 = io_pipe_phv_in_data_190; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_191 = io_pipe_phv_in_data_191; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_192 = io_pipe_phv_in_data_192; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_193 = io_pipe_phv_in_data_193; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_194 = io_pipe_phv_in_data_194; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_195 = io_pipe_phv_in_data_195; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_196 = io_pipe_phv_in_data_196; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_197 = io_pipe_phv_in_data_197; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_198 = io_pipe_phv_in_data_198; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_199 = io_pipe_phv_in_data_199; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_200 = io_pipe_phv_in_data_200; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_201 = io_pipe_phv_in_data_201; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_202 = io_pipe_phv_in_data_202; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_203 = io_pipe_phv_in_data_203; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_204 = io_pipe_phv_in_data_204; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_205 = io_pipe_phv_in_data_205; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_206 = io_pipe_phv_in_data_206; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_207 = io_pipe_phv_in_data_207; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_208 = io_pipe_phv_in_data_208; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_209 = io_pipe_phv_in_data_209; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_210 = io_pipe_phv_in_data_210; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_211 = io_pipe_phv_in_data_211; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_212 = io_pipe_phv_in_data_212; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_213 = io_pipe_phv_in_data_213; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_214 = io_pipe_phv_in_data_214; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_215 = io_pipe_phv_in_data_215; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_216 = io_pipe_phv_in_data_216; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_217 = io_pipe_phv_in_data_217; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_218 = io_pipe_phv_in_data_218; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_219 = io_pipe_phv_in_data_219; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_220 = io_pipe_phv_in_data_220; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_221 = io_pipe_phv_in_data_221; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_222 = io_pipe_phv_in_data_222; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_223 = io_pipe_phv_in_data_223; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_224 = io_pipe_phv_in_data_224; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_225 = io_pipe_phv_in_data_225; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_226 = io_pipe_phv_in_data_226; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_227 = io_pipe_phv_in_data_227; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_228 = io_pipe_phv_in_data_228; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_229 = io_pipe_phv_in_data_229; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_230 = io_pipe_phv_in_data_230; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_231 = io_pipe_phv_in_data_231; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_232 = io_pipe_phv_in_data_232; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_233 = io_pipe_phv_in_data_233; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_234 = io_pipe_phv_in_data_234; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_235 = io_pipe_phv_in_data_235; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_236 = io_pipe_phv_in_data_236; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_237 = io_pipe_phv_in_data_237; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_238 = io_pipe_phv_in_data_238; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_239 = io_pipe_phv_in_data_239; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_240 = io_pipe_phv_in_data_240; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_241 = io_pipe_phv_in_data_241; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_242 = io_pipe_phv_in_data_242; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_243 = io_pipe_phv_in_data_243; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_244 = io_pipe_phv_in_data_244; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_245 = io_pipe_phv_in_data_245; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_246 = io_pipe_phv_in_data_246; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_247 = io_pipe_phv_in_data_247; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_248 = io_pipe_phv_in_data_248; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_249 = io_pipe_phv_in_data_249; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_250 = io_pipe_phv_in_data_250; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_251 = io_pipe_phv_in_data_251; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_252 = io_pipe_phv_in_data_252; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_253 = io_pipe_phv_in_data_253; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_254 = io_pipe_phv_in_data_254; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_255 = io_pipe_phv_in_data_255; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[hash.scala 136:27]
  assign pipe1_io_key_in = io_key_in; // @[hash.scala 137:27]
  assign pipe1_io_sum_in = pipe1_io_key_in; // @[hash.scala 138:27]
  assign pipe2_clock = clock;
  assign pipe2_io_pipe_phv_in_data_0 = pipe1_io_pipe_phv_out_data_0; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_1 = pipe1_io_pipe_phv_out_data_1; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_2 = pipe1_io_pipe_phv_out_data_2; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_3 = pipe1_io_pipe_phv_out_data_3; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_4 = pipe1_io_pipe_phv_out_data_4; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_5 = pipe1_io_pipe_phv_out_data_5; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_6 = pipe1_io_pipe_phv_out_data_6; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_7 = pipe1_io_pipe_phv_out_data_7; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_8 = pipe1_io_pipe_phv_out_data_8; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_9 = pipe1_io_pipe_phv_out_data_9; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_10 = pipe1_io_pipe_phv_out_data_10; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_11 = pipe1_io_pipe_phv_out_data_11; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_12 = pipe1_io_pipe_phv_out_data_12; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_13 = pipe1_io_pipe_phv_out_data_13; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_14 = pipe1_io_pipe_phv_out_data_14; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_15 = pipe1_io_pipe_phv_out_data_15; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_16 = pipe1_io_pipe_phv_out_data_16; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_17 = pipe1_io_pipe_phv_out_data_17; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_18 = pipe1_io_pipe_phv_out_data_18; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_19 = pipe1_io_pipe_phv_out_data_19; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_20 = pipe1_io_pipe_phv_out_data_20; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_21 = pipe1_io_pipe_phv_out_data_21; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_22 = pipe1_io_pipe_phv_out_data_22; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_23 = pipe1_io_pipe_phv_out_data_23; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_24 = pipe1_io_pipe_phv_out_data_24; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_25 = pipe1_io_pipe_phv_out_data_25; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_26 = pipe1_io_pipe_phv_out_data_26; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_27 = pipe1_io_pipe_phv_out_data_27; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_28 = pipe1_io_pipe_phv_out_data_28; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_29 = pipe1_io_pipe_phv_out_data_29; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_30 = pipe1_io_pipe_phv_out_data_30; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_31 = pipe1_io_pipe_phv_out_data_31; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_32 = pipe1_io_pipe_phv_out_data_32; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_33 = pipe1_io_pipe_phv_out_data_33; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_34 = pipe1_io_pipe_phv_out_data_34; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_35 = pipe1_io_pipe_phv_out_data_35; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_36 = pipe1_io_pipe_phv_out_data_36; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_37 = pipe1_io_pipe_phv_out_data_37; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_38 = pipe1_io_pipe_phv_out_data_38; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_39 = pipe1_io_pipe_phv_out_data_39; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_40 = pipe1_io_pipe_phv_out_data_40; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_41 = pipe1_io_pipe_phv_out_data_41; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_42 = pipe1_io_pipe_phv_out_data_42; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_43 = pipe1_io_pipe_phv_out_data_43; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_44 = pipe1_io_pipe_phv_out_data_44; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_45 = pipe1_io_pipe_phv_out_data_45; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_46 = pipe1_io_pipe_phv_out_data_46; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_47 = pipe1_io_pipe_phv_out_data_47; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_48 = pipe1_io_pipe_phv_out_data_48; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_49 = pipe1_io_pipe_phv_out_data_49; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_50 = pipe1_io_pipe_phv_out_data_50; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_51 = pipe1_io_pipe_phv_out_data_51; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_52 = pipe1_io_pipe_phv_out_data_52; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_53 = pipe1_io_pipe_phv_out_data_53; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_54 = pipe1_io_pipe_phv_out_data_54; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_55 = pipe1_io_pipe_phv_out_data_55; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_56 = pipe1_io_pipe_phv_out_data_56; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_57 = pipe1_io_pipe_phv_out_data_57; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_58 = pipe1_io_pipe_phv_out_data_58; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_59 = pipe1_io_pipe_phv_out_data_59; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_60 = pipe1_io_pipe_phv_out_data_60; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_61 = pipe1_io_pipe_phv_out_data_61; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_62 = pipe1_io_pipe_phv_out_data_62; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_63 = pipe1_io_pipe_phv_out_data_63; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_64 = pipe1_io_pipe_phv_out_data_64; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_65 = pipe1_io_pipe_phv_out_data_65; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_66 = pipe1_io_pipe_phv_out_data_66; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_67 = pipe1_io_pipe_phv_out_data_67; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_68 = pipe1_io_pipe_phv_out_data_68; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_69 = pipe1_io_pipe_phv_out_data_69; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_70 = pipe1_io_pipe_phv_out_data_70; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_71 = pipe1_io_pipe_phv_out_data_71; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_72 = pipe1_io_pipe_phv_out_data_72; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_73 = pipe1_io_pipe_phv_out_data_73; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_74 = pipe1_io_pipe_phv_out_data_74; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_75 = pipe1_io_pipe_phv_out_data_75; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_76 = pipe1_io_pipe_phv_out_data_76; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_77 = pipe1_io_pipe_phv_out_data_77; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_78 = pipe1_io_pipe_phv_out_data_78; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_79 = pipe1_io_pipe_phv_out_data_79; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_80 = pipe1_io_pipe_phv_out_data_80; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_81 = pipe1_io_pipe_phv_out_data_81; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_82 = pipe1_io_pipe_phv_out_data_82; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_83 = pipe1_io_pipe_phv_out_data_83; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_84 = pipe1_io_pipe_phv_out_data_84; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_85 = pipe1_io_pipe_phv_out_data_85; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_86 = pipe1_io_pipe_phv_out_data_86; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_87 = pipe1_io_pipe_phv_out_data_87; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_88 = pipe1_io_pipe_phv_out_data_88; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_89 = pipe1_io_pipe_phv_out_data_89; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_90 = pipe1_io_pipe_phv_out_data_90; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_91 = pipe1_io_pipe_phv_out_data_91; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_92 = pipe1_io_pipe_phv_out_data_92; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_93 = pipe1_io_pipe_phv_out_data_93; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_94 = pipe1_io_pipe_phv_out_data_94; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_95 = pipe1_io_pipe_phv_out_data_95; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_96 = pipe1_io_pipe_phv_out_data_96; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_97 = pipe1_io_pipe_phv_out_data_97; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_98 = pipe1_io_pipe_phv_out_data_98; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_99 = pipe1_io_pipe_phv_out_data_99; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_100 = pipe1_io_pipe_phv_out_data_100; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_101 = pipe1_io_pipe_phv_out_data_101; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_102 = pipe1_io_pipe_phv_out_data_102; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_103 = pipe1_io_pipe_phv_out_data_103; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_104 = pipe1_io_pipe_phv_out_data_104; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_105 = pipe1_io_pipe_phv_out_data_105; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_106 = pipe1_io_pipe_phv_out_data_106; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_107 = pipe1_io_pipe_phv_out_data_107; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_108 = pipe1_io_pipe_phv_out_data_108; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_109 = pipe1_io_pipe_phv_out_data_109; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_110 = pipe1_io_pipe_phv_out_data_110; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_111 = pipe1_io_pipe_phv_out_data_111; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_112 = pipe1_io_pipe_phv_out_data_112; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_113 = pipe1_io_pipe_phv_out_data_113; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_114 = pipe1_io_pipe_phv_out_data_114; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_115 = pipe1_io_pipe_phv_out_data_115; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_116 = pipe1_io_pipe_phv_out_data_116; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_117 = pipe1_io_pipe_phv_out_data_117; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_118 = pipe1_io_pipe_phv_out_data_118; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_119 = pipe1_io_pipe_phv_out_data_119; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_120 = pipe1_io_pipe_phv_out_data_120; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_121 = pipe1_io_pipe_phv_out_data_121; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_122 = pipe1_io_pipe_phv_out_data_122; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_123 = pipe1_io_pipe_phv_out_data_123; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_124 = pipe1_io_pipe_phv_out_data_124; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_125 = pipe1_io_pipe_phv_out_data_125; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_126 = pipe1_io_pipe_phv_out_data_126; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_127 = pipe1_io_pipe_phv_out_data_127; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_128 = pipe1_io_pipe_phv_out_data_128; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_129 = pipe1_io_pipe_phv_out_data_129; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_130 = pipe1_io_pipe_phv_out_data_130; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_131 = pipe1_io_pipe_phv_out_data_131; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_132 = pipe1_io_pipe_phv_out_data_132; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_133 = pipe1_io_pipe_phv_out_data_133; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_134 = pipe1_io_pipe_phv_out_data_134; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_135 = pipe1_io_pipe_phv_out_data_135; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_136 = pipe1_io_pipe_phv_out_data_136; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_137 = pipe1_io_pipe_phv_out_data_137; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_138 = pipe1_io_pipe_phv_out_data_138; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_139 = pipe1_io_pipe_phv_out_data_139; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_140 = pipe1_io_pipe_phv_out_data_140; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_141 = pipe1_io_pipe_phv_out_data_141; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_142 = pipe1_io_pipe_phv_out_data_142; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_143 = pipe1_io_pipe_phv_out_data_143; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_144 = pipe1_io_pipe_phv_out_data_144; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_145 = pipe1_io_pipe_phv_out_data_145; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_146 = pipe1_io_pipe_phv_out_data_146; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_147 = pipe1_io_pipe_phv_out_data_147; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_148 = pipe1_io_pipe_phv_out_data_148; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_149 = pipe1_io_pipe_phv_out_data_149; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_150 = pipe1_io_pipe_phv_out_data_150; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_151 = pipe1_io_pipe_phv_out_data_151; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_152 = pipe1_io_pipe_phv_out_data_152; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_153 = pipe1_io_pipe_phv_out_data_153; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_154 = pipe1_io_pipe_phv_out_data_154; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_155 = pipe1_io_pipe_phv_out_data_155; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_156 = pipe1_io_pipe_phv_out_data_156; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_157 = pipe1_io_pipe_phv_out_data_157; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_158 = pipe1_io_pipe_phv_out_data_158; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_159 = pipe1_io_pipe_phv_out_data_159; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_160 = pipe1_io_pipe_phv_out_data_160; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_161 = pipe1_io_pipe_phv_out_data_161; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_162 = pipe1_io_pipe_phv_out_data_162; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_163 = pipe1_io_pipe_phv_out_data_163; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_164 = pipe1_io_pipe_phv_out_data_164; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_165 = pipe1_io_pipe_phv_out_data_165; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_166 = pipe1_io_pipe_phv_out_data_166; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_167 = pipe1_io_pipe_phv_out_data_167; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_168 = pipe1_io_pipe_phv_out_data_168; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_169 = pipe1_io_pipe_phv_out_data_169; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_170 = pipe1_io_pipe_phv_out_data_170; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_171 = pipe1_io_pipe_phv_out_data_171; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_172 = pipe1_io_pipe_phv_out_data_172; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_173 = pipe1_io_pipe_phv_out_data_173; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_174 = pipe1_io_pipe_phv_out_data_174; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_175 = pipe1_io_pipe_phv_out_data_175; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_176 = pipe1_io_pipe_phv_out_data_176; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_177 = pipe1_io_pipe_phv_out_data_177; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_178 = pipe1_io_pipe_phv_out_data_178; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_179 = pipe1_io_pipe_phv_out_data_179; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_180 = pipe1_io_pipe_phv_out_data_180; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_181 = pipe1_io_pipe_phv_out_data_181; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_182 = pipe1_io_pipe_phv_out_data_182; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_183 = pipe1_io_pipe_phv_out_data_183; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_184 = pipe1_io_pipe_phv_out_data_184; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_185 = pipe1_io_pipe_phv_out_data_185; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_186 = pipe1_io_pipe_phv_out_data_186; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_187 = pipe1_io_pipe_phv_out_data_187; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_188 = pipe1_io_pipe_phv_out_data_188; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_189 = pipe1_io_pipe_phv_out_data_189; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_190 = pipe1_io_pipe_phv_out_data_190; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_191 = pipe1_io_pipe_phv_out_data_191; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_192 = pipe1_io_pipe_phv_out_data_192; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_193 = pipe1_io_pipe_phv_out_data_193; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_194 = pipe1_io_pipe_phv_out_data_194; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_195 = pipe1_io_pipe_phv_out_data_195; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_196 = pipe1_io_pipe_phv_out_data_196; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_197 = pipe1_io_pipe_phv_out_data_197; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_198 = pipe1_io_pipe_phv_out_data_198; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_199 = pipe1_io_pipe_phv_out_data_199; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_200 = pipe1_io_pipe_phv_out_data_200; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_201 = pipe1_io_pipe_phv_out_data_201; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_202 = pipe1_io_pipe_phv_out_data_202; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_203 = pipe1_io_pipe_phv_out_data_203; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_204 = pipe1_io_pipe_phv_out_data_204; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_205 = pipe1_io_pipe_phv_out_data_205; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_206 = pipe1_io_pipe_phv_out_data_206; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_207 = pipe1_io_pipe_phv_out_data_207; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_208 = pipe1_io_pipe_phv_out_data_208; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_209 = pipe1_io_pipe_phv_out_data_209; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_210 = pipe1_io_pipe_phv_out_data_210; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_211 = pipe1_io_pipe_phv_out_data_211; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_212 = pipe1_io_pipe_phv_out_data_212; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_213 = pipe1_io_pipe_phv_out_data_213; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_214 = pipe1_io_pipe_phv_out_data_214; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_215 = pipe1_io_pipe_phv_out_data_215; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_216 = pipe1_io_pipe_phv_out_data_216; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_217 = pipe1_io_pipe_phv_out_data_217; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_218 = pipe1_io_pipe_phv_out_data_218; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_219 = pipe1_io_pipe_phv_out_data_219; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_220 = pipe1_io_pipe_phv_out_data_220; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_221 = pipe1_io_pipe_phv_out_data_221; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_222 = pipe1_io_pipe_phv_out_data_222; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_223 = pipe1_io_pipe_phv_out_data_223; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_224 = pipe1_io_pipe_phv_out_data_224; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_225 = pipe1_io_pipe_phv_out_data_225; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_226 = pipe1_io_pipe_phv_out_data_226; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_227 = pipe1_io_pipe_phv_out_data_227; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_228 = pipe1_io_pipe_phv_out_data_228; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_229 = pipe1_io_pipe_phv_out_data_229; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_230 = pipe1_io_pipe_phv_out_data_230; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_231 = pipe1_io_pipe_phv_out_data_231; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_232 = pipe1_io_pipe_phv_out_data_232; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_233 = pipe1_io_pipe_phv_out_data_233; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_234 = pipe1_io_pipe_phv_out_data_234; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_235 = pipe1_io_pipe_phv_out_data_235; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_236 = pipe1_io_pipe_phv_out_data_236; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_237 = pipe1_io_pipe_phv_out_data_237; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_238 = pipe1_io_pipe_phv_out_data_238; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_239 = pipe1_io_pipe_phv_out_data_239; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_240 = pipe1_io_pipe_phv_out_data_240; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_241 = pipe1_io_pipe_phv_out_data_241; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_242 = pipe1_io_pipe_phv_out_data_242; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_243 = pipe1_io_pipe_phv_out_data_243; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_244 = pipe1_io_pipe_phv_out_data_244; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_245 = pipe1_io_pipe_phv_out_data_245; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_246 = pipe1_io_pipe_phv_out_data_246; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_247 = pipe1_io_pipe_phv_out_data_247; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_248 = pipe1_io_pipe_phv_out_data_248; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_249 = pipe1_io_pipe_phv_out_data_249; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_250 = pipe1_io_pipe_phv_out_data_250; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_251 = pipe1_io_pipe_phv_out_data_251; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_252 = pipe1_io_pipe_phv_out_data_252; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_253 = pipe1_io_pipe_phv_out_data_253; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_254 = pipe1_io_pipe_phv_out_data_254; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_255 = pipe1_io_pipe_phv_out_data_255; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_0 = pipe1_io_pipe_phv_out_header_0; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_1 = pipe1_io_pipe_phv_out_header_1; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_2 = pipe1_io_pipe_phv_out_header_2; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_3 = pipe1_io_pipe_phv_out_header_3; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_4 = pipe1_io_pipe_phv_out_header_4; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_5 = pipe1_io_pipe_phv_out_header_5; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_6 = pipe1_io_pipe_phv_out_header_6; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_7 = pipe1_io_pipe_phv_out_header_7; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_8 = pipe1_io_pipe_phv_out_header_8; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_9 = pipe1_io_pipe_phv_out_header_9; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_10 = pipe1_io_pipe_phv_out_header_10; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_11 = pipe1_io_pipe_phv_out_header_11; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_12 = pipe1_io_pipe_phv_out_header_12; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_13 = pipe1_io_pipe_phv_out_header_13; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_14 = pipe1_io_pipe_phv_out_header_14; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_15 = pipe1_io_pipe_phv_out_header_15; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_parse_current_state = pipe1_io_pipe_phv_out_parse_current_state; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_parse_current_offset = pipe1_io_pipe_phv_out_parse_current_offset; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_parse_transition_field = pipe1_io_pipe_phv_out_parse_transition_field; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_next_processor_id = pipe1_io_pipe_phv_out_next_processor_id; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_next_config_id = pipe1_io_pipe_phv_out_next_config_id; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_is_valid_processor = pipe1_io_pipe_phv_out_is_valid_processor; // @[hash.scala 140:27]
  assign pipe2_io_key_in = pipe1_io_key_out; // @[hash.scala 141:27]
  assign pipe2_io_sum_in = pipe1_io_sum_out; // @[hash.scala 142:27]
  assign pipe3_clock = clock;
  assign pipe3_io_pipe_phv_in_data_0 = pipe2_io_pipe_phv_out_data_0; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_1 = pipe2_io_pipe_phv_out_data_1; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_2 = pipe2_io_pipe_phv_out_data_2; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_3 = pipe2_io_pipe_phv_out_data_3; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_4 = pipe2_io_pipe_phv_out_data_4; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_5 = pipe2_io_pipe_phv_out_data_5; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_6 = pipe2_io_pipe_phv_out_data_6; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_7 = pipe2_io_pipe_phv_out_data_7; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_8 = pipe2_io_pipe_phv_out_data_8; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_9 = pipe2_io_pipe_phv_out_data_9; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_10 = pipe2_io_pipe_phv_out_data_10; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_11 = pipe2_io_pipe_phv_out_data_11; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_12 = pipe2_io_pipe_phv_out_data_12; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_13 = pipe2_io_pipe_phv_out_data_13; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_14 = pipe2_io_pipe_phv_out_data_14; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_15 = pipe2_io_pipe_phv_out_data_15; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_16 = pipe2_io_pipe_phv_out_data_16; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_17 = pipe2_io_pipe_phv_out_data_17; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_18 = pipe2_io_pipe_phv_out_data_18; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_19 = pipe2_io_pipe_phv_out_data_19; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_20 = pipe2_io_pipe_phv_out_data_20; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_21 = pipe2_io_pipe_phv_out_data_21; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_22 = pipe2_io_pipe_phv_out_data_22; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_23 = pipe2_io_pipe_phv_out_data_23; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_24 = pipe2_io_pipe_phv_out_data_24; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_25 = pipe2_io_pipe_phv_out_data_25; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_26 = pipe2_io_pipe_phv_out_data_26; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_27 = pipe2_io_pipe_phv_out_data_27; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_28 = pipe2_io_pipe_phv_out_data_28; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_29 = pipe2_io_pipe_phv_out_data_29; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_30 = pipe2_io_pipe_phv_out_data_30; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_31 = pipe2_io_pipe_phv_out_data_31; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_32 = pipe2_io_pipe_phv_out_data_32; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_33 = pipe2_io_pipe_phv_out_data_33; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_34 = pipe2_io_pipe_phv_out_data_34; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_35 = pipe2_io_pipe_phv_out_data_35; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_36 = pipe2_io_pipe_phv_out_data_36; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_37 = pipe2_io_pipe_phv_out_data_37; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_38 = pipe2_io_pipe_phv_out_data_38; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_39 = pipe2_io_pipe_phv_out_data_39; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_40 = pipe2_io_pipe_phv_out_data_40; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_41 = pipe2_io_pipe_phv_out_data_41; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_42 = pipe2_io_pipe_phv_out_data_42; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_43 = pipe2_io_pipe_phv_out_data_43; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_44 = pipe2_io_pipe_phv_out_data_44; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_45 = pipe2_io_pipe_phv_out_data_45; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_46 = pipe2_io_pipe_phv_out_data_46; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_47 = pipe2_io_pipe_phv_out_data_47; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_48 = pipe2_io_pipe_phv_out_data_48; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_49 = pipe2_io_pipe_phv_out_data_49; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_50 = pipe2_io_pipe_phv_out_data_50; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_51 = pipe2_io_pipe_phv_out_data_51; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_52 = pipe2_io_pipe_phv_out_data_52; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_53 = pipe2_io_pipe_phv_out_data_53; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_54 = pipe2_io_pipe_phv_out_data_54; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_55 = pipe2_io_pipe_phv_out_data_55; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_56 = pipe2_io_pipe_phv_out_data_56; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_57 = pipe2_io_pipe_phv_out_data_57; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_58 = pipe2_io_pipe_phv_out_data_58; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_59 = pipe2_io_pipe_phv_out_data_59; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_60 = pipe2_io_pipe_phv_out_data_60; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_61 = pipe2_io_pipe_phv_out_data_61; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_62 = pipe2_io_pipe_phv_out_data_62; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_63 = pipe2_io_pipe_phv_out_data_63; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_64 = pipe2_io_pipe_phv_out_data_64; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_65 = pipe2_io_pipe_phv_out_data_65; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_66 = pipe2_io_pipe_phv_out_data_66; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_67 = pipe2_io_pipe_phv_out_data_67; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_68 = pipe2_io_pipe_phv_out_data_68; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_69 = pipe2_io_pipe_phv_out_data_69; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_70 = pipe2_io_pipe_phv_out_data_70; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_71 = pipe2_io_pipe_phv_out_data_71; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_72 = pipe2_io_pipe_phv_out_data_72; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_73 = pipe2_io_pipe_phv_out_data_73; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_74 = pipe2_io_pipe_phv_out_data_74; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_75 = pipe2_io_pipe_phv_out_data_75; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_76 = pipe2_io_pipe_phv_out_data_76; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_77 = pipe2_io_pipe_phv_out_data_77; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_78 = pipe2_io_pipe_phv_out_data_78; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_79 = pipe2_io_pipe_phv_out_data_79; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_80 = pipe2_io_pipe_phv_out_data_80; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_81 = pipe2_io_pipe_phv_out_data_81; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_82 = pipe2_io_pipe_phv_out_data_82; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_83 = pipe2_io_pipe_phv_out_data_83; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_84 = pipe2_io_pipe_phv_out_data_84; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_85 = pipe2_io_pipe_phv_out_data_85; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_86 = pipe2_io_pipe_phv_out_data_86; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_87 = pipe2_io_pipe_phv_out_data_87; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_88 = pipe2_io_pipe_phv_out_data_88; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_89 = pipe2_io_pipe_phv_out_data_89; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_90 = pipe2_io_pipe_phv_out_data_90; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_91 = pipe2_io_pipe_phv_out_data_91; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_92 = pipe2_io_pipe_phv_out_data_92; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_93 = pipe2_io_pipe_phv_out_data_93; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_94 = pipe2_io_pipe_phv_out_data_94; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_95 = pipe2_io_pipe_phv_out_data_95; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_96 = pipe2_io_pipe_phv_out_data_96; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_97 = pipe2_io_pipe_phv_out_data_97; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_98 = pipe2_io_pipe_phv_out_data_98; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_99 = pipe2_io_pipe_phv_out_data_99; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_100 = pipe2_io_pipe_phv_out_data_100; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_101 = pipe2_io_pipe_phv_out_data_101; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_102 = pipe2_io_pipe_phv_out_data_102; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_103 = pipe2_io_pipe_phv_out_data_103; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_104 = pipe2_io_pipe_phv_out_data_104; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_105 = pipe2_io_pipe_phv_out_data_105; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_106 = pipe2_io_pipe_phv_out_data_106; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_107 = pipe2_io_pipe_phv_out_data_107; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_108 = pipe2_io_pipe_phv_out_data_108; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_109 = pipe2_io_pipe_phv_out_data_109; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_110 = pipe2_io_pipe_phv_out_data_110; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_111 = pipe2_io_pipe_phv_out_data_111; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_112 = pipe2_io_pipe_phv_out_data_112; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_113 = pipe2_io_pipe_phv_out_data_113; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_114 = pipe2_io_pipe_phv_out_data_114; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_115 = pipe2_io_pipe_phv_out_data_115; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_116 = pipe2_io_pipe_phv_out_data_116; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_117 = pipe2_io_pipe_phv_out_data_117; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_118 = pipe2_io_pipe_phv_out_data_118; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_119 = pipe2_io_pipe_phv_out_data_119; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_120 = pipe2_io_pipe_phv_out_data_120; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_121 = pipe2_io_pipe_phv_out_data_121; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_122 = pipe2_io_pipe_phv_out_data_122; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_123 = pipe2_io_pipe_phv_out_data_123; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_124 = pipe2_io_pipe_phv_out_data_124; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_125 = pipe2_io_pipe_phv_out_data_125; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_126 = pipe2_io_pipe_phv_out_data_126; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_127 = pipe2_io_pipe_phv_out_data_127; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_128 = pipe2_io_pipe_phv_out_data_128; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_129 = pipe2_io_pipe_phv_out_data_129; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_130 = pipe2_io_pipe_phv_out_data_130; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_131 = pipe2_io_pipe_phv_out_data_131; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_132 = pipe2_io_pipe_phv_out_data_132; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_133 = pipe2_io_pipe_phv_out_data_133; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_134 = pipe2_io_pipe_phv_out_data_134; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_135 = pipe2_io_pipe_phv_out_data_135; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_136 = pipe2_io_pipe_phv_out_data_136; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_137 = pipe2_io_pipe_phv_out_data_137; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_138 = pipe2_io_pipe_phv_out_data_138; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_139 = pipe2_io_pipe_phv_out_data_139; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_140 = pipe2_io_pipe_phv_out_data_140; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_141 = pipe2_io_pipe_phv_out_data_141; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_142 = pipe2_io_pipe_phv_out_data_142; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_143 = pipe2_io_pipe_phv_out_data_143; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_144 = pipe2_io_pipe_phv_out_data_144; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_145 = pipe2_io_pipe_phv_out_data_145; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_146 = pipe2_io_pipe_phv_out_data_146; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_147 = pipe2_io_pipe_phv_out_data_147; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_148 = pipe2_io_pipe_phv_out_data_148; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_149 = pipe2_io_pipe_phv_out_data_149; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_150 = pipe2_io_pipe_phv_out_data_150; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_151 = pipe2_io_pipe_phv_out_data_151; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_152 = pipe2_io_pipe_phv_out_data_152; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_153 = pipe2_io_pipe_phv_out_data_153; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_154 = pipe2_io_pipe_phv_out_data_154; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_155 = pipe2_io_pipe_phv_out_data_155; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_156 = pipe2_io_pipe_phv_out_data_156; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_157 = pipe2_io_pipe_phv_out_data_157; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_158 = pipe2_io_pipe_phv_out_data_158; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_159 = pipe2_io_pipe_phv_out_data_159; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_160 = pipe2_io_pipe_phv_out_data_160; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_161 = pipe2_io_pipe_phv_out_data_161; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_162 = pipe2_io_pipe_phv_out_data_162; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_163 = pipe2_io_pipe_phv_out_data_163; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_164 = pipe2_io_pipe_phv_out_data_164; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_165 = pipe2_io_pipe_phv_out_data_165; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_166 = pipe2_io_pipe_phv_out_data_166; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_167 = pipe2_io_pipe_phv_out_data_167; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_168 = pipe2_io_pipe_phv_out_data_168; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_169 = pipe2_io_pipe_phv_out_data_169; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_170 = pipe2_io_pipe_phv_out_data_170; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_171 = pipe2_io_pipe_phv_out_data_171; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_172 = pipe2_io_pipe_phv_out_data_172; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_173 = pipe2_io_pipe_phv_out_data_173; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_174 = pipe2_io_pipe_phv_out_data_174; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_175 = pipe2_io_pipe_phv_out_data_175; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_176 = pipe2_io_pipe_phv_out_data_176; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_177 = pipe2_io_pipe_phv_out_data_177; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_178 = pipe2_io_pipe_phv_out_data_178; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_179 = pipe2_io_pipe_phv_out_data_179; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_180 = pipe2_io_pipe_phv_out_data_180; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_181 = pipe2_io_pipe_phv_out_data_181; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_182 = pipe2_io_pipe_phv_out_data_182; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_183 = pipe2_io_pipe_phv_out_data_183; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_184 = pipe2_io_pipe_phv_out_data_184; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_185 = pipe2_io_pipe_phv_out_data_185; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_186 = pipe2_io_pipe_phv_out_data_186; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_187 = pipe2_io_pipe_phv_out_data_187; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_188 = pipe2_io_pipe_phv_out_data_188; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_189 = pipe2_io_pipe_phv_out_data_189; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_190 = pipe2_io_pipe_phv_out_data_190; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_191 = pipe2_io_pipe_phv_out_data_191; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_192 = pipe2_io_pipe_phv_out_data_192; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_193 = pipe2_io_pipe_phv_out_data_193; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_194 = pipe2_io_pipe_phv_out_data_194; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_195 = pipe2_io_pipe_phv_out_data_195; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_196 = pipe2_io_pipe_phv_out_data_196; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_197 = pipe2_io_pipe_phv_out_data_197; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_198 = pipe2_io_pipe_phv_out_data_198; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_199 = pipe2_io_pipe_phv_out_data_199; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_200 = pipe2_io_pipe_phv_out_data_200; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_201 = pipe2_io_pipe_phv_out_data_201; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_202 = pipe2_io_pipe_phv_out_data_202; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_203 = pipe2_io_pipe_phv_out_data_203; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_204 = pipe2_io_pipe_phv_out_data_204; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_205 = pipe2_io_pipe_phv_out_data_205; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_206 = pipe2_io_pipe_phv_out_data_206; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_207 = pipe2_io_pipe_phv_out_data_207; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_208 = pipe2_io_pipe_phv_out_data_208; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_209 = pipe2_io_pipe_phv_out_data_209; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_210 = pipe2_io_pipe_phv_out_data_210; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_211 = pipe2_io_pipe_phv_out_data_211; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_212 = pipe2_io_pipe_phv_out_data_212; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_213 = pipe2_io_pipe_phv_out_data_213; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_214 = pipe2_io_pipe_phv_out_data_214; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_215 = pipe2_io_pipe_phv_out_data_215; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_216 = pipe2_io_pipe_phv_out_data_216; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_217 = pipe2_io_pipe_phv_out_data_217; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_218 = pipe2_io_pipe_phv_out_data_218; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_219 = pipe2_io_pipe_phv_out_data_219; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_220 = pipe2_io_pipe_phv_out_data_220; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_221 = pipe2_io_pipe_phv_out_data_221; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_222 = pipe2_io_pipe_phv_out_data_222; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_223 = pipe2_io_pipe_phv_out_data_223; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_224 = pipe2_io_pipe_phv_out_data_224; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_225 = pipe2_io_pipe_phv_out_data_225; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_226 = pipe2_io_pipe_phv_out_data_226; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_227 = pipe2_io_pipe_phv_out_data_227; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_228 = pipe2_io_pipe_phv_out_data_228; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_229 = pipe2_io_pipe_phv_out_data_229; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_230 = pipe2_io_pipe_phv_out_data_230; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_231 = pipe2_io_pipe_phv_out_data_231; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_232 = pipe2_io_pipe_phv_out_data_232; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_233 = pipe2_io_pipe_phv_out_data_233; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_234 = pipe2_io_pipe_phv_out_data_234; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_235 = pipe2_io_pipe_phv_out_data_235; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_236 = pipe2_io_pipe_phv_out_data_236; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_237 = pipe2_io_pipe_phv_out_data_237; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_238 = pipe2_io_pipe_phv_out_data_238; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_239 = pipe2_io_pipe_phv_out_data_239; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_240 = pipe2_io_pipe_phv_out_data_240; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_241 = pipe2_io_pipe_phv_out_data_241; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_242 = pipe2_io_pipe_phv_out_data_242; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_243 = pipe2_io_pipe_phv_out_data_243; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_244 = pipe2_io_pipe_phv_out_data_244; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_245 = pipe2_io_pipe_phv_out_data_245; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_246 = pipe2_io_pipe_phv_out_data_246; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_247 = pipe2_io_pipe_phv_out_data_247; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_248 = pipe2_io_pipe_phv_out_data_248; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_249 = pipe2_io_pipe_phv_out_data_249; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_250 = pipe2_io_pipe_phv_out_data_250; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_251 = pipe2_io_pipe_phv_out_data_251; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_252 = pipe2_io_pipe_phv_out_data_252; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_253 = pipe2_io_pipe_phv_out_data_253; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_254 = pipe2_io_pipe_phv_out_data_254; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_255 = pipe2_io_pipe_phv_out_data_255; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_0 = pipe2_io_pipe_phv_out_header_0; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_1 = pipe2_io_pipe_phv_out_header_1; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_2 = pipe2_io_pipe_phv_out_header_2; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_3 = pipe2_io_pipe_phv_out_header_3; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_4 = pipe2_io_pipe_phv_out_header_4; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_5 = pipe2_io_pipe_phv_out_header_5; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_6 = pipe2_io_pipe_phv_out_header_6; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_7 = pipe2_io_pipe_phv_out_header_7; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_8 = pipe2_io_pipe_phv_out_header_8; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_9 = pipe2_io_pipe_phv_out_header_9; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_10 = pipe2_io_pipe_phv_out_header_10; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_11 = pipe2_io_pipe_phv_out_header_11; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_12 = pipe2_io_pipe_phv_out_header_12; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_13 = pipe2_io_pipe_phv_out_header_13; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_14 = pipe2_io_pipe_phv_out_header_14; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_15 = pipe2_io_pipe_phv_out_header_15; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_parse_current_state = pipe2_io_pipe_phv_out_parse_current_state; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_parse_current_offset = pipe2_io_pipe_phv_out_parse_current_offset; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_parse_transition_field = pipe2_io_pipe_phv_out_parse_transition_field; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_next_processor_id = pipe2_io_pipe_phv_out_next_processor_id; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_next_config_id = pipe2_io_pipe_phv_out_next_config_id; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_is_valid_processor = pipe2_io_pipe_phv_out_is_valid_processor; // @[hash.scala 144:27]
  assign pipe3_io_key_in = pipe2_io_key_out; // @[hash.scala 145:27]
  assign pipe3_io_sum_in = pipe2_io_sum_out; // @[hash.scala 146:27]
  assign pipe4_clock = clock;
  assign pipe4_io_pipe_phv_in_data_0 = pipe3_io_pipe_phv_out_data_0; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_1 = pipe3_io_pipe_phv_out_data_1; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_2 = pipe3_io_pipe_phv_out_data_2; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_3 = pipe3_io_pipe_phv_out_data_3; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_4 = pipe3_io_pipe_phv_out_data_4; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_5 = pipe3_io_pipe_phv_out_data_5; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_6 = pipe3_io_pipe_phv_out_data_6; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_7 = pipe3_io_pipe_phv_out_data_7; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_8 = pipe3_io_pipe_phv_out_data_8; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_9 = pipe3_io_pipe_phv_out_data_9; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_10 = pipe3_io_pipe_phv_out_data_10; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_11 = pipe3_io_pipe_phv_out_data_11; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_12 = pipe3_io_pipe_phv_out_data_12; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_13 = pipe3_io_pipe_phv_out_data_13; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_14 = pipe3_io_pipe_phv_out_data_14; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_15 = pipe3_io_pipe_phv_out_data_15; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_16 = pipe3_io_pipe_phv_out_data_16; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_17 = pipe3_io_pipe_phv_out_data_17; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_18 = pipe3_io_pipe_phv_out_data_18; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_19 = pipe3_io_pipe_phv_out_data_19; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_20 = pipe3_io_pipe_phv_out_data_20; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_21 = pipe3_io_pipe_phv_out_data_21; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_22 = pipe3_io_pipe_phv_out_data_22; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_23 = pipe3_io_pipe_phv_out_data_23; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_24 = pipe3_io_pipe_phv_out_data_24; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_25 = pipe3_io_pipe_phv_out_data_25; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_26 = pipe3_io_pipe_phv_out_data_26; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_27 = pipe3_io_pipe_phv_out_data_27; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_28 = pipe3_io_pipe_phv_out_data_28; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_29 = pipe3_io_pipe_phv_out_data_29; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_30 = pipe3_io_pipe_phv_out_data_30; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_31 = pipe3_io_pipe_phv_out_data_31; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_32 = pipe3_io_pipe_phv_out_data_32; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_33 = pipe3_io_pipe_phv_out_data_33; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_34 = pipe3_io_pipe_phv_out_data_34; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_35 = pipe3_io_pipe_phv_out_data_35; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_36 = pipe3_io_pipe_phv_out_data_36; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_37 = pipe3_io_pipe_phv_out_data_37; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_38 = pipe3_io_pipe_phv_out_data_38; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_39 = pipe3_io_pipe_phv_out_data_39; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_40 = pipe3_io_pipe_phv_out_data_40; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_41 = pipe3_io_pipe_phv_out_data_41; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_42 = pipe3_io_pipe_phv_out_data_42; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_43 = pipe3_io_pipe_phv_out_data_43; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_44 = pipe3_io_pipe_phv_out_data_44; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_45 = pipe3_io_pipe_phv_out_data_45; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_46 = pipe3_io_pipe_phv_out_data_46; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_47 = pipe3_io_pipe_phv_out_data_47; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_48 = pipe3_io_pipe_phv_out_data_48; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_49 = pipe3_io_pipe_phv_out_data_49; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_50 = pipe3_io_pipe_phv_out_data_50; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_51 = pipe3_io_pipe_phv_out_data_51; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_52 = pipe3_io_pipe_phv_out_data_52; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_53 = pipe3_io_pipe_phv_out_data_53; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_54 = pipe3_io_pipe_phv_out_data_54; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_55 = pipe3_io_pipe_phv_out_data_55; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_56 = pipe3_io_pipe_phv_out_data_56; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_57 = pipe3_io_pipe_phv_out_data_57; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_58 = pipe3_io_pipe_phv_out_data_58; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_59 = pipe3_io_pipe_phv_out_data_59; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_60 = pipe3_io_pipe_phv_out_data_60; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_61 = pipe3_io_pipe_phv_out_data_61; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_62 = pipe3_io_pipe_phv_out_data_62; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_63 = pipe3_io_pipe_phv_out_data_63; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_64 = pipe3_io_pipe_phv_out_data_64; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_65 = pipe3_io_pipe_phv_out_data_65; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_66 = pipe3_io_pipe_phv_out_data_66; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_67 = pipe3_io_pipe_phv_out_data_67; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_68 = pipe3_io_pipe_phv_out_data_68; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_69 = pipe3_io_pipe_phv_out_data_69; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_70 = pipe3_io_pipe_phv_out_data_70; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_71 = pipe3_io_pipe_phv_out_data_71; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_72 = pipe3_io_pipe_phv_out_data_72; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_73 = pipe3_io_pipe_phv_out_data_73; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_74 = pipe3_io_pipe_phv_out_data_74; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_75 = pipe3_io_pipe_phv_out_data_75; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_76 = pipe3_io_pipe_phv_out_data_76; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_77 = pipe3_io_pipe_phv_out_data_77; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_78 = pipe3_io_pipe_phv_out_data_78; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_79 = pipe3_io_pipe_phv_out_data_79; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_80 = pipe3_io_pipe_phv_out_data_80; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_81 = pipe3_io_pipe_phv_out_data_81; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_82 = pipe3_io_pipe_phv_out_data_82; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_83 = pipe3_io_pipe_phv_out_data_83; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_84 = pipe3_io_pipe_phv_out_data_84; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_85 = pipe3_io_pipe_phv_out_data_85; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_86 = pipe3_io_pipe_phv_out_data_86; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_87 = pipe3_io_pipe_phv_out_data_87; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_88 = pipe3_io_pipe_phv_out_data_88; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_89 = pipe3_io_pipe_phv_out_data_89; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_90 = pipe3_io_pipe_phv_out_data_90; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_91 = pipe3_io_pipe_phv_out_data_91; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_92 = pipe3_io_pipe_phv_out_data_92; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_93 = pipe3_io_pipe_phv_out_data_93; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_94 = pipe3_io_pipe_phv_out_data_94; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_95 = pipe3_io_pipe_phv_out_data_95; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_96 = pipe3_io_pipe_phv_out_data_96; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_97 = pipe3_io_pipe_phv_out_data_97; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_98 = pipe3_io_pipe_phv_out_data_98; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_99 = pipe3_io_pipe_phv_out_data_99; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_100 = pipe3_io_pipe_phv_out_data_100; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_101 = pipe3_io_pipe_phv_out_data_101; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_102 = pipe3_io_pipe_phv_out_data_102; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_103 = pipe3_io_pipe_phv_out_data_103; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_104 = pipe3_io_pipe_phv_out_data_104; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_105 = pipe3_io_pipe_phv_out_data_105; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_106 = pipe3_io_pipe_phv_out_data_106; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_107 = pipe3_io_pipe_phv_out_data_107; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_108 = pipe3_io_pipe_phv_out_data_108; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_109 = pipe3_io_pipe_phv_out_data_109; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_110 = pipe3_io_pipe_phv_out_data_110; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_111 = pipe3_io_pipe_phv_out_data_111; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_112 = pipe3_io_pipe_phv_out_data_112; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_113 = pipe3_io_pipe_phv_out_data_113; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_114 = pipe3_io_pipe_phv_out_data_114; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_115 = pipe3_io_pipe_phv_out_data_115; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_116 = pipe3_io_pipe_phv_out_data_116; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_117 = pipe3_io_pipe_phv_out_data_117; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_118 = pipe3_io_pipe_phv_out_data_118; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_119 = pipe3_io_pipe_phv_out_data_119; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_120 = pipe3_io_pipe_phv_out_data_120; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_121 = pipe3_io_pipe_phv_out_data_121; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_122 = pipe3_io_pipe_phv_out_data_122; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_123 = pipe3_io_pipe_phv_out_data_123; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_124 = pipe3_io_pipe_phv_out_data_124; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_125 = pipe3_io_pipe_phv_out_data_125; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_126 = pipe3_io_pipe_phv_out_data_126; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_127 = pipe3_io_pipe_phv_out_data_127; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_128 = pipe3_io_pipe_phv_out_data_128; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_129 = pipe3_io_pipe_phv_out_data_129; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_130 = pipe3_io_pipe_phv_out_data_130; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_131 = pipe3_io_pipe_phv_out_data_131; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_132 = pipe3_io_pipe_phv_out_data_132; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_133 = pipe3_io_pipe_phv_out_data_133; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_134 = pipe3_io_pipe_phv_out_data_134; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_135 = pipe3_io_pipe_phv_out_data_135; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_136 = pipe3_io_pipe_phv_out_data_136; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_137 = pipe3_io_pipe_phv_out_data_137; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_138 = pipe3_io_pipe_phv_out_data_138; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_139 = pipe3_io_pipe_phv_out_data_139; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_140 = pipe3_io_pipe_phv_out_data_140; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_141 = pipe3_io_pipe_phv_out_data_141; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_142 = pipe3_io_pipe_phv_out_data_142; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_143 = pipe3_io_pipe_phv_out_data_143; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_144 = pipe3_io_pipe_phv_out_data_144; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_145 = pipe3_io_pipe_phv_out_data_145; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_146 = pipe3_io_pipe_phv_out_data_146; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_147 = pipe3_io_pipe_phv_out_data_147; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_148 = pipe3_io_pipe_phv_out_data_148; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_149 = pipe3_io_pipe_phv_out_data_149; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_150 = pipe3_io_pipe_phv_out_data_150; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_151 = pipe3_io_pipe_phv_out_data_151; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_152 = pipe3_io_pipe_phv_out_data_152; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_153 = pipe3_io_pipe_phv_out_data_153; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_154 = pipe3_io_pipe_phv_out_data_154; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_155 = pipe3_io_pipe_phv_out_data_155; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_156 = pipe3_io_pipe_phv_out_data_156; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_157 = pipe3_io_pipe_phv_out_data_157; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_158 = pipe3_io_pipe_phv_out_data_158; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_159 = pipe3_io_pipe_phv_out_data_159; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_160 = pipe3_io_pipe_phv_out_data_160; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_161 = pipe3_io_pipe_phv_out_data_161; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_162 = pipe3_io_pipe_phv_out_data_162; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_163 = pipe3_io_pipe_phv_out_data_163; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_164 = pipe3_io_pipe_phv_out_data_164; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_165 = pipe3_io_pipe_phv_out_data_165; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_166 = pipe3_io_pipe_phv_out_data_166; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_167 = pipe3_io_pipe_phv_out_data_167; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_168 = pipe3_io_pipe_phv_out_data_168; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_169 = pipe3_io_pipe_phv_out_data_169; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_170 = pipe3_io_pipe_phv_out_data_170; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_171 = pipe3_io_pipe_phv_out_data_171; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_172 = pipe3_io_pipe_phv_out_data_172; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_173 = pipe3_io_pipe_phv_out_data_173; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_174 = pipe3_io_pipe_phv_out_data_174; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_175 = pipe3_io_pipe_phv_out_data_175; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_176 = pipe3_io_pipe_phv_out_data_176; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_177 = pipe3_io_pipe_phv_out_data_177; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_178 = pipe3_io_pipe_phv_out_data_178; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_179 = pipe3_io_pipe_phv_out_data_179; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_180 = pipe3_io_pipe_phv_out_data_180; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_181 = pipe3_io_pipe_phv_out_data_181; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_182 = pipe3_io_pipe_phv_out_data_182; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_183 = pipe3_io_pipe_phv_out_data_183; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_184 = pipe3_io_pipe_phv_out_data_184; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_185 = pipe3_io_pipe_phv_out_data_185; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_186 = pipe3_io_pipe_phv_out_data_186; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_187 = pipe3_io_pipe_phv_out_data_187; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_188 = pipe3_io_pipe_phv_out_data_188; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_189 = pipe3_io_pipe_phv_out_data_189; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_190 = pipe3_io_pipe_phv_out_data_190; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_191 = pipe3_io_pipe_phv_out_data_191; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_192 = pipe3_io_pipe_phv_out_data_192; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_193 = pipe3_io_pipe_phv_out_data_193; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_194 = pipe3_io_pipe_phv_out_data_194; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_195 = pipe3_io_pipe_phv_out_data_195; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_196 = pipe3_io_pipe_phv_out_data_196; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_197 = pipe3_io_pipe_phv_out_data_197; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_198 = pipe3_io_pipe_phv_out_data_198; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_199 = pipe3_io_pipe_phv_out_data_199; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_200 = pipe3_io_pipe_phv_out_data_200; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_201 = pipe3_io_pipe_phv_out_data_201; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_202 = pipe3_io_pipe_phv_out_data_202; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_203 = pipe3_io_pipe_phv_out_data_203; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_204 = pipe3_io_pipe_phv_out_data_204; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_205 = pipe3_io_pipe_phv_out_data_205; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_206 = pipe3_io_pipe_phv_out_data_206; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_207 = pipe3_io_pipe_phv_out_data_207; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_208 = pipe3_io_pipe_phv_out_data_208; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_209 = pipe3_io_pipe_phv_out_data_209; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_210 = pipe3_io_pipe_phv_out_data_210; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_211 = pipe3_io_pipe_phv_out_data_211; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_212 = pipe3_io_pipe_phv_out_data_212; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_213 = pipe3_io_pipe_phv_out_data_213; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_214 = pipe3_io_pipe_phv_out_data_214; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_215 = pipe3_io_pipe_phv_out_data_215; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_216 = pipe3_io_pipe_phv_out_data_216; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_217 = pipe3_io_pipe_phv_out_data_217; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_218 = pipe3_io_pipe_phv_out_data_218; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_219 = pipe3_io_pipe_phv_out_data_219; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_220 = pipe3_io_pipe_phv_out_data_220; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_221 = pipe3_io_pipe_phv_out_data_221; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_222 = pipe3_io_pipe_phv_out_data_222; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_223 = pipe3_io_pipe_phv_out_data_223; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_224 = pipe3_io_pipe_phv_out_data_224; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_225 = pipe3_io_pipe_phv_out_data_225; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_226 = pipe3_io_pipe_phv_out_data_226; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_227 = pipe3_io_pipe_phv_out_data_227; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_228 = pipe3_io_pipe_phv_out_data_228; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_229 = pipe3_io_pipe_phv_out_data_229; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_230 = pipe3_io_pipe_phv_out_data_230; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_231 = pipe3_io_pipe_phv_out_data_231; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_232 = pipe3_io_pipe_phv_out_data_232; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_233 = pipe3_io_pipe_phv_out_data_233; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_234 = pipe3_io_pipe_phv_out_data_234; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_235 = pipe3_io_pipe_phv_out_data_235; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_236 = pipe3_io_pipe_phv_out_data_236; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_237 = pipe3_io_pipe_phv_out_data_237; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_238 = pipe3_io_pipe_phv_out_data_238; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_239 = pipe3_io_pipe_phv_out_data_239; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_240 = pipe3_io_pipe_phv_out_data_240; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_241 = pipe3_io_pipe_phv_out_data_241; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_242 = pipe3_io_pipe_phv_out_data_242; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_243 = pipe3_io_pipe_phv_out_data_243; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_244 = pipe3_io_pipe_phv_out_data_244; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_245 = pipe3_io_pipe_phv_out_data_245; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_246 = pipe3_io_pipe_phv_out_data_246; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_247 = pipe3_io_pipe_phv_out_data_247; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_248 = pipe3_io_pipe_phv_out_data_248; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_249 = pipe3_io_pipe_phv_out_data_249; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_250 = pipe3_io_pipe_phv_out_data_250; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_251 = pipe3_io_pipe_phv_out_data_251; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_252 = pipe3_io_pipe_phv_out_data_252; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_253 = pipe3_io_pipe_phv_out_data_253; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_254 = pipe3_io_pipe_phv_out_data_254; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_255 = pipe3_io_pipe_phv_out_data_255; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_0 = pipe3_io_pipe_phv_out_header_0; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_1 = pipe3_io_pipe_phv_out_header_1; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_2 = pipe3_io_pipe_phv_out_header_2; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_3 = pipe3_io_pipe_phv_out_header_3; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_4 = pipe3_io_pipe_phv_out_header_4; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_5 = pipe3_io_pipe_phv_out_header_5; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_6 = pipe3_io_pipe_phv_out_header_6; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_7 = pipe3_io_pipe_phv_out_header_7; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_8 = pipe3_io_pipe_phv_out_header_8; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_9 = pipe3_io_pipe_phv_out_header_9; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_10 = pipe3_io_pipe_phv_out_header_10; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_11 = pipe3_io_pipe_phv_out_header_11; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_12 = pipe3_io_pipe_phv_out_header_12; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_13 = pipe3_io_pipe_phv_out_header_13; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_14 = pipe3_io_pipe_phv_out_header_14; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_15 = pipe3_io_pipe_phv_out_header_15; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_parse_current_state = pipe3_io_pipe_phv_out_parse_current_state; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_parse_current_offset = pipe3_io_pipe_phv_out_parse_current_offset; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_parse_transition_field = pipe3_io_pipe_phv_out_parse_transition_field; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_next_processor_id = pipe3_io_pipe_phv_out_next_processor_id; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_next_config_id = pipe3_io_pipe_phv_out_next_config_id; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_is_valid_processor = pipe3_io_pipe_phv_out_is_valid_processor; // @[hash.scala 148:27]
  assign pipe4_io_key_in = pipe3_io_key_out; // @[hash.scala 149:27]
  assign pipe4_io_sum_in = pipe3_io_sum_out; // @[hash.scala 150:27]
  assign pipe5_clock = clock;
  assign pipe5_io_pipe_phv_in_data_0 = pipe4_io_pipe_phv_out_data_0; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_1 = pipe4_io_pipe_phv_out_data_1; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_2 = pipe4_io_pipe_phv_out_data_2; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_3 = pipe4_io_pipe_phv_out_data_3; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_4 = pipe4_io_pipe_phv_out_data_4; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_5 = pipe4_io_pipe_phv_out_data_5; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_6 = pipe4_io_pipe_phv_out_data_6; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_7 = pipe4_io_pipe_phv_out_data_7; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_8 = pipe4_io_pipe_phv_out_data_8; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_9 = pipe4_io_pipe_phv_out_data_9; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_10 = pipe4_io_pipe_phv_out_data_10; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_11 = pipe4_io_pipe_phv_out_data_11; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_12 = pipe4_io_pipe_phv_out_data_12; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_13 = pipe4_io_pipe_phv_out_data_13; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_14 = pipe4_io_pipe_phv_out_data_14; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_15 = pipe4_io_pipe_phv_out_data_15; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_16 = pipe4_io_pipe_phv_out_data_16; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_17 = pipe4_io_pipe_phv_out_data_17; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_18 = pipe4_io_pipe_phv_out_data_18; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_19 = pipe4_io_pipe_phv_out_data_19; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_20 = pipe4_io_pipe_phv_out_data_20; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_21 = pipe4_io_pipe_phv_out_data_21; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_22 = pipe4_io_pipe_phv_out_data_22; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_23 = pipe4_io_pipe_phv_out_data_23; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_24 = pipe4_io_pipe_phv_out_data_24; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_25 = pipe4_io_pipe_phv_out_data_25; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_26 = pipe4_io_pipe_phv_out_data_26; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_27 = pipe4_io_pipe_phv_out_data_27; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_28 = pipe4_io_pipe_phv_out_data_28; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_29 = pipe4_io_pipe_phv_out_data_29; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_30 = pipe4_io_pipe_phv_out_data_30; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_31 = pipe4_io_pipe_phv_out_data_31; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_32 = pipe4_io_pipe_phv_out_data_32; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_33 = pipe4_io_pipe_phv_out_data_33; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_34 = pipe4_io_pipe_phv_out_data_34; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_35 = pipe4_io_pipe_phv_out_data_35; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_36 = pipe4_io_pipe_phv_out_data_36; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_37 = pipe4_io_pipe_phv_out_data_37; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_38 = pipe4_io_pipe_phv_out_data_38; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_39 = pipe4_io_pipe_phv_out_data_39; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_40 = pipe4_io_pipe_phv_out_data_40; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_41 = pipe4_io_pipe_phv_out_data_41; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_42 = pipe4_io_pipe_phv_out_data_42; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_43 = pipe4_io_pipe_phv_out_data_43; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_44 = pipe4_io_pipe_phv_out_data_44; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_45 = pipe4_io_pipe_phv_out_data_45; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_46 = pipe4_io_pipe_phv_out_data_46; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_47 = pipe4_io_pipe_phv_out_data_47; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_48 = pipe4_io_pipe_phv_out_data_48; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_49 = pipe4_io_pipe_phv_out_data_49; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_50 = pipe4_io_pipe_phv_out_data_50; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_51 = pipe4_io_pipe_phv_out_data_51; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_52 = pipe4_io_pipe_phv_out_data_52; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_53 = pipe4_io_pipe_phv_out_data_53; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_54 = pipe4_io_pipe_phv_out_data_54; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_55 = pipe4_io_pipe_phv_out_data_55; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_56 = pipe4_io_pipe_phv_out_data_56; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_57 = pipe4_io_pipe_phv_out_data_57; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_58 = pipe4_io_pipe_phv_out_data_58; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_59 = pipe4_io_pipe_phv_out_data_59; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_60 = pipe4_io_pipe_phv_out_data_60; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_61 = pipe4_io_pipe_phv_out_data_61; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_62 = pipe4_io_pipe_phv_out_data_62; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_63 = pipe4_io_pipe_phv_out_data_63; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_64 = pipe4_io_pipe_phv_out_data_64; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_65 = pipe4_io_pipe_phv_out_data_65; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_66 = pipe4_io_pipe_phv_out_data_66; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_67 = pipe4_io_pipe_phv_out_data_67; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_68 = pipe4_io_pipe_phv_out_data_68; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_69 = pipe4_io_pipe_phv_out_data_69; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_70 = pipe4_io_pipe_phv_out_data_70; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_71 = pipe4_io_pipe_phv_out_data_71; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_72 = pipe4_io_pipe_phv_out_data_72; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_73 = pipe4_io_pipe_phv_out_data_73; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_74 = pipe4_io_pipe_phv_out_data_74; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_75 = pipe4_io_pipe_phv_out_data_75; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_76 = pipe4_io_pipe_phv_out_data_76; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_77 = pipe4_io_pipe_phv_out_data_77; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_78 = pipe4_io_pipe_phv_out_data_78; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_79 = pipe4_io_pipe_phv_out_data_79; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_80 = pipe4_io_pipe_phv_out_data_80; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_81 = pipe4_io_pipe_phv_out_data_81; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_82 = pipe4_io_pipe_phv_out_data_82; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_83 = pipe4_io_pipe_phv_out_data_83; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_84 = pipe4_io_pipe_phv_out_data_84; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_85 = pipe4_io_pipe_phv_out_data_85; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_86 = pipe4_io_pipe_phv_out_data_86; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_87 = pipe4_io_pipe_phv_out_data_87; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_88 = pipe4_io_pipe_phv_out_data_88; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_89 = pipe4_io_pipe_phv_out_data_89; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_90 = pipe4_io_pipe_phv_out_data_90; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_91 = pipe4_io_pipe_phv_out_data_91; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_92 = pipe4_io_pipe_phv_out_data_92; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_93 = pipe4_io_pipe_phv_out_data_93; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_94 = pipe4_io_pipe_phv_out_data_94; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_95 = pipe4_io_pipe_phv_out_data_95; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_96 = pipe4_io_pipe_phv_out_data_96; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_97 = pipe4_io_pipe_phv_out_data_97; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_98 = pipe4_io_pipe_phv_out_data_98; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_99 = pipe4_io_pipe_phv_out_data_99; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_100 = pipe4_io_pipe_phv_out_data_100; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_101 = pipe4_io_pipe_phv_out_data_101; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_102 = pipe4_io_pipe_phv_out_data_102; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_103 = pipe4_io_pipe_phv_out_data_103; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_104 = pipe4_io_pipe_phv_out_data_104; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_105 = pipe4_io_pipe_phv_out_data_105; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_106 = pipe4_io_pipe_phv_out_data_106; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_107 = pipe4_io_pipe_phv_out_data_107; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_108 = pipe4_io_pipe_phv_out_data_108; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_109 = pipe4_io_pipe_phv_out_data_109; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_110 = pipe4_io_pipe_phv_out_data_110; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_111 = pipe4_io_pipe_phv_out_data_111; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_112 = pipe4_io_pipe_phv_out_data_112; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_113 = pipe4_io_pipe_phv_out_data_113; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_114 = pipe4_io_pipe_phv_out_data_114; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_115 = pipe4_io_pipe_phv_out_data_115; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_116 = pipe4_io_pipe_phv_out_data_116; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_117 = pipe4_io_pipe_phv_out_data_117; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_118 = pipe4_io_pipe_phv_out_data_118; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_119 = pipe4_io_pipe_phv_out_data_119; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_120 = pipe4_io_pipe_phv_out_data_120; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_121 = pipe4_io_pipe_phv_out_data_121; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_122 = pipe4_io_pipe_phv_out_data_122; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_123 = pipe4_io_pipe_phv_out_data_123; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_124 = pipe4_io_pipe_phv_out_data_124; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_125 = pipe4_io_pipe_phv_out_data_125; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_126 = pipe4_io_pipe_phv_out_data_126; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_127 = pipe4_io_pipe_phv_out_data_127; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_128 = pipe4_io_pipe_phv_out_data_128; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_129 = pipe4_io_pipe_phv_out_data_129; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_130 = pipe4_io_pipe_phv_out_data_130; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_131 = pipe4_io_pipe_phv_out_data_131; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_132 = pipe4_io_pipe_phv_out_data_132; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_133 = pipe4_io_pipe_phv_out_data_133; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_134 = pipe4_io_pipe_phv_out_data_134; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_135 = pipe4_io_pipe_phv_out_data_135; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_136 = pipe4_io_pipe_phv_out_data_136; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_137 = pipe4_io_pipe_phv_out_data_137; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_138 = pipe4_io_pipe_phv_out_data_138; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_139 = pipe4_io_pipe_phv_out_data_139; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_140 = pipe4_io_pipe_phv_out_data_140; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_141 = pipe4_io_pipe_phv_out_data_141; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_142 = pipe4_io_pipe_phv_out_data_142; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_143 = pipe4_io_pipe_phv_out_data_143; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_144 = pipe4_io_pipe_phv_out_data_144; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_145 = pipe4_io_pipe_phv_out_data_145; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_146 = pipe4_io_pipe_phv_out_data_146; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_147 = pipe4_io_pipe_phv_out_data_147; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_148 = pipe4_io_pipe_phv_out_data_148; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_149 = pipe4_io_pipe_phv_out_data_149; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_150 = pipe4_io_pipe_phv_out_data_150; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_151 = pipe4_io_pipe_phv_out_data_151; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_152 = pipe4_io_pipe_phv_out_data_152; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_153 = pipe4_io_pipe_phv_out_data_153; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_154 = pipe4_io_pipe_phv_out_data_154; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_155 = pipe4_io_pipe_phv_out_data_155; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_156 = pipe4_io_pipe_phv_out_data_156; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_157 = pipe4_io_pipe_phv_out_data_157; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_158 = pipe4_io_pipe_phv_out_data_158; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_159 = pipe4_io_pipe_phv_out_data_159; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_160 = pipe4_io_pipe_phv_out_data_160; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_161 = pipe4_io_pipe_phv_out_data_161; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_162 = pipe4_io_pipe_phv_out_data_162; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_163 = pipe4_io_pipe_phv_out_data_163; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_164 = pipe4_io_pipe_phv_out_data_164; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_165 = pipe4_io_pipe_phv_out_data_165; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_166 = pipe4_io_pipe_phv_out_data_166; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_167 = pipe4_io_pipe_phv_out_data_167; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_168 = pipe4_io_pipe_phv_out_data_168; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_169 = pipe4_io_pipe_phv_out_data_169; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_170 = pipe4_io_pipe_phv_out_data_170; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_171 = pipe4_io_pipe_phv_out_data_171; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_172 = pipe4_io_pipe_phv_out_data_172; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_173 = pipe4_io_pipe_phv_out_data_173; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_174 = pipe4_io_pipe_phv_out_data_174; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_175 = pipe4_io_pipe_phv_out_data_175; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_176 = pipe4_io_pipe_phv_out_data_176; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_177 = pipe4_io_pipe_phv_out_data_177; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_178 = pipe4_io_pipe_phv_out_data_178; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_179 = pipe4_io_pipe_phv_out_data_179; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_180 = pipe4_io_pipe_phv_out_data_180; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_181 = pipe4_io_pipe_phv_out_data_181; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_182 = pipe4_io_pipe_phv_out_data_182; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_183 = pipe4_io_pipe_phv_out_data_183; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_184 = pipe4_io_pipe_phv_out_data_184; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_185 = pipe4_io_pipe_phv_out_data_185; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_186 = pipe4_io_pipe_phv_out_data_186; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_187 = pipe4_io_pipe_phv_out_data_187; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_188 = pipe4_io_pipe_phv_out_data_188; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_189 = pipe4_io_pipe_phv_out_data_189; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_190 = pipe4_io_pipe_phv_out_data_190; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_191 = pipe4_io_pipe_phv_out_data_191; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_192 = pipe4_io_pipe_phv_out_data_192; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_193 = pipe4_io_pipe_phv_out_data_193; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_194 = pipe4_io_pipe_phv_out_data_194; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_195 = pipe4_io_pipe_phv_out_data_195; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_196 = pipe4_io_pipe_phv_out_data_196; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_197 = pipe4_io_pipe_phv_out_data_197; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_198 = pipe4_io_pipe_phv_out_data_198; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_199 = pipe4_io_pipe_phv_out_data_199; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_200 = pipe4_io_pipe_phv_out_data_200; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_201 = pipe4_io_pipe_phv_out_data_201; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_202 = pipe4_io_pipe_phv_out_data_202; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_203 = pipe4_io_pipe_phv_out_data_203; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_204 = pipe4_io_pipe_phv_out_data_204; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_205 = pipe4_io_pipe_phv_out_data_205; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_206 = pipe4_io_pipe_phv_out_data_206; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_207 = pipe4_io_pipe_phv_out_data_207; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_208 = pipe4_io_pipe_phv_out_data_208; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_209 = pipe4_io_pipe_phv_out_data_209; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_210 = pipe4_io_pipe_phv_out_data_210; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_211 = pipe4_io_pipe_phv_out_data_211; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_212 = pipe4_io_pipe_phv_out_data_212; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_213 = pipe4_io_pipe_phv_out_data_213; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_214 = pipe4_io_pipe_phv_out_data_214; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_215 = pipe4_io_pipe_phv_out_data_215; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_216 = pipe4_io_pipe_phv_out_data_216; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_217 = pipe4_io_pipe_phv_out_data_217; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_218 = pipe4_io_pipe_phv_out_data_218; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_219 = pipe4_io_pipe_phv_out_data_219; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_220 = pipe4_io_pipe_phv_out_data_220; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_221 = pipe4_io_pipe_phv_out_data_221; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_222 = pipe4_io_pipe_phv_out_data_222; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_223 = pipe4_io_pipe_phv_out_data_223; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_224 = pipe4_io_pipe_phv_out_data_224; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_225 = pipe4_io_pipe_phv_out_data_225; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_226 = pipe4_io_pipe_phv_out_data_226; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_227 = pipe4_io_pipe_phv_out_data_227; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_228 = pipe4_io_pipe_phv_out_data_228; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_229 = pipe4_io_pipe_phv_out_data_229; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_230 = pipe4_io_pipe_phv_out_data_230; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_231 = pipe4_io_pipe_phv_out_data_231; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_232 = pipe4_io_pipe_phv_out_data_232; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_233 = pipe4_io_pipe_phv_out_data_233; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_234 = pipe4_io_pipe_phv_out_data_234; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_235 = pipe4_io_pipe_phv_out_data_235; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_236 = pipe4_io_pipe_phv_out_data_236; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_237 = pipe4_io_pipe_phv_out_data_237; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_238 = pipe4_io_pipe_phv_out_data_238; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_239 = pipe4_io_pipe_phv_out_data_239; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_240 = pipe4_io_pipe_phv_out_data_240; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_241 = pipe4_io_pipe_phv_out_data_241; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_242 = pipe4_io_pipe_phv_out_data_242; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_243 = pipe4_io_pipe_phv_out_data_243; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_244 = pipe4_io_pipe_phv_out_data_244; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_245 = pipe4_io_pipe_phv_out_data_245; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_246 = pipe4_io_pipe_phv_out_data_246; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_247 = pipe4_io_pipe_phv_out_data_247; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_248 = pipe4_io_pipe_phv_out_data_248; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_249 = pipe4_io_pipe_phv_out_data_249; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_250 = pipe4_io_pipe_phv_out_data_250; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_251 = pipe4_io_pipe_phv_out_data_251; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_252 = pipe4_io_pipe_phv_out_data_252; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_253 = pipe4_io_pipe_phv_out_data_253; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_254 = pipe4_io_pipe_phv_out_data_254; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_255 = pipe4_io_pipe_phv_out_data_255; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_0 = pipe4_io_pipe_phv_out_header_0; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_1 = pipe4_io_pipe_phv_out_header_1; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_2 = pipe4_io_pipe_phv_out_header_2; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_3 = pipe4_io_pipe_phv_out_header_3; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_4 = pipe4_io_pipe_phv_out_header_4; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_5 = pipe4_io_pipe_phv_out_header_5; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_6 = pipe4_io_pipe_phv_out_header_6; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_7 = pipe4_io_pipe_phv_out_header_7; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_8 = pipe4_io_pipe_phv_out_header_8; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_9 = pipe4_io_pipe_phv_out_header_9; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_10 = pipe4_io_pipe_phv_out_header_10; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_11 = pipe4_io_pipe_phv_out_header_11; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_12 = pipe4_io_pipe_phv_out_header_12; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_13 = pipe4_io_pipe_phv_out_header_13; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_14 = pipe4_io_pipe_phv_out_header_14; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_15 = pipe4_io_pipe_phv_out_header_15; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_parse_current_state = pipe4_io_pipe_phv_out_parse_current_state; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_parse_current_offset = pipe4_io_pipe_phv_out_parse_current_offset; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_parse_transition_field = pipe4_io_pipe_phv_out_parse_transition_field; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_next_processor_id = pipe4_io_pipe_phv_out_next_processor_id; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_next_config_id = pipe4_io_pipe_phv_out_next_config_id; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_is_valid_processor = pipe4_io_pipe_phv_out_is_valid_processor; // @[hash.scala 152:27]
  assign pipe5_io_hash_depth_0 = hash_depth_0; // @[hash.scala 156:27]
  assign pipe5_io_hash_depth_1 = hash_depth_1; // @[hash.scala 156:27]
  assign pipe5_io_key_in = pipe4_io_key_out; // @[hash.scala 153:27]
  assign pipe5_io_sum_in = pipe4_io_sum_out[15:0]; // @[hash.scala 154:27]
  assign pipe6_clock = clock;
  assign pipe6_io_pipe_phv_in_data_0 = pipe5_io_pipe_phv_out_data_0; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_1 = pipe5_io_pipe_phv_out_data_1; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_2 = pipe5_io_pipe_phv_out_data_2; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_3 = pipe5_io_pipe_phv_out_data_3; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_4 = pipe5_io_pipe_phv_out_data_4; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_5 = pipe5_io_pipe_phv_out_data_5; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_6 = pipe5_io_pipe_phv_out_data_6; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_7 = pipe5_io_pipe_phv_out_data_7; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_8 = pipe5_io_pipe_phv_out_data_8; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_9 = pipe5_io_pipe_phv_out_data_9; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_10 = pipe5_io_pipe_phv_out_data_10; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_11 = pipe5_io_pipe_phv_out_data_11; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_12 = pipe5_io_pipe_phv_out_data_12; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_13 = pipe5_io_pipe_phv_out_data_13; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_14 = pipe5_io_pipe_phv_out_data_14; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_15 = pipe5_io_pipe_phv_out_data_15; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_16 = pipe5_io_pipe_phv_out_data_16; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_17 = pipe5_io_pipe_phv_out_data_17; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_18 = pipe5_io_pipe_phv_out_data_18; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_19 = pipe5_io_pipe_phv_out_data_19; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_20 = pipe5_io_pipe_phv_out_data_20; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_21 = pipe5_io_pipe_phv_out_data_21; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_22 = pipe5_io_pipe_phv_out_data_22; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_23 = pipe5_io_pipe_phv_out_data_23; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_24 = pipe5_io_pipe_phv_out_data_24; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_25 = pipe5_io_pipe_phv_out_data_25; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_26 = pipe5_io_pipe_phv_out_data_26; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_27 = pipe5_io_pipe_phv_out_data_27; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_28 = pipe5_io_pipe_phv_out_data_28; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_29 = pipe5_io_pipe_phv_out_data_29; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_30 = pipe5_io_pipe_phv_out_data_30; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_31 = pipe5_io_pipe_phv_out_data_31; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_32 = pipe5_io_pipe_phv_out_data_32; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_33 = pipe5_io_pipe_phv_out_data_33; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_34 = pipe5_io_pipe_phv_out_data_34; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_35 = pipe5_io_pipe_phv_out_data_35; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_36 = pipe5_io_pipe_phv_out_data_36; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_37 = pipe5_io_pipe_phv_out_data_37; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_38 = pipe5_io_pipe_phv_out_data_38; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_39 = pipe5_io_pipe_phv_out_data_39; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_40 = pipe5_io_pipe_phv_out_data_40; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_41 = pipe5_io_pipe_phv_out_data_41; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_42 = pipe5_io_pipe_phv_out_data_42; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_43 = pipe5_io_pipe_phv_out_data_43; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_44 = pipe5_io_pipe_phv_out_data_44; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_45 = pipe5_io_pipe_phv_out_data_45; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_46 = pipe5_io_pipe_phv_out_data_46; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_47 = pipe5_io_pipe_phv_out_data_47; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_48 = pipe5_io_pipe_phv_out_data_48; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_49 = pipe5_io_pipe_phv_out_data_49; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_50 = pipe5_io_pipe_phv_out_data_50; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_51 = pipe5_io_pipe_phv_out_data_51; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_52 = pipe5_io_pipe_phv_out_data_52; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_53 = pipe5_io_pipe_phv_out_data_53; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_54 = pipe5_io_pipe_phv_out_data_54; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_55 = pipe5_io_pipe_phv_out_data_55; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_56 = pipe5_io_pipe_phv_out_data_56; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_57 = pipe5_io_pipe_phv_out_data_57; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_58 = pipe5_io_pipe_phv_out_data_58; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_59 = pipe5_io_pipe_phv_out_data_59; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_60 = pipe5_io_pipe_phv_out_data_60; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_61 = pipe5_io_pipe_phv_out_data_61; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_62 = pipe5_io_pipe_phv_out_data_62; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_63 = pipe5_io_pipe_phv_out_data_63; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_64 = pipe5_io_pipe_phv_out_data_64; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_65 = pipe5_io_pipe_phv_out_data_65; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_66 = pipe5_io_pipe_phv_out_data_66; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_67 = pipe5_io_pipe_phv_out_data_67; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_68 = pipe5_io_pipe_phv_out_data_68; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_69 = pipe5_io_pipe_phv_out_data_69; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_70 = pipe5_io_pipe_phv_out_data_70; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_71 = pipe5_io_pipe_phv_out_data_71; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_72 = pipe5_io_pipe_phv_out_data_72; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_73 = pipe5_io_pipe_phv_out_data_73; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_74 = pipe5_io_pipe_phv_out_data_74; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_75 = pipe5_io_pipe_phv_out_data_75; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_76 = pipe5_io_pipe_phv_out_data_76; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_77 = pipe5_io_pipe_phv_out_data_77; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_78 = pipe5_io_pipe_phv_out_data_78; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_79 = pipe5_io_pipe_phv_out_data_79; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_80 = pipe5_io_pipe_phv_out_data_80; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_81 = pipe5_io_pipe_phv_out_data_81; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_82 = pipe5_io_pipe_phv_out_data_82; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_83 = pipe5_io_pipe_phv_out_data_83; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_84 = pipe5_io_pipe_phv_out_data_84; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_85 = pipe5_io_pipe_phv_out_data_85; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_86 = pipe5_io_pipe_phv_out_data_86; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_87 = pipe5_io_pipe_phv_out_data_87; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_88 = pipe5_io_pipe_phv_out_data_88; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_89 = pipe5_io_pipe_phv_out_data_89; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_90 = pipe5_io_pipe_phv_out_data_90; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_91 = pipe5_io_pipe_phv_out_data_91; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_92 = pipe5_io_pipe_phv_out_data_92; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_93 = pipe5_io_pipe_phv_out_data_93; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_94 = pipe5_io_pipe_phv_out_data_94; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_95 = pipe5_io_pipe_phv_out_data_95; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_96 = pipe5_io_pipe_phv_out_data_96; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_97 = pipe5_io_pipe_phv_out_data_97; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_98 = pipe5_io_pipe_phv_out_data_98; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_99 = pipe5_io_pipe_phv_out_data_99; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_100 = pipe5_io_pipe_phv_out_data_100; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_101 = pipe5_io_pipe_phv_out_data_101; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_102 = pipe5_io_pipe_phv_out_data_102; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_103 = pipe5_io_pipe_phv_out_data_103; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_104 = pipe5_io_pipe_phv_out_data_104; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_105 = pipe5_io_pipe_phv_out_data_105; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_106 = pipe5_io_pipe_phv_out_data_106; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_107 = pipe5_io_pipe_phv_out_data_107; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_108 = pipe5_io_pipe_phv_out_data_108; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_109 = pipe5_io_pipe_phv_out_data_109; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_110 = pipe5_io_pipe_phv_out_data_110; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_111 = pipe5_io_pipe_phv_out_data_111; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_112 = pipe5_io_pipe_phv_out_data_112; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_113 = pipe5_io_pipe_phv_out_data_113; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_114 = pipe5_io_pipe_phv_out_data_114; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_115 = pipe5_io_pipe_phv_out_data_115; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_116 = pipe5_io_pipe_phv_out_data_116; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_117 = pipe5_io_pipe_phv_out_data_117; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_118 = pipe5_io_pipe_phv_out_data_118; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_119 = pipe5_io_pipe_phv_out_data_119; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_120 = pipe5_io_pipe_phv_out_data_120; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_121 = pipe5_io_pipe_phv_out_data_121; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_122 = pipe5_io_pipe_phv_out_data_122; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_123 = pipe5_io_pipe_phv_out_data_123; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_124 = pipe5_io_pipe_phv_out_data_124; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_125 = pipe5_io_pipe_phv_out_data_125; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_126 = pipe5_io_pipe_phv_out_data_126; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_127 = pipe5_io_pipe_phv_out_data_127; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_128 = pipe5_io_pipe_phv_out_data_128; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_129 = pipe5_io_pipe_phv_out_data_129; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_130 = pipe5_io_pipe_phv_out_data_130; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_131 = pipe5_io_pipe_phv_out_data_131; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_132 = pipe5_io_pipe_phv_out_data_132; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_133 = pipe5_io_pipe_phv_out_data_133; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_134 = pipe5_io_pipe_phv_out_data_134; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_135 = pipe5_io_pipe_phv_out_data_135; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_136 = pipe5_io_pipe_phv_out_data_136; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_137 = pipe5_io_pipe_phv_out_data_137; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_138 = pipe5_io_pipe_phv_out_data_138; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_139 = pipe5_io_pipe_phv_out_data_139; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_140 = pipe5_io_pipe_phv_out_data_140; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_141 = pipe5_io_pipe_phv_out_data_141; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_142 = pipe5_io_pipe_phv_out_data_142; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_143 = pipe5_io_pipe_phv_out_data_143; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_144 = pipe5_io_pipe_phv_out_data_144; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_145 = pipe5_io_pipe_phv_out_data_145; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_146 = pipe5_io_pipe_phv_out_data_146; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_147 = pipe5_io_pipe_phv_out_data_147; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_148 = pipe5_io_pipe_phv_out_data_148; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_149 = pipe5_io_pipe_phv_out_data_149; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_150 = pipe5_io_pipe_phv_out_data_150; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_151 = pipe5_io_pipe_phv_out_data_151; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_152 = pipe5_io_pipe_phv_out_data_152; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_153 = pipe5_io_pipe_phv_out_data_153; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_154 = pipe5_io_pipe_phv_out_data_154; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_155 = pipe5_io_pipe_phv_out_data_155; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_156 = pipe5_io_pipe_phv_out_data_156; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_157 = pipe5_io_pipe_phv_out_data_157; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_158 = pipe5_io_pipe_phv_out_data_158; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_159 = pipe5_io_pipe_phv_out_data_159; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_160 = pipe5_io_pipe_phv_out_data_160; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_161 = pipe5_io_pipe_phv_out_data_161; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_162 = pipe5_io_pipe_phv_out_data_162; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_163 = pipe5_io_pipe_phv_out_data_163; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_164 = pipe5_io_pipe_phv_out_data_164; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_165 = pipe5_io_pipe_phv_out_data_165; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_166 = pipe5_io_pipe_phv_out_data_166; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_167 = pipe5_io_pipe_phv_out_data_167; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_168 = pipe5_io_pipe_phv_out_data_168; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_169 = pipe5_io_pipe_phv_out_data_169; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_170 = pipe5_io_pipe_phv_out_data_170; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_171 = pipe5_io_pipe_phv_out_data_171; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_172 = pipe5_io_pipe_phv_out_data_172; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_173 = pipe5_io_pipe_phv_out_data_173; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_174 = pipe5_io_pipe_phv_out_data_174; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_175 = pipe5_io_pipe_phv_out_data_175; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_176 = pipe5_io_pipe_phv_out_data_176; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_177 = pipe5_io_pipe_phv_out_data_177; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_178 = pipe5_io_pipe_phv_out_data_178; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_179 = pipe5_io_pipe_phv_out_data_179; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_180 = pipe5_io_pipe_phv_out_data_180; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_181 = pipe5_io_pipe_phv_out_data_181; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_182 = pipe5_io_pipe_phv_out_data_182; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_183 = pipe5_io_pipe_phv_out_data_183; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_184 = pipe5_io_pipe_phv_out_data_184; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_185 = pipe5_io_pipe_phv_out_data_185; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_186 = pipe5_io_pipe_phv_out_data_186; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_187 = pipe5_io_pipe_phv_out_data_187; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_188 = pipe5_io_pipe_phv_out_data_188; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_189 = pipe5_io_pipe_phv_out_data_189; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_190 = pipe5_io_pipe_phv_out_data_190; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_191 = pipe5_io_pipe_phv_out_data_191; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_192 = pipe5_io_pipe_phv_out_data_192; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_193 = pipe5_io_pipe_phv_out_data_193; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_194 = pipe5_io_pipe_phv_out_data_194; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_195 = pipe5_io_pipe_phv_out_data_195; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_196 = pipe5_io_pipe_phv_out_data_196; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_197 = pipe5_io_pipe_phv_out_data_197; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_198 = pipe5_io_pipe_phv_out_data_198; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_199 = pipe5_io_pipe_phv_out_data_199; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_200 = pipe5_io_pipe_phv_out_data_200; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_201 = pipe5_io_pipe_phv_out_data_201; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_202 = pipe5_io_pipe_phv_out_data_202; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_203 = pipe5_io_pipe_phv_out_data_203; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_204 = pipe5_io_pipe_phv_out_data_204; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_205 = pipe5_io_pipe_phv_out_data_205; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_206 = pipe5_io_pipe_phv_out_data_206; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_207 = pipe5_io_pipe_phv_out_data_207; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_208 = pipe5_io_pipe_phv_out_data_208; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_209 = pipe5_io_pipe_phv_out_data_209; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_210 = pipe5_io_pipe_phv_out_data_210; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_211 = pipe5_io_pipe_phv_out_data_211; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_212 = pipe5_io_pipe_phv_out_data_212; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_213 = pipe5_io_pipe_phv_out_data_213; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_214 = pipe5_io_pipe_phv_out_data_214; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_215 = pipe5_io_pipe_phv_out_data_215; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_216 = pipe5_io_pipe_phv_out_data_216; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_217 = pipe5_io_pipe_phv_out_data_217; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_218 = pipe5_io_pipe_phv_out_data_218; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_219 = pipe5_io_pipe_phv_out_data_219; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_220 = pipe5_io_pipe_phv_out_data_220; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_221 = pipe5_io_pipe_phv_out_data_221; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_222 = pipe5_io_pipe_phv_out_data_222; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_223 = pipe5_io_pipe_phv_out_data_223; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_224 = pipe5_io_pipe_phv_out_data_224; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_225 = pipe5_io_pipe_phv_out_data_225; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_226 = pipe5_io_pipe_phv_out_data_226; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_227 = pipe5_io_pipe_phv_out_data_227; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_228 = pipe5_io_pipe_phv_out_data_228; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_229 = pipe5_io_pipe_phv_out_data_229; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_230 = pipe5_io_pipe_phv_out_data_230; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_231 = pipe5_io_pipe_phv_out_data_231; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_232 = pipe5_io_pipe_phv_out_data_232; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_233 = pipe5_io_pipe_phv_out_data_233; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_234 = pipe5_io_pipe_phv_out_data_234; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_235 = pipe5_io_pipe_phv_out_data_235; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_236 = pipe5_io_pipe_phv_out_data_236; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_237 = pipe5_io_pipe_phv_out_data_237; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_238 = pipe5_io_pipe_phv_out_data_238; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_239 = pipe5_io_pipe_phv_out_data_239; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_240 = pipe5_io_pipe_phv_out_data_240; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_241 = pipe5_io_pipe_phv_out_data_241; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_242 = pipe5_io_pipe_phv_out_data_242; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_243 = pipe5_io_pipe_phv_out_data_243; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_244 = pipe5_io_pipe_phv_out_data_244; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_245 = pipe5_io_pipe_phv_out_data_245; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_246 = pipe5_io_pipe_phv_out_data_246; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_247 = pipe5_io_pipe_phv_out_data_247; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_248 = pipe5_io_pipe_phv_out_data_248; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_249 = pipe5_io_pipe_phv_out_data_249; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_250 = pipe5_io_pipe_phv_out_data_250; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_251 = pipe5_io_pipe_phv_out_data_251; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_252 = pipe5_io_pipe_phv_out_data_252; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_253 = pipe5_io_pipe_phv_out_data_253; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_254 = pipe5_io_pipe_phv_out_data_254; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_255 = pipe5_io_pipe_phv_out_data_255; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_0 = pipe5_io_pipe_phv_out_header_0; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_1 = pipe5_io_pipe_phv_out_header_1; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_2 = pipe5_io_pipe_phv_out_header_2; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_3 = pipe5_io_pipe_phv_out_header_3; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_4 = pipe5_io_pipe_phv_out_header_4; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_5 = pipe5_io_pipe_phv_out_header_5; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_6 = pipe5_io_pipe_phv_out_header_6; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_7 = pipe5_io_pipe_phv_out_header_7; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_8 = pipe5_io_pipe_phv_out_header_8; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_9 = pipe5_io_pipe_phv_out_header_9; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_10 = pipe5_io_pipe_phv_out_header_10; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_11 = pipe5_io_pipe_phv_out_header_11; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_12 = pipe5_io_pipe_phv_out_header_12; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_13 = pipe5_io_pipe_phv_out_header_13; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_14 = pipe5_io_pipe_phv_out_header_14; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_15 = pipe5_io_pipe_phv_out_header_15; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_parse_current_state = pipe5_io_pipe_phv_out_parse_current_state; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_parse_current_offset = pipe5_io_pipe_phv_out_parse_current_offset; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_parse_transition_field = pipe5_io_pipe_phv_out_parse_transition_field; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_next_processor_id = pipe5_io_pipe_phv_out_next_processor_id; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_next_config_id = pipe5_io_pipe_phv_out_next_config_id; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_is_valid_processor = pipe5_io_pipe_phv_out_is_valid_processor; // @[hash.scala 158:27]
  assign pipe6_io_hash_depth_0 = hash_depth_0; // @[hash.scala 162:27]
  assign pipe6_io_hash_depth_1 = hash_depth_1; // @[hash.scala 162:27]
  assign pipe6_io_key_in = pipe5_io_key_out; // @[hash.scala 159:27]
  assign pipe6_io_sum_in = pipe5_io_sum_out; // @[hash.scala 160:27]
  assign pipe6_io_val_in = pipe5_io_val_out; // @[hash.scala 161:27]
  assign pipe7_clock = clock;
  assign pipe7_io_pipe_phv_in_data_0 = pipe6_io_pipe_phv_out_data_0; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_1 = pipe6_io_pipe_phv_out_data_1; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_2 = pipe6_io_pipe_phv_out_data_2; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_3 = pipe6_io_pipe_phv_out_data_3; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_4 = pipe6_io_pipe_phv_out_data_4; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_5 = pipe6_io_pipe_phv_out_data_5; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_6 = pipe6_io_pipe_phv_out_data_6; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_7 = pipe6_io_pipe_phv_out_data_7; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_8 = pipe6_io_pipe_phv_out_data_8; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_9 = pipe6_io_pipe_phv_out_data_9; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_10 = pipe6_io_pipe_phv_out_data_10; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_11 = pipe6_io_pipe_phv_out_data_11; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_12 = pipe6_io_pipe_phv_out_data_12; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_13 = pipe6_io_pipe_phv_out_data_13; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_14 = pipe6_io_pipe_phv_out_data_14; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_15 = pipe6_io_pipe_phv_out_data_15; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_16 = pipe6_io_pipe_phv_out_data_16; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_17 = pipe6_io_pipe_phv_out_data_17; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_18 = pipe6_io_pipe_phv_out_data_18; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_19 = pipe6_io_pipe_phv_out_data_19; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_20 = pipe6_io_pipe_phv_out_data_20; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_21 = pipe6_io_pipe_phv_out_data_21; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_22 = pipe6_io_pipe_phv_out_data_22; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_23 = pipe6_io_pipe_phv_out_data_23; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_24 = pipe6_io_pipe_phv_out_data_24; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_25 = pipe6_io_pipe_phv_out_data_25; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_26 = pipe6_io_pipe_phv_out_data_26; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_27 = pipe6_io_pipe_phv_out_data_27; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_28 = pipe6_io_pipe_phv_out_data_28; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_29 = pipe6_io_pipe_phv_out_data_29; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_30 = pipe6_io_pipe_phv_out_data_30; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_31 = pipe6_io_pipe_phv_out_data_31; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_32 = pipe6_io_pipe_phv_out_data_32; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_33 = pipe6_io_pipe_phv_out_data_33; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_34 = pipe6_io_pipe_phv_out_data_34; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_35 = pipe6_io_pipe_phv_out_data_35; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_36 = pipe6_io_pipe_phv_out_data_36; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_37 = pipe6_io_pipe_phv_out_data_37; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_38 = pipe6_io_pipe_phv_out_data_38; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_39 = pipe6_io_pipe_phv_out_data_39; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_40 = pipe6_io_pipe_phv_out_data_40; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_41 = pipe6_io_pipe_phv_out_data_41; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_42 = pipe6_io_pipe_phv_out_data_42; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_43 = pipe6_io_pipe_phv_out_data_43; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_44 = pipe6_io_pipe_phv_out_data_44; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_45 = pipe6_io_pipe_phv_out_data_45; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_46 = pipe6_io_pipe_phv_out_data_46; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_47 = pipe6_io_pipe_phv_out_data_47; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_48 = pipe6_io_pipe_phv_out_data_48; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_49 = pipe6_io_pipe_phv_out_data_49; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_50 = pipe6_io_pipe_phv_out_data_50; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_51 = pipe6_io_pipe_phv_out_data_51; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_52 = pipe6_io_pipe_phv_out_data_52; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_53 = pipe6_io_pipe_phv_out_data_53; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_54 = pipe6_io_pipe_phv_out_data_54; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_55 = pipe6_io_pipe_phv_out_data_55; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_56 = pipe6_io_pipe_phv_out_data_56; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_57 = pipe6_io_pipe_phv_out_data_57; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_58 = pipe6_io_pipe_phv_out_data_58; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_59 = pipe6_io_pipe_phv_out_data_59; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_60 = pipe6_io_pipe_phv_out_data_60; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_61 = pipe6_io_pipe_phv_out_data_61; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_62 = pipe6_io_pipe_phv_out_data_62; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_63 = pipe6_io_pipe_phv_out_data_63; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_64 = pipe6_io_pipe_phv_out_data_64; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_65 = pipe6_io_pipe_phv_out_data_65; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_66 = pipe6_io_pipe_phv_out_data_66; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_67 = pipe6_io_pipe_phv_out_data_67; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_68 = pipe6_io_pipe_phv_out_data_68; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_69 = pipe6_io_pipe_phv_out_data_69; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_70 = pipe6_io_pipe_phv_out_data_70; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_71 = pipe6_io_pipe_phv_out_data_71; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_72 = pipe6_io_pipe_phv_out_data_72; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_73 = pipe6_io_pipe_phv_out_data_73; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_74 = pipe6_io_pipe_phv_out_data_74; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_75 = pipe6_io_pipe_phv_out_data_75; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_76 = pipe6_io_pipe_phv_out_data_76; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_77 = pipe6_io_pipe_phv_out_data_77; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_78 = pipe6_io_pipe_phv_out_data_78; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_79 = pipe6_io_pipe_phv_out_data_79; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_80 = pipe6_io_pipe_phv_out_data_80; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_81 = pipe6_io_pipe_phv_out_data_81; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_82 = pipe6_io_pipe_phv_out_data_82; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_83 = pipe6_io_pipe_phv_out_data_83; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_84 = pipe6_io_pipe_phv_out_data_84; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_85 = pipe6_io_pipe_phv_out_data_85; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_86 = pipe6_io_pipe_phv_out_data_86; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_87 = pipe6_io_pipe_phv_out_data_87; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_88 = pipe6_io_pipe_phv_out_data_88; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_89 = pipe6_io_pipe_phv_out_data_89; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_90 = pipe6_io_pipe_phv_out_data_90; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_91 = pipe6_io_pipe_phv_out_data_91; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_92 = pipe6_io_pipe_phv_out_data_92; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_93 = pipe6_io_pipe_phv_out_data_93; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_94 = pipe6_io_pipe_phv_out_data_94; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_95 = pipe6_io_pipe_phv_out_data_95; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_96 = pipe6_io_pipe_phv_out_data_96; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_97 = pipe6_io_pipe_phv_out_data_97; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_98 = pipe6_io_pipe_phv_out_data_98; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_99 = pipe6_io_pipe_phv_out_data_99; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_100 = pipe6_io_pipe_phv_out_data_100; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_101 = pipe6_io_pipe_phv_out_data_101; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_102 = pipe6_io_pipe_phv_out_data_102; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_103 = pipe6_io_pipe_phv_out_data_103; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_104 = pipe6_io_pipe_phv_out_data_104; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_105 = pipe6_io_pipe_phv_out_data_105; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_106 = pipe6_io_pipe_phv_out_data_106; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_107 = pipe6_io_pipe_phv_out_data_107; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_108 = pipe6_io_pipe_phv_out_data_108; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_109 = pipe6_io_pipe_phv_out_data_109; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_110 = pipe6_io_pipe_phv_out_data_110; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_111 = pipe6_io_pipe_phv_out_data_111; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_112 = pipe6_io_pipe_phv_out_data_112; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_113 = pipe6_io_pipe_phv_out_data_113; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_114 = pipe6_io_pipe_phv_out_data_114; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_115 = pipe6_io_pipe_phv_out_data_115; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_116 = pipe6_io_pipe_phv_out_data_116; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_117 = pipe6_io_pipe_phv_out_data_117; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_118 = pipe6_io_pipe_phv_out_data_118; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_119 = pipe6_io_pipe_phv_out_data_119; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_120 = pipe6_io_pipe_phv_out_data_120; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_121 = pipe6_io_pipe_phv_out_data_121; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_122 = pipe6_io_pipe_phv_out_data_122; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_123 = pipe6_io_pipe_phv_out_data_123; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_124 = pipe6_io_pipe_phv_out_data_124; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_125 = pipe6_io_pipe_phv_out_data_125; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_126 = pipe6_io_pipe_phv_out_data_126; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_127 = pipe6_io_pipe_phv_out_data_127; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_128 = pipe6_io_pipe_phv_out_data_128; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_129 = pipe6_io_pipe_phv_out_data_129; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_130 = pipe6_io_pipe_phv_out_data_130; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_131 = pipe6_io_pipe_phv_out_data_131; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_132 = pipe6_io_pipe_phv_out_data_132; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_133 = pipe6_io_pipe_phv_out_data_133; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_134 = pipe6_io_pipe_phv_out_data_134; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_135 = pipe6_io_pipe_phv_out_data_135; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_136 = pipe6_io_pipe_phv_out_data_136; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_137 = pipe6_io_pipe_phv_out_data_137; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_138 = pipe6_io_pipe_phv_out_data_138; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_139 = pipe6_io_pipe_phv_out_data_139; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_140 = pipe6_io_pipe_phv_out_data_140; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_141 = pipe6_io_pipe_phv_out_data_141; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_142 = pipe6_io_pipe_phv_out_data_142; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_143 = pipe6_io_pipe_phv_out_data_143; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_144 = pipe6_io_pipe_phv_out_data_144; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_145 = pipe6_io_pipe_phv_out_data_145; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_146 = pipe6_io_pipe_phv_out_data_146; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_147 = pipe6_io_pipe_phv_out_data_147; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_148 = pipe6_io_pipe_phv_out_data_148; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_149 = pipe6_io_pipe_phv_out_data_149; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_150 = pipe6_io_pipe_phv_out_data_150; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_151 = pipe6_io_pipe_phv_out_data_151; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_152 = pipe6_io_pipe_phv_out_data_152; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_153 = pipe6_io_pipe_phv_out_data_153; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_154 = pipe6_io_pipe_phv_out_data_154; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_155 = pipe6_io_pipe_phv_out_data_155; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_156 = pipe6_io_pipe_phv_out_data_156; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_157 = pipe6_io_pipe_phv_out_data_157; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_158 = pipe6_io_pipe_phv_out_data_158; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_159 = pipe6_io_pipe_phv_out_data_159; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_160 = pipe6_io_pipe_phv_out_data_160; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_161 = pipe6_io_pipe_phv_out_data_161; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_162 = pipe6_io_pipe_phv_out_data_162; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_163 = pipe6_io_pipe_phv_out_data_163; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_164 = pipe6_io_pipe_phv_out_data_164; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_165 = pipe6_io_pipe_phv_out_data_165; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_166 = pipe6_io_pipe_phv_out_data_166; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_167 = pipe6_io_pipe_phv_out_data_167; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_168 = pipe6_io_pipe_phv_out_data_168; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_169 = pipe6_io_pipe_phv_out_data_169; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_170 = pipe6_io_pipe_phv_out_data_170; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_171 = pipe6_io_pipe_phv_out_data_171; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_172 = pipe6_io_pipe_phv_out_data_172; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_173 = pipe6_io_pipe_phv_out_data_173; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_174 = pipe6_io_pipe_phv_out_data_174; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_175 = pipe6_io_pipe_phv_out_data_175; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_176 = pipe6_io_pipe_phv_out_data_176; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_177 = pipe6_io_pipe_phv_out_data_177; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_178 = pipe6_io_pipe_phv_out_data_178; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_179 = pipe6_io_pipe_phv_out_data_179; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_180 = pipe6_io_pipe_phv_out_data_180; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_181 = pipe6_io_pipe_phv_out_data_181; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_182 = pipe6_io_pipe_phv_out_data_182; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_183 = pipe6_io_pipe_phv_out_data_183; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_184 = pipe6_io_pipe_phv_out_data_184; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_185 = pipe6_io_pipe_phv_out_data_185; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_186 = pipe6_io_pipe_phv_out_data_186; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_187 = pipe6_io_pipe_phv_out_data_187; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_188 = pipe6_io_pipe_phv_out_data_188; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_189 = pipe6_io_pipe_phv_out_data_189; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_190 = pipe6_io_pipe_phv_out_data_190; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_191 = pipe6_io_pipe_phv_out_data_191; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_192 = pipe6_io_pipe_phv_out_data_192; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_193 = pipe6_io_pipe_phv_out_data_193; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_194 = pipe6_io_pipe_phv_out_data_194; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_195 = pipe6_io_pipe_phv_out_data_195; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_196 = pipe6_io_pipe_phv_out_data_196; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_197 = pipe6_io_pipe_phv_out_data_197; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_198 = pipe6_io_pipe_phv_out_data_198; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_199 = pipe6_io_pipe_phv_out_data_199; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_200 = pipe6_io_pipe_phv_out_data_200; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_201 = pipe6_io_pipe_phv_out_data_201; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_202 = pipe6_io_pipe_phv_out_data_202; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_203 = pipe6_io_pipe_phv_out_data_203; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_204 = pipe6_io_pipe_phv_out_data_204; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_205 = pipe6_io_pipe_phv_out_data_205; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_206 = pipe6_io_pipe_phv_out_data_206; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_207 = pipe6_io_pipe_phv_out_data_207; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_208 = pipe6_io_pipe_phv_out_data_208; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_209 = pipe6_io_pipe_phv_out_data_209; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_210 = pipe6_io_pipe_phv_out_data_210; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_211 = pipe6_io_pipe_phv_out_data_211; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_212 = pipe6_io_pipe_phv_out_data_212; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_213 = pipe6_io_pipe_phv_out_data_213; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_214 = pipe6_io_pipe_phv_out_data_214; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_215 = pipe6_io_pipe_phv_out_data_215; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_216 = pipe6_io_pipe_phv_out_data_216; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_217 = pipe6_io_pipe_phv_out_data_217; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_218 = pipe6_io_pipe_phv_out_data_218; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_219 = pipe6_io_pipe_phv_out_data_219; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_220 = pipe6_io_pipe_phv_out_data_220; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_221 = pipe6_io_pipe_phv_out_data_221; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_222 = pipe6_io_pipe_phv_out_data_222; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_223 = pipe6_io_pipe_phv_out_data_223; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_224 = pipe6_io_pipe_phv_out_data_224; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_225 = pipe6_io_pipe_phv_out_data_225; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_226 = pipe6_io_pipe_phv_out_data_226; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_227 = pipe6_io_pipe_phv_out_data_227; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_228 = pipe6_io_pipe_phv_out_data_228; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_229 = pipe6_io_pipe_phv_out_data_229; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_230 = pipe6_io_pipe_phv_out_data_230; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_231 = pipe6_io_pipe_phv_out_data_231; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_232 = pipe6_io_pipe_phv_out_data_232; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_233 = pipe6_io_pipe_phv_out_data_233; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_234 = pipe6_io_pipe_phv_out_data_234; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_235 = pipe6_io_pipe_phv_out_data_235; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_236 = pipe6_io_pipe_phv_out_data_236; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_237 = pipe6_io_pipe_phv_out_data_237; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_238 = pipe6_io_pipe_phv_out_data_238; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_239 = pipe6_io_pipe_phv_out_data_239; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_240 = pipe6_io_pipe_phv_out_data_240; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_241 = pipe6_io_pipe_phv_out_data_241; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_242 = pipe6_io_pipe_phv_out_data_242; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_243 = pipe6_io_pipe_phv_out_data_243; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_244 = pipe6_io_pipe_phv_out_data_244; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_245 = pipe6_io_pipe_phv_out_data_245; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_246 = pipe6_io_pipe_phv_out_data_246; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_247 = pipe6_io_pipe_phv_out_data_247; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_248 = pipe6_io_pipe_phv_out_data_248; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_249 = pipe6_io_pipe_phv_out_data_249; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_250 = pipe6_io_pipe_phv_out_data_250; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_251 = pipe6_io_pipe_phv_out_data_251; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_252 = pipe6_io_pipe_phv_out_data_252; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_253 = pipe6_io_pipe_phv_out_data_253; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_254 = pipe6_io_pipe_phv_out_data_254; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_255 = pipe6_io_pipe_phv_out_data_255; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_0 = pipe6_io_pipe_phv_out_header_0; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_1 = pipe6_io_pipe_phv_out_header_1; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_2 = pipe6_io_pipe_phv_out_header_2; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_3 = pipe6_io_pipe_phv_out_header_3; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_4 = pipe6_io_pipe_phv_out_header_4; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_5 = pipe6_io_pipe_phv_out_header_5; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_6 = pipe6_io_pipe_phv_out_header_6; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_7 = pipe6_io_pipe_phv_out_header_7; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_8 = pipe6_io_pipe_phv_out_header_8; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_9 = pipe6_io_pipe_phv_out_header_9; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_10 = pipe6_io_pipe_phv_out_header_10; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_11 = pipe6_io_pipe_phv_out_header_11; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_12 = pipe6_io_pipe_phv_out_header_12; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_13 = pipe6_io_pipe_phv_out_header_13; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_14 = pipe6_io_pipe_phv_out_header_14; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_15 = pipe6_io_pipe_phv_out_header_15; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_parse_current_state = pipe6_io_pipe_phv_out_parse_current_state; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_parse_current_offset = pipe6_io_pipe_phv_out_parse_current_offset; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_parse_transition_field = pipe6_io_pipe_phv_out_parse_transition_field; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_next_processor_id = pipe6_io_pipe_phv_out_next_processor_id; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_next_config_id = pipe6_io_pipe_phv_out_next_config_id; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_is_valid_processor = pipe6_io_pipe_phv_out_is_valid_processor; // @[hash.scala 164:27]
  assign pipe7_io_hash_depth_0 = hash_depth_0; // @[hash.scala 168:27]
  assign pipe7_io_hash_depth_1 = hash_depth_1; // @[hash.scala 168:27]
  assign pipe7_io_key_in = pipe6_io_key_out; // @[hash.scala 165:27]
  assign pipe7_io_sum_in = pipe6_io_sum_out; // @[hash.scala 166:27]
  assign pipe7_io_val_in = pipe6_io_val_out; // @[hash.scala 167:27]
  assign pipe8_clock = clock;
  assign pipe8_io_pipe_phv_in_data_0 = pipe7_io_pipe_phv_out_data_0; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_1 = pipe7_io_pipe_phv_out_data_1; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_2 = pipe7_io_pipe_phv_out_data_2; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_3 = pipe7_io_pipe_phv_out_data_3; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_4 = pipe7_io_pipe_phv_out_data_4; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_5 = pipe7_io_pipe_phv_out_data_5; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_6 = pipe7_io_pipe_phv_out_data_6; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_7 = pipe7_io_pipe_phv_out_data_7; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_8 = pipe7_io_pipe_phv_out_data_8; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_9 = pipe7_io_pipe_phv_out_data_9; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_10 = pipe7_io_pipe_phv_out_data_10; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_11 = pipe7_io_pipe_phv_out_data_11; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_12 = pipe7_io_pipe_phv_out_data_12; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_13 = pipe7_io_pipe_phv_out_data_13; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_14 = pipe7_io_pipe_phv_out_data_14; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_15 = pipe7_io_pipe_phv_out_data_15; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_16 = pipe7_io_pipe_phv_out_data_16; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_17 = pipe7_io_pipe_phv_out_data_17; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_18 = pipe7_io_pipe_phv_out_data_18; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_19 = pipe7_io_pipe_phv_out_data_19; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_20 = pipe7_io_pipe_phv_out_data_20; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_21 = pipe7_io_pipe_phv_out_data_21; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_22 = pipe7_io_pipe_phv_out_data_22; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_23 = pipe7_io_pipe_phv_out_data_23; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_24 = pipe7_io_pipe_phv_out_data_24; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_25 = pipe7_io_pipe_phv_out_data_25; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_26 = pipe7_io_pipe_phv_out_data_26; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_27 = pipe7_io_pipe_phv_out_data_27; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_28 = pipe7_io_pipe_phv_out_data_28; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_29 = pipe7_io_pipe_phv_out_data_29; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_30 = pipe7_io_pipe_phv_out_data_30; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_31 = pipe7_io_pipe_phv_out_data_31; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_32 = pipe7_io_pipe_phv_out_data_32; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_33 = pipe7_io_pipe_phv_out_data_33; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_34 = pipe7_io_pipe_phv_out_data_34; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_35 = pipe7_io_pipe_phv_out_data_35; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_36 = pipe7_io_pipe_phv_out_data_36; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_37 = pipe7_io_pipe_phv_out_data_37; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_38 = pipe7_io_pipe_phv_out_data_38; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_39 = pipe7_io_pipe_phv_out_data_39; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_40 = pipe7_io_pipe_phv_out_data_40; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_41 = pipe7_io_pipe_phv_out_data_41; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_42 = pipe7_io_pipe_phv_out_data_42; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_43 = pipe7_io_pipe_phv_out_data_43; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_44 = pipe7_io_pipe_phv_out_data_44; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_45 = pipe7_io_pipe_phv_out_data_45; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_46 = pipe7_io_pipe_phv_out_data_46; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_47 = pipe7_io_pipe_phv_out_data_47; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_48 = pipe7_io_pipe_phv_out_data_48; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_49 = pipe7_io_pipe_phv_out_data_49; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_50 = pipe7_io_pipe_phv_out_data_50; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_51 = pipe7_io_pipe_phv_out_data_51; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_52 = pipe7_io_pipe_phv_out_data_52; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_53 = pipe7_io_pipe_phv_out_data_53; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_54 = pipe7_io_pipe_phv_out_data_54; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_55 = pipe7_io_pipe_phv_out_data_55; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_56 = pipe7_io_pipe_phv_out_data_56; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_57 = pipe7_io_pipe_phv_out_data_57; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_58 = pipe7_io_pipe_phv_out_data_58; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_59 = pipe7_io_pipe_phv_out_data_59; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_60 = pipe7_io_pipe_phv_out_data_60; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_61 = pipe7_io_pipe_phv_out_data_61; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_62 = pipe7_io_pipe_phv_out_data_62; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_63 = pipe7_io_pipe_phv_out_data_63; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_64 = pipe7_io_pipe_phv_out_data_64; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_65 = pipe7_io_pipe_phv_out_data_65; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_66 = pipe7_io_pipe_phv_out_data_66; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_67 = pipe7_io_pipe_phv_out_data_67; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_68 = pipe7_io_pipe_phv_out_data_68; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_69 = pipe7_io_pipe_phv_out_data_69; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_70 = pipe7_io_pipe_phv_out_data_70; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_71 = pipe7_io_pipe_phv_out_data_71; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_72 = pipe7_io_pipe_phv_out_data_72; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_73 = pipe7_io_pipe_phv_out_data_73; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_74 = pipe7_io_pipe_phv_out_data_74; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_75 = pipe7_io_pipe_phv_out_data_75; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_76 = pipe7_io_pipe_phv_out_data_76; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_77 = pipe7_io_pipe_phv_out_data_77; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_78 = pipe7_io_pipe_phv_out_data_78; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_79 = pipe7_io_pipe_phv_out_data_79; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_80 = pipe7_io_pipe_phv_out_data_80; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_81 = pipe7_io_pipe_phv_out_data_81; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_82 = pipe7_io_pipe_phv_out_data_82; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_83 = pipe7_io_pipe_phv_out_data_83; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_84 = pipe7_io_pipe_phv_out_data_84; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_85 = pipe7_io_pipe_phv_out_data_85; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_86 = pipe7_io_pipe_phv_out_data_86; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_87 = pipe7_io_pipe_phv_out_data_87; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_88 = pipe7_io_pipe_phv_out_data_88; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_89 = pipe7_io_pipe_phv_out_data_89; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_90 = pipe7_io_pipe_phv_out_data_90; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_91 = pipe7_io_pipe_phv_out_data_91; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_92 = pipe7_io_pipe_phv_out_data_92; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_93 = pipe7_io_pipe_phv_out_data_93; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_94 = pipe7_io_pipe_phv_out_data_94; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_95 = pipe7_io_pipe_phv_out_data_95; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_96 = pipe7_io_pipe_phv_out_data_96; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_97 = pipe7_io_pipe_phv_out_data_97; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_98 = pipe7_io_pipe_phv_out_data_98; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_99 = pipe7_io_pipe_phv_out_data_99; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_100 = pipe7_io_pipe_phv_out_data_100; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_101 = pipe7_io_pipe_phv_out_data_101; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_102 = pipe7_io_pipe_phv_out_data_102; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_103 = pipe7_io_pipe_phv_out_data_103; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_104 = pipe7_io_pipe_phv_out_data_104; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_105 = pipe7_io_pipe_phv_out_data_105; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_106 = pipe7_io_pipe_phv_out_data_106; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_107 = pipe7_io_pipe_phv_out_data_107; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_108 = pipe7_io_pipe_phv_out_data_108; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_109 = pipe7_io_pipe_phv_out_data_109; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_110 = pipe7_io_pipe_phv_out_data_110; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_111 = pipe7_io_pipe_phv_out_data_111; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_112 = pipe7_io_pipe_phv_out_data_112; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_113 = pipe7_io_pipe_phv_out_data_113; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_114 = pipe7_io_pipe_phv_out_data_114; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_115 = pipe7_io_pipe_phv_out_data_115; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_116 = pipe7_io_pipe_phv_out_data_116; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_117 = pipe7_io_pipe_phv_out_data_117; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_118 = pipe7_io_pipe_phv_out_data_118; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_119 = pipe7_io_pipe_phv_out_data_119; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_120 = pipe7_io_pipe_phv_out_data_120; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_121 = pipe7_io_pipe_phv_out_data_121; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_122 = pipe7_io_pipe_phv_out_data_122; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_123 = pipe7_io_pipe_phv_out_data_123; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_124 = pipe7_io_pipe_phv_out_data_124; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_125 = pipe7_io_pipe_phv_out_data_125; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_126 = pipe7_io_pipe_phv_out_data_126; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_127 = pipe7_io_pipe_phv_out_data_127; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_128 = pipe7_io_pipe_phv_out_data_128; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_129 = pipe7_io_pipe_phv_out_data_129; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_130 = pipe7_io_pipe_phv_out_data_130; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_131 = pipe7_io_pipe_phv_out_data_131; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_132 = pipe7_io_pipe_phv_out_data_132; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_133 = pipe7_io_pipe_phv_out_data_133; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_134 = pipe7_io_pipe_phv_out_data_134; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_135 = pipe7_io_pipe_phv_out_data_135; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_136 = pipe7_io_pipe_phv_out_data_136; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_137 = pipe7_io_pipe_phv_out_data_137; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_138 = pipe7_io_pipe_phv_out_data_138; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_139 = pipe7_io_pipe_phv_out_data_139; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_140 = pipe7_io_pipe_phv_out_data_140; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_141 = pipe7_io_pipe_phv_out_data_141; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_142 = pipe7_io_pipe_phv_out_data_142; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_143 = pipe7_io_pipe_phv_out_data_143; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_144 = pipe7_io_pipe_phv_out_data_144; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_145 = pipe7_io_pipe_phv_out_data_145; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_146 = pipe7_io_pipe_phv_out_data_146; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_147 = pipe7_io_pipe_phv_out_data_147; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_148 = pipe7_io_pipe_phv_out_data_148; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_149 = pipe7_io_pipe_phv_out_data_149; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_150 = pipe7_io_pipe_phv_out_data_150; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_151 = pipe7_io_pipe_phv_out_data_151; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_152 = pipe7_io_pipe_phv_out_data_152; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_153 = pipe7_io_pipe_phv_out_data_153; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_154 = pipe7_io_pipe_phv_out_data_154; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_155 = pipe7_io_pipe_phv_out_data_155; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_156 = pipe7_io_pipe_phv_out_data_156; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_157 = pipe7_io_pipe_phv_out_data_157; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_158 = pipe7_io_pipe_phv_out_data_158; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_159 = pipe7_io_pipe_phv_out_data_159; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_160 = pipe7_io_pipe_phv_out_data_160; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_161 = pipe7_io_pipe_phv_out_data_161; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_162 = pipe7_io_pipe_phv_out_data_162; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_163 = pipe7_io_pipe_phv_out_data_163; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_164 = pipe7_io_pipe_phv_out_data_164; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_165 = pipe7_io_pipe_phv_out_data_165; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_166 = pipe7_io_pipe_phv_out_data_166; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_167 = pipe7_io_pipe_phv_out_data_167; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_168 = pipe7_io_pipe_phv_out_data_168; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_169 = pipe7_io_pipe_phv_out_data_169; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_170 = pipe7_io_pipe_phv_out_data_170; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_171 = pipe7_io_pipe_phv_out_data_171; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_172 = pipe7_io_pipe_phv_out_data_172; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_173 = pipe7_io_pipe_phv_out_data_173; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_174 = pipe7_io_pipe_phv_out_data_174; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_175 = pipe7_io_pipe_phv_out_data_175; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_176 = pipe7_io_pipe_phv_out_data_176; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_177 = pipe7_io_pipe_phv_out_data_177; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_178 = pipe7_io_pipe_phv_out_data_178; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_179 = pipe7_io_pipe_phv_out_data_179; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_180 = pipe7_io_pipe_phv_out_data_180; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_181 = pipe7_io_pipe_phv_out_data_181; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_182 = pipe7_io_pipe_phv_out_data_182; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_183 = pipe7_io_pipe_phv_out_data_183; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_184 = pipe7_io_pipe_phv_out_data_184; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_185 = pipe7_io_pipe_phv_out_data_185; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_186 = pipe7_io_pipe_phv_out_data_186; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_187 = pipe7_io_pipe_phv_out_data_187; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_188 = pipe7_io_pipe_phv_out_data_188; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_189 = pipe7_io_pipe_phv_out_data_189; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_190 = pipe7_io_pipe_phv_out_data_190; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_191 = pipe7_io_pipe_phv_out_data_191; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_192 = pipe7_io_pipe_phv_out_data_192; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_193 = pipe7_io_pipe_phv_out_data_193; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_194 = pipe7_io_pipe_phv_out_data_194; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_195 = pipe7_io_pipe_phv_out_data_195; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_196 = pipe7_io_pipe_phv_out_data_196; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_197 = pipe7_io_pipe_phv_out_data_197; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_198 = pipe7_io_pipe_phv_out_data_198; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_199 = pipe7_io_pipe_phv_out_data_199; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_200 = pipe7_io_pipe_phv_out_data_200; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_201 = pipe7_io_pipe_phv_out_data_201; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_202 = pipe7_io_pipe_phv_out_data_202; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_203 = pipe7_io_pipe_phv_out_data_203; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_204 = pipe7_io_pipe_phv_out_data_204; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_205 = pipe7_io_pipe_phv_out_data_205; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_206 = pipe7_io_pipe_phv_out_data_206; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_207 = pipe7_io_pipe_phv_out_data_207; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_208 = pipe7_io_pipe_phv_out_data_208; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_209 = pipe7_io_pipe_phv_out_data_209; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_210 = pipe7_io_pipe_phv_out_data_210; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_211 = pipe7_io_pipe_phv_out_data_211; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_212 = pipe7_io_pipe_phv_out_data_212; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_213 = pipe7_io_pipe_phv_out_data_213; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_214 = pipe7_io_pipe_phv_out_data_214; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_215 = pipe7_io_pipe_phv_out_data_215; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_216 = pipe7_io_pipe_phv_out_data_216; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_217 = pipe7_io_pipe_phv_out_data_217; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_218 = pipe7_io_pipe_phv_out_data_218; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_219 = pipe7_io_pipe_phv_out_data_219; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_220 = pipe7_io_pipe_phv_out_data_220; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_221 = pipe7_io_pipe_phv_out_data_221; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_222 = pipe7_io_pipe_phv_out_data_222; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_223 = pipe7_io_pipe_phv_out_data_223; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_224 = pipe7_io_pipe_phv_out_data_224; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_225 = pipe7_io_pipe_phv_out_data_225; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_226 = pipe7_io_pipe_phv_out_data_226; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_227 = pipe7_io_pipe_phv_out_data_227; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_228 = pipe7_io_pipe_phv_out_data_228; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_229 = pipe7_io_pipe_phv_out_data_229; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_230 = pipe7_io_pipe_phv_out_data_230; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_231 = pipe7_io_pipe_phv_out_data_231; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_232 = pipe7_io_pipe_phv_out_data_232; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_233 = pipe7_io_pipe_phv_out_data_233; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_234 = pipe7_io_pipe_phv_out_data_234; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_235 = pipe7_io_pipe_phv_out_data_235; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_236 = pipe7_io_pipe_phv_out_data_236; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_237 = pipe7_io_pipe_phv_out_data_237; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_238 = pipe7_io_pipe_phv_out_data_238; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_239 = pipe7_io_pipe_phv_out_data_239; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_240 = pipe7_io_pipe_phv_out_data_240; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_241 = pipe7_io_pipe_phv_out_data_241; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_242 = pipe7_io_pipe_phv_out_data_242; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_243 = pipe7_io_pipe_phv_out_data_243; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_244 = pipe7_io_pipe_phv_out_data_244; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_245 = pipe7_io_pipe_phv_out_data_245; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_246 = pipe7_io_pipe_phv_out_data_246; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_247 = pipe7_io_pipe_phv_out_data_247; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_248 = pipe7_io_pipe_phv_out_data_248; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_249 = pipe7_io_pipe_phv_out_data_249; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_250 = pipe7_io_pipe_phv_out_data_250; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_251 = pipe7_io_pipe_phv_out_data_251; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_252 = pipe7_io_pipe_phv_out_data_252; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_253 = pipe7_io_pipe_phv_out_data_253; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_254 = pipe7_io_pipe_phv_out_data_254; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_255 = pipe7_io_pipe_phv_out_data_255; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_0 = pipe7_io_pipe_phv_out_header_0; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_1 = pipe7_io_pipe_phv_out_header_1; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_2 = pipe7_io_pipe_phv_out_header_2; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_3 = pipe7_io_pipe_phv_out_header_3; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_4 = pipe7_io_pipe_phv_out_header_4; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_5 = pipe7_io_pipe_phv_out_header_5; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_6 = pipe7_io_pipe_phv_out_header_6; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_7 = pipe7_io_pipe_phv_out_header_7; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_8 = pipe7_io_pipe_phv_out_header_8; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_9 = pipe7_io_pipe_phv_out_header_9; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_10 = pipe7_io_pipe_phv_out_header_10; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_11 = pipe7_io_pipe_phv_out_header_11; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_12 = pipe7_io_pipe_phv_out_header_12; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_13 = pipe7_io_pipe_phv_out_header_13; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_14 = pipe7_io_pipe_phv_out_header_14; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_15 = pipe7_io_pipe_phv_out_header_15; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_parse_current_state = pipe7_io_pipe_phv_out_parse_current_state; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_parse_current_offset = pipe7_io_pipe_phv_out_parse_current_offset; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_parse_transition_field = pipe7_io_pipe_phv_out_parse_transition_field; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_next_processor_id = pipe7_io_pipe_phv_out_next_processor_id; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_next_config_id = pipe7_io_pipe_phv_out_next_config_id; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_is_valid_processor = pipe7_io_pipe_phv_out_is_valid_processor; // @[hash.scala 170:27]
  assign pipe8_io_hash_depth_0 = hash_depth_0; // @[hash.scala 174:27]
  assign pipe8_io_hash_depth_1 = hash_depth_1; // @[hash.scala 174:27]
  assign pipe8_io_key_in = pipe7_io_key_out; // @[hash.scala 171:27]
  assign pipe8_io_sum_in = pipe7_io_sum_out; // @[hash.scala 172:27]
  assign pipe8_io_val_in = pipe7_io_val_out; // @[hash.scala 173:27]
  always @(posedge clock) begin
    if (io_mod_hash_depth_mod) begin // @[hash.scala 19:34]
      if (~io_mod_config_id) begin // @[hash.scala 20:38]
        hash_depth_0 <= io_mod_hash_depth; // @[hash.scala 20:38]
      end
    end
    if (io_mod_hash_depth_mod) begin // @[hash.scala 19:34]
      if (io_mod_config_id) begin // @[hash.scala 20:38]
        hash_depth_1 <= io_mod_hash_depth; // @[hash.scala 20:38]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  hash_depth_0 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  hash_depth_1 = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
