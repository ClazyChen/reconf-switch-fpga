module Processor(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [7:0]  io_pipe_phv_in_data_256,
  input  [7:0]  io_pipe_phv_in_data_257,
  input  [7:0]  io_pipe_phv_in_data_258,
  input  [7:0]  io_pipe_phv_in_data_259,
  input  [7:0]  io_pipe_phv_in_data_260,
  input  [7:0]  io_pipe_phv_in_data_261,
  input  [7:0]  io_pipe_phv_in_data_262,
  input  [7:0]  io_pipe_phv_in_data_263,
  input  [7:0]  io_pipe_phv_in_data_264,
  input  [7:0]  io_pipe_phv_in_data_265,
  input  [7:0]  io_pipe_phv_in_data_266,
  input  [7:0]  io_pipe_phv_in_data_267,
  input  [7:0]  io_pipe_phv_in_data_268,
  input  [7:0]  io_pipe_phv_in_data_269,
  input  [7:0]  io_pipe_phv_in_data_270,
  input  [7:0]  io_pipe_phv_in_data_271,
  input  [7:0]  io_pipe_phv_in_data_272,
  input  [7:0]  io_pipe_phv_in_data_273,
  input  [7:0]  io_pipe_phv_in_data_274,
  input  [7:0]  io_pipe_phv_in_data_275,
  input  [7:0]  io_pipe_phv_in_data_276,
  input  [7:0]  io_pipe_phv_in_data_277,
  input  [7:0]  io_pipe_phv_in_data_278,
  input  [7:0]  io_pipe_phv_in_data_279,
  input  [7:0]  io_pipe_phv_in_data_280,
  input  [7:0]  io_pipe_phv_in_data_281,
  input  [7:0]  io_pipe_phv_in_data_282,
  input  [7:0]  io_pipe_phv_in_data_283,
  input  [7:0]  io_pipe_phv_in_data_284,
  input  [7:0]  io_pipe_phv_in_data_285,
  input  [7:0]  io_pipe_phv_in_data_286,
  input  [7:0]  io_pipe_phv_in_data_287,
  input  [7:0]  io_pipe_phv_in_data_288,
  input  [7:0]  io_pipe_phv_in_data_289,
  input  [7:0]  io_pipe_phv_in_data_290,
  input  [7:0]  io_pipe_phv_in_data_291,
  input  [7:0]  io_pipe_phv_in_data_292,
  input  [7:0]  io_pipe_phv_in_data_293,
  input  [7:0]  io_pipe_phv_in_data_294,
  input  [7:0]  io_pipe_phv_in_data_295,
  input  [7:0]  io_pipe_phv_in_data_296,
  input  [7:0]  io_pipe_phv_in_data_297,
  input  [7:0]  io_pipe_phv_in_data_298,
  input  [7:0]  io_pipe_phv_in_data_299,
  input  [7:0]  io_pipe_phv_in_data_300,
  input  [7:0]  io_pipe_phv_in_data_301,
  input  [7:0]  io_pipe_phv_in_data_302,
  input  [7:0]  io_pipe_phv_in_data_303,
  input  [7:0]  io_pipe_phv_in_data_304,
  input  [7:0]  io_pipe_phv_in_data_305,
  input  [7:0]  io_pipe_phv_in_data_306,
  input  [7:0]  io_pipe_phv_in_data_307,
  input  [7:0]  io_pipe_phv_in_data_308,
  input  [7:0]  io_pipe_phv_in_data_309,
  input  [7:0]  io_pipe_phv_in_data_310,
  input  [7:0]  io_pipe_phv_in_data_311,
  input  [7:0]  io_pipe_phv_in_data_312,
  input  [7:0]  io_pipe_phv_in_data_313,
  input  [7:0]  io_pipe_phv_in_data_314,
  input  [7:0]  io_pipe_phv_in_data_315,
  input  [7:0]  io_pipe_phv_in_data_316,
  input  [7:0]  io_pipe_phv_in_data_317,
  input  [7:0]  io_pipe_phv_in_data_318,
  input  [7:0]  io_pipe_phv_in_data_319,
  input  [7:0]  io_pipe_phv_in_data_320,
  input  [7:0]  io_pipe_phv_in_data_321,
  input  [7:0]  io_pipe_phv_in_data_322,
  input  [7:0]  io_pipe_phv_in_data_323,
  input  [7:0]  io_pipe_phv_in_data_324,
  input  [7:0]  io_pipe_phv_in_data_325,
  input  [7:0]  io_pipe_phv_in_data_326,
  input  [7:0]  io_pipe_phv_in_data_327,
  input  [7:0]  io_pipe_phv_in_data_328,
  input  [7:0]  io_pipe_phv_in_data_329,
  input  [7:0]  io_pipe_phv_in_data_330,
  input  [7:0]  io_pipe_phv_in_data_331,
  input  [7:0]  io_pipe_phv_in_data_332,
  input  [7:0]  io_pipe_phv_in_data_333,
  input  [7:0]  io_pipe_phv_in_data_334,
  input  [7:0]  io_pipe_phv_in_data_335,
  input  [7:0]  io_pipe_phv_in_data_336,
  input  [7:0]  io_pipe_phv_in_data_337,
  input  [7:0]  io_pipe_phv_in_data_338,
  input  [7:0]  io_pipe_phv_in_data_339,
  input  [7:0]  io_pipe_phv_in_data_340,
  input  [7:0]  io_pipe_phv_in_data_341,
  input  [7:0]  io_pipe_phv_in_data_342,
  input  [7:0]  io_pipe_phv_in_data_343,
  input  [7:0]  io_pipe_phv_in_data_344,
  input  [7:0]  io_pipe_phv_in_data_345,
  input  [7:0]  io_pipe_phv_in_data_346,
  input  [7:0]  io_pipe_phv_in_data_347,
  input  [7:0]  io_pipe_phv_in_data_348,
  input  [7:0]  io_pipe_phv_in_data_349,
  input  [7:0]  io_pipe_phv_in_data_350,
  input  [7:0]  io_pipe_phv_in_data_351,
  input  [7:0]  io_pipe_phv_in_data_352,
  input  [7:0]  io_pipe_phv_in_data_353,
  input  [7:0]  io_pipe_phv_in_data_354,
  input  [7:0]  io_pipe_phv_in_data_355,
  input  [7:0]  io_pipe_phv_in_data_356,
  input  [7:0]  io_pipe_phv_in_data_357,
  input  [7:0]  io_pipe_phv_in_data_358,
  input  [7:0]  io_pipe_phv_in_data_359,
  input  [7:0]  io_pipe_phv_in_data_360,
  input  [7:0]  io_pipe_phv_in_data_361,
  input  [7:0]  io_pipe_phv_in_data_362,
  input  [7:0]  io_pipe_phv_in_data_363,
  input  [7:0]  io_pipe_phv_in_data_364,
  input  [7:0]  io_pipe_phv_in_data_365,
  input  [7:0]  io_pipe_phv_in_data_366,
  input  [7:0]  io_pipe_phv_in_data_367,
  input  [7:0]  io_pipe_phv_in_data_368,
  input  [7:0]  io_pipe_phv_in_data_369,
  input  [7:0]  io_pipe_phv_in_data_370,
  input  [7:0]  io_pipe_phv_in_data_371,
  input  [7:0]  io_pipe_phv_in_data_372,
  input  [7:0]  io_pipe_phv_in_data_373,
  input  [7:0]  io_pipe_phv_in_data_374,
  input  [7:0]  io_pipe_phv_in_data_375,
  input  [7:0]  io_pipe_phv_in_data_376,
  input  [7:0]  io_pipe_phv_in_data_377,
  input  [7:0]  io_pipe_phv_in_data_378,
  input  [7:0]  io_pipe_phv_in_data_379,
  input  [7:0]  io_pipe_phv_in_data_380,
  input  [7:0]  io_pipe_phv_in_data_381,
  input  [7:0]  io_pipe_phv_in_data_382,
  input  [7:0]  io_pipe_phv_in_data_383,
  input  [7:0]  io_pipe_phv_in_data_384,
  input  [7:0]  io_pipe_phv_in_data_385,
  input  [7:0]  io_pipe_phv_in_data_386,
  input  [7:0]  io_pipe_phv_in_data_387,
  input  [7:0]  io_pipe_phv_in_data_388,
  input  [7:0]  io_pipe_phv_in_data_389,
  input  [7:0]  io_pipe_phv_in_data_390,
  input  [7:0]  io_pipe_phv_in_data_391,
  input  [7:0]  io_pipe_phv_in_data_392,
  input  [7:0]  io_pipe_phv_in_data_393,
  input  [7:0]  io_pipe_phv_in_data_394,
  input  [7:0]  io_pipe_phv_in_data_395,
  input  [7:0]  io_pipe_phv_in_data_396,
  input  [7:0]  io_pipe_phv_in_data_397,
  input  [7:0]  io_pipe_phv_in_data_398,
  input  [7:0]  io_pipe_phv_in_data_399,
  input  [7:0]  io_pipe_phv_in_data_400,
  input  [7:0]  io_pipe_phv_in_data_401,
  input  [7:0]  io_pipe_phv_in_data_402,
  input  [7:0]  io_pipe_phv_in_data_403,
  input  [7:0]  io_pipe_phv_in_data_404,
  input  [7:0]  io_pipe_phv_in_data_405,
  input  [7:0]  io_pipe_phv_in_data_406,
  input  [7:0]  io_pipe_phv_in_data_407,
  input  [7:0]  io_pipe_phv_in_data_408,
  input  [7:0]  io_pipe_phv_in_data_409,
  input  [7:0]  io_pipe_phv_in_data_410,
  input  [7:0]  io_pipe_phv_in_data_411,
  input  [7:0]  io_pipe_phv_in_data_412,
  input  [7:0]  io_pipe_phv_in_data_413,
  input  [7:0]  io_pipe_phv_in_data_414,
  input  [7:0]  io_pipe_phv_in_data_415,
  input  [7:0]  io_pipe_phv_in_data_416,
  input  [7:0]  io_pipe_phv_in_data_417,
  input  [7:0]  io_pipe_phv_in_data_418,
  input  [7:0]  io_pipe_phv_in_data_419,
  input  [7:0]  io_pipe_phv_in_data_420,
  input  [7:0]  io_pipe_phv_in_data_421,
  input  [7:0]  io_pipe_phv_in_data_422,
  input  [7:0]  io_pipe_phv_in_data_423,
  input  [7:0]  io_pipe_phv_in_data_424,
  input  [7:0]  io_pipe_phv_in_data_425,
  input  [7:0]  io_pipe_phv_in_data_426,
  input  [7:0]  io_pipe_phv_in_data_427,
  input  [7:0]  io_pipe_phv_in_data_428,
  input  [7:0]  io_pipe_phv_in_data_429,
  input  [7:0]  io_pipe_phv_in_data_430,
  input  [7:0]  io_pipe_phv_in_data_431,
  input  [7:0]  io_pipe_phv_in_data_432,
  input  [7:0]  io_pipe_phv_in_data_433,
  input  [7:0]  io_pipe_phv_in_data_434,
  input  [7:0]  io_pipe_phv_in_data_435,
  input  [7:0]  io_pipe_phv_in_data_436,
  input  [7:0]  io_pipe_phv_in_data_437,
  input  [7:0]  io_pipe_phv_in_data_438,
  input  [7:0]  io_pipe_phv_in_data_439,
  input  [7:0]  io_pipe_phv_in_data_440,
  input  [7:0]  io_pipe_phv_in_data_441,
  input  [7:0]  io_pipe_phv_in_data_442,
  input  [7:0]  io_pipe_phv_in_data_443,
  input  [7:0]  io_pipe_phv_in_data_444,
  input  [7:0]  io_pipe_phv_in_data_445,
  input  [7:0]  io_pipe_phv_in_data_446,
  input  [7:0]  io_pipe_phv_in_data_447,
  input  [7:0]  io_pipe_phv_in_data_448,
  input  [7:0]  io_pipe_phv_in_data_449,
  input  [7:0]  io_pipe_phv_in_data_450,
  input  [7:0]  io_pipe_phv_in_data_451,
  input  [7:0]  io_pipe_phv_in_data_452,
  input  [7:0]  io_pipe_phv_in_data_453,
  input  [7:0]  io_pipe_phv_in_data_454,
  input  [7:0]  io_pipe_phv_in_data_455,
  input  [7:0]  io_pipe_phv_in_data_456,
  input  [7:0]  io_pipe_phv_in_data_457,
  input  [7:0]  io_pipe_phv_in_data_458,
  input  [7:0]  io_pipe_phv_in_data_459,
  input  [7:0]  io_pipe_phv_in_data_460,
  input  [7:0]  io_pipe_phv_in_data_461,
  input  [7:0]  io_pipe_phv_in_data_462,
  input  [7:0]  io_pipe_phv_in_data_463,
  input  [7:0]  io_pipe_phv_in_data_464,
  input  [7:0]  io_pipe_phv_in_data_465,
  input  [7:0]  io_pipe_phv_in_data_466,
  input  [7:0]  io_pipe_phv_in_data_467,
  input  [7:0]  io_pipe_phv_in_data_468,
  input  [7:0]  io_pipe_phv_in_data_469,
  input  [7:0]  io_pipe_phv_in_data_470,
  input  [7:0]  io_pipe_phv_in_data_471,
  input  [7:0]  io_pipe_phv_in_data_472,
  input  [7:0]  io_pipe_phv_in_data_473,
  input  [7:0]  io_pipe_phv_in_data_474,
  input  [7:0]  io_pipe_phv_in_data_475,
  input  [7:0]  io_pipe_phv_in_data_476,
  input  [7:0]  io_pipe_phv_in_data_477,
  input  [7:0]  io_pipe_phv_in_data_478,
  input  [7:0]  io_pipe_phv_in_data_479,
  input  [7:0]  io_pipe_phv_in_data_480,
  input  [7:0]  io_pipe_phv_in_data_481,
  input  [7:0]  io_pipe_phv_in_data_482,
  input  [7:0]  io_pipe_phv_in_data_483,
  input  [7:0]  io_pipe_phv_in_data_484,
  input  [7:0]  io_pipe_phv_in_data_485,
  input  [7:0]  io_pipe_phv_in_data_486,
  input  [7:0]  io_pipe_phv_in_data_487,
  input  [7:0]  io_pipe_phv_in_data_488,
  input  [7:0]  io_pipe_phv_in_data_489,
  input  [7:0]  io_pipe_phv_in_data_490,
  input  [7:0]  io_pipe_phv_in_data_491,
  input  [7:0]  io_pipe_phv_in_data_492,
  input  [7:0]  io_pipe_phv_in_data_493,
  input  [7:0]  io_pipe_phv_in_data_494,
  input  [7:0]  io_pipe_phv_in_data_495,
  input  [7:0]  io_pipe_phv_in_data_496,
  input  [7:0]  io_pipe_phv_in_data_497,
  input  [7:0]  io_pipe_phv_in_data_498,
  input  [7:0]  io_pipe_phv_in_data_499,
  input  [7:0]  io_pipe_phv_in_data_500,
  input  [7:0]  io_pipe_phv_in_data_501,
  input  [7:0]  io_pipe_phv_in_data_502,
  input  [7:0]  io_pipe_phv_in_data_503,
  input  [7:0]  io_pipe_phv_in_data_504,
  input  [7:0]  io_pipe_phv_in_data_505,
  input  [7:0]  io_pipe_phv_in_data_506,
  input  [7:0]  io_pipe_phv_in_data_507,
  input  [7:0]  io_pipe_phv_in_data_508,
  input  [7:0]  io_pipe_phv_in_data_509,
  input  [7:0]  io_pipe_phv_in_data_510,
  input  [7:0]  io_pipe_phv_in_data_511,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [7:0]  io_pipe_phv_out_data_256,
  output [7:0]  io_pipe_phv_out_data_257,
  output [7:0]  io_pipe_phv_out_data_258,
  output [7:0]  io_pipe_phv_out_data_259,
  output [7:0]  io_pipe_phv_out_data_260,
  output [7:0]  io_pipe_phv_out_data_261,
  output [7:0]  io_pipe_phv_out_data_262,
  output [7:0]  io_pipe_phv_out_data_263,
  output [7:0]  io_pipe_phv_out_data_264,
  output [7:0]  io_pipe_phv_out_data_265,
  output [7:0]  io_pipe_phv_out_data_266,
  output [7:0]  io_pipe_phv_out_data_267,
  output [7:0]  io_pipe_phv_out_data_268,
  output [7:0]  io_pipe_phv_out_data_269,
  output [7:0]  io_pipe_phv_out_data_270,
  output [7:0]  io_pipe_phv_out_data_271,
  output [7:0]  io_pipe_phv_out_data_272,
  output [7:0]  io_pipe_phv_out_data_273,
  output [7:0]  io_pipe_phv_out_data_274,
  output [7:0]  io_pipe_phv_out_data_275,
  output [7:0]  io_pipe_phv_out_data_276,
  output [7:0]  io_pipe_phv_out_data_277,
  output [7:0]  io_pipe_phv_out_data_278,
  output [7:0]  io_pipe_phv_out_data_279,
  output [7:0]  io_pipe_phv_out_data_280,
  output [7:0]  io_pipe_phv_out_data_281,
  output [7:0]  io_pipe_phv_out_data_282,
  output [7:0]  io_pipe_phv_out_data_283,
  output [7:0]  io_pipe_phv_out_data_284,
  output [7:0]  io_pipe_phv_out_data_285,
  output [7:0]  io_pipe_phv_out_data_286,
  output [7:0]  io_pipe_phv_out_data_287,
  output [7:0]  io_pipe_phv_out_data_288,
  output [7:0]  io_pipe_phv_out_data_289,
  output [7:0]  io_pipe_phv_out_data_290,
  output [7:0]  io_pipe_phv_out_data_291,
  output [7:0]  io_pipe_phv_out_data_292,
  output [7:0]  io_pipe_phv_out_data_293,
  output [7:0]  io_pipe_phv_out_data_294,
  output [7:0]  io_pipe_phv_out_data_295,
  output [7:0]  io_pipe_phv_out_data_296,
  output [7:0]  io_pipe_phv_out_data_297,
  output [7:0]  io_pipe_phv_out_data_298,
  output [7:0]  io_pipe_phv_out_data_299,
  output [7:0]  io_pipe_phv_out_data_300,
  output [7:0]  io_pipe_phv_out_data_301,
  output [7:0]  io_pipe_phv_out_data_302,
  output [7:0]  io_pipe_phv_out_data_303,
  output [7:0]  io_pipe_phv_out_data_304,
  output [7:0]  io_pipe_phv_out_data_305,
  output [7:0]  io_pipe_phv_out_data_306,
  output [7:0]  io_pipe_phv_out_data_307,
  output [7:0]  io_pipe_phv_out_data_308,
  output [7:0]  io_pipe_phv_out_data_309,
  output [7:0]  io_pipe_phv_out_data_310,
  output [7:0]  io_pipe_phv_out_data_311,
  output [7:0]  io_pipe_phv_out_data_312,
  output [7:0]  io_pipe_phv_out_data_313,
  output [7:0]  io_pipe_phv_out_data_314,
  output [7:0]  io_pipe_phv_out_data_315,
  output [7:0]  io_pipe_phv_out_data_316,
  output [7:0]  io_pipe_phv_out_data_317,
  output [7:0]  io_pipe_phv_out_data_318,
  output [7:0]  io_pipe_phv_out_data_319,
  output [7:0]  io_pipe_phv_out_data_320,
  output [7:0]  io_pipe_phv_out_data_321,
  output [7:0]  io_pipe_phv_out_data_322,
  output [7:0]  io_pipe_phv_out_data_323,
  output [7:0]  io_pipe_phv_out_data_324,
  output [7:0]  io_pipe_phv_out_data_325,
  output [7:0]  io_pipe_phv_out_data_326,
  output [7:0]  io_pipe_phv_out_data_327,
  output [7:0]  io_pipe_phv_out_data_328,
  output [7:0]  io_pipe_phv_out_data_329,
  output [7:0]  io_pipe_phv_out_data_330,
  output [7:0]  io_pipe_phv_out_data_331,
  output [7:0]  io_pipe_phv_out_data_332,
  output [7:0]  io_pipe_phv_out_data_333,
  output [7:0]  io_pipe_phv_out_data_334,
  output [7:0]  io_pipe_phv_out_data_335,
  output [7:0]  io_pipe_phv_out_data_336,
  output [7:0]  io_pipe_phv_out_data_337,
  output [7:0]  io_pipe_phv_out_data_338,
  output [7:0]  io_pipe_phv_out_data_339,
  output [7:0]  io_pipe_phv_out_data_340,
  output [7:0]  io_pipe_phv_out_data_341,
  output [7:0]  io_pipe_phv_out_data_342,
  output [7:0]  io_pipe_phv_out_data_343,
  output [7:0]  io_pipe_phv_out_data_344,
  output [7:0]  io_pipe_phv_out_data_345,
  output [7:0]  io_pipe_phv_out_data_346,
  output [7:0]  io_pipe_phv_out_data_347,
  output [7:0]  io_pipe_phv_out_data_348,
  output [7:0]  io_pipe_phv_out_data_349,
  output [7:0]  io_pipe_phv_out_data_350,
  output [7:0]  io_pipe_phv_out_data_351,
  output [7:0]  io_pipe_phv_out_data_352,
  output [7:0]  io_pipe_phv_out_data_353,
  output [7:0]  io_pipe_phv_out_data_354,
  output [7:0]  io_pipe_phv_out_data_355,
  output [7:0]  io_pipe_phv_out_data_356,
  output [7:0]  io_pipe_phv_out_data_357,
  output [7:0]  io_pipe_phv_out_data_358,
  output [7:0]  io_pipe_phv_out_data_359,
  output [7:0]  io_pipe_phv_out_data_360,
  output [7:0]  io_pipe_phv_out_data_361,
  output [7:0]  io_pipe_phv_out_data_362,
  output [7:0]  io_pipe_phv_out_data_363,
  output [7:0]  io_pipe_phv_out_data_364,
  output [7:0]  io_pipe_phv_out_data_365,
  output [7:0]  io_pipe_phv_out_data_366,
  output [7:0]  io_pipe_phv_out_data_367,
  output [7:0]  io_pipe_phv_out_data_368,
  output [7:0]  io_pipe_phv_out_data_369,
  output [7:0]  io_pipe_phv_out_data_370,
  output [7:0]  io_pipe_phv_out_data_371,
  output [7:0]  io_pipe_phv_out_data_372,
  output [7:0]  io_pipe_phv_out_data_373,
  output [7:0]  io_pipe_phv_out_data_374,
  output [7:0]  io_pipe_phv_out_data_375,
  output [7:0]  io_pipe_phv_out_data_376,
  output [7:0]  io_pipe_phv_out_data_377,
  output [7:0]  io_pipe_phv_out_data_378,
  output [7:0]  io_pipe_phv_out_data_379,
  output [7:0]  io_pipe_phv_out_data_380,
  output [7:0]  io_pipe_phv_out_data_381,
  output [7:0]  io_pipe_phv_out_data_382,
  output [7:0]  io_pipe_phv_out_data_383,
  output [7:0]  io_pipe_phv_out_data_384,
  output [7:0]  io_pipe_phv_out_data_385,
  output [7:0]  io_pipe_phv_out_data_386,
  output [7:0]  io_pipe_phv_out_data_387,
  output [7:0]  io_pipe_phv_out_data_388,
  output [7:0]  io_pipe_phv_out_data_389,
  output [7:0]  io_pipe_phv_out_data_390,
  output [7:0]  io_pipe_phv_out_data_391,
  output [7:0]  io_pipe_phv_out_data_392,
  output [7:0]  io_pipe_phv_out_data_393,
  output [7:0]  io_pipe_phv_out_data_394,
  output [7:0]  io_pipe_phv_out_data_395,
  output [7:0]  io_pipe_phv_out_data_396,
  output [7:0]  io_pipe_phv_out_data_397,
  output [7:0]  io_pipe_phv_out_data_398,
  output [7:0]  io_pipe_phv_out_data_399,
  output [7:0]  io_pipe_phv_out_data_400,
  output [7:0]  io_pipe_phv_out_data_401,
  output [7:0]  io_pipe_phv_out_data_402,
  output [7:0]  io_pipe_phv_out_data_403,
  output [7:0]  io_pipe_phv_out_data_404,
  output [7:0]  io_pipe_phv_out_data_405,
  output [7:0]  io_pipe_phv_out_data_406,
  output [7:0]  io_pipe_phv_out_data_407,
  output [7:0]  io_pipe_phv_out_data_408,
  output [7:0]  io_pipe_phv_out_data_409,
  output [7:0]  io_pipe_phv_out_data_410,
  output [7:0]  io_pipe_phv_out_data_411,
  output [7:0]  io_pipe_phv_out_data_412,
  output [7:0]  io_pipe_phv_out_data_413,
  output [7:0]  io_pipe_phv_out_data_414,
  output [7:0]  io_pipe_phv_out_data_415,
  output [7:0]  io_pipe_phv_out_data_416,
  output [7:0]  io_pipe_phv_out_data_417,
  output [7:0]  io_pipe_phv_out_data_418,
  output [7:0]  io_pipe_phv_out_data_419,
  output [7:0]  io_pipe_phv_out_data_420,
  output [7:0]  io_pipe_phv_out_data_421,
  output [7:0]  io_pipe_phv_out_data_422,
  output [7:0]  io_pipe_phv_out_data_423,
  output [7:0]  io_pipe_phv_out_data_424,
  output [7:0]  io_pipe_phv_out_data_425,
  output [7:0]  io_pipe_phv_out_data_426,
  output [7:0]  io_pipe_phv_out_data_427,
  output [7:0]  io_pipe_phv_out_data_428,
  output [7:0]  io_pipe_phv_out_data_429,
  output [7:0]  io_pipe_phv_out_data_430,
  output [7:0]  io_pipe_phv_out_data_431,
  output [7:0]  io_pipe_phv_out_data_432,
  output [7:0]  io_pipe_phv_out_data_433,
  output [7:0]  io_pipe_phv_out_data_434,
  output [7:0]  io_pipe_phv_out_data_435,
  output [7:0]  io_pipe_phv_out_data_436,
  output [7:0]  io_pipe_phv_out_data_437,
  output [7:0]  io_pipe_phv_out_data_438,
  output [7:0]  io_pipe_phv_out_data_439,
  output [7:0]  io_pipe_phv_out_data_440,
  output [7:0]  io_pipe_phv_out_data_441,
  output [7:0]  io_pipe_phv_out_data_442,
  output [7:0]  io_pipe_phv_out_data_443,
  output [7:0]  io_pipe_phv_out_data_444,
  output [7:0]  io_pipe_phv_out_data_445,
  output [7:0]  io_pipe_phv_out_data_446,
  output [7:0]  io_pipe_phv_out_data_447,
  output [7:0]  io_pipe_phv_out_data_448,
  output [7:0]  io_pipe_phv_out_data_449,
  output [7:0]  io_pipe_phv_out_data_450,
  output [7:0]  io_pipe_phv_out_data_451,
  output [7:0]  io_pipe_phv_out_data_452,
  output [7:0]  io_pipe_phv_out_data_453,
  output [7:0]  io_pipe_phv_out_data_454,
  output [7:0]  io_pipe_phv_out_data_455,
  output [7:0]  io_pipe_phv_out_data_456,
  output [7:0]  io_pipe_phv_out_data_457,
  output [7:0]  io_pipe_phv_out_data_458,
  output [7:0]  io_pipe_phv_out_data_459,
  output [7:0]  io_pipe_phv_out_data_460,
  output [7:0]  io_pipe_phv_out_data_461,
  output [7:0]  io_pipe_phv_out_data_462,
  output [7:0]  io_pipe_phv_out_data_463,
  output [7:0]  io_pipe_phv_out_data_464,
  output [7:0]  io_pipe_phv_out_data_465,
  output [7:0]  io_pipe_phv_out_data_466,
  output [7:0]  io_pipe_phv_out_data_467,
  output [7:0]  io_pipe_phv_out_data_468,
  output [7:0]  io_pipe_phv_out_data_469,
  output [7:0]  io_pipe_phv_out_data_470,
  output [7:0]  io_pipe_phv_out_data_471,
  output [7:0]  io_pipe_phv_out_data_472,
  output [7:0]  io_pipe_phv_out_data_473,
  output [7:0]  io_pipe_phv_out_data_474,
  output [7:0]  io_pipe_phv_out_data_475,
  output [7:0]  io_pipe_phv_out_data_476,
  output [7:0]  io_pipe_phv_out_data_477,
  output [7:0]  io_pipe_phv_out_data_478,
  output [7:0]  io_pipe_phv_out_data_479,
  output [7:0]  io_pipe_phv_out_data_480,
  output [7:0]  io_pipe_phv_out_data_481,
  output [7:0]  io_pipe_phv_out_data_482,
  output [7:0]  io_pipe_phv_out_data_483,
  output [7:0]  io_pipe_phv_out_data_484,
  output [7:0]  io_pipe_phv_out_data_485,
  output [7:0]  io_pipe_phv_out_data_486,
  output [7:0]  io_pipe_phv_out_data_487,
  output [7:0]  io_pipe_phv_out_data_488,
  output [7:0]  io_pipe_phv_out_data_489,
  output [7:0]  io_pipe_phv_out_data_490,
  output [7:0]  io_pipe_phv_out_data_491,
  output [7:0]  io_pipe_phv_out_data_492,
  output [7:0]  io_pipe_phv_out_data_493,
  output [7:0]  io_pipe_phv_out_data_494,
  output [7:0]  io_pipe_phv_out_data_495,
  output [7:0]  io_pipe_phv_out_data_496,
  output [7:0]  io_pipe_phv_out_data_497,
  output [7:0]  io_pipe_phv_out_data_498,
  output [7:0]  io_pipe_phv_out_data_499,
  output [7:0]  io_pipe_phv_out_data_500,
  output [7:0]  io_pipe_phv_out_data_501,
  output [7:0]  io_pipe_phv_out_data_502,
  output [7:0]  io_pipe_phv_out_data_503,
  output [7:0]  io_pipe_phv_out_data_504,
  output [7:0]  io_pipe_phv_out_data_505,
  output [7:0]  io_pipe_phv_out_data_506,
  output [7:0]  io_pipe_phv_out_data_507,
  output [7:0]  io_pipe_phv_out_data_508,
  output [7:0]  io_pipe_phv_out_data_509,
  output [7:0]  io_pipe_phv_out_data_510,
  output [7:0]  io_pipe_phv_out_data_511,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  input         io_mod_par_mod_en,
  input         io_mod_par_mod_last_mau_id_mod,
  input  [1:0]  io_mod_par_mod_last_mau_id,
  input  [1:0]  io_mod_par_mod_cs,
  input         io_mod_par_mod_module_mod_state_id_mod,
  input  [7:0]  io_mod_par_mod_module_mod_state_id,
  input         io_mod_par_mod_module_mod_sram_w_cs,
  input         io_mod_par_mod_module_mod_sram_w_en,
  input  [7:0]  io_mod_par_mod_module_mod_sram_w_addr,
  input  [63:0] io_mod_par_mod_module_mod_sram_w_data,
  input         io_mod_mat_mod_en,
  input         io_mod_mat_mod_config_id,
  input  [7:0]  io_mod_mat_mod_key_mod_header_id,
  input  [7:0]  io_mod_mat_mod_key_mod_internal_offset,
  input  [7:0]  io_mod_mat_mod_key_mod_key_length,
  input  [4:0]  io_mod_mat_mod_table_mod_table_width,
  input  [4:0]  io_mod_mat_mod_table_mod_table_depth,
  input         io_mod_act_mod_en_0,
  input         io_mod_act_mod_en_1,
  input  [7:0]  io_mod_act_mod_addr,
  input  [63:0] io_mod_act_mod_data_0,
  input  [63:0] io_mod_act_mod_data_1,
  output        io_mem_cluster_0_en,
  output [7:0]  io_mem_cluster_0_addr,
  input  [63:0] io_mem_cluster_0_data,
  output        io_mem_cluster_1_en,
  output [7:0]  io_mem_cluster_1_addr,
  input  [63:0] io_mem_cluster_1_data,
  output        io_mem_cluster_2_en,
  output [7:0]  io_mem_cluster_2_addr,
  input  [63:0] io_mem_cluster_2_data,
  output        io_mem_cluster_3_en,
  output [7:0]  io_mem_cluster_3_addr,
  input  [63:0] io_mem_cluster_3_data,
  output        io_mem_cluster_4_en,
  output [7:0]  io_mem_cluster_4_addr,
  input  [63:0] io_mem_cluster_4_data,
  output        io_mem_cluster_5_en,
  output [7:0]  io_mem_cluster_5_addr,
  input  [63:0] io_mem_cluster_5_data,
  output        io_mem_cluster_6_en,
  output [7:0]  io_mem_cluster_6_addr,
  input  [63:0] io_mem_cluster_6_data,
  output        io_mem_cluster_7_en,
  output [7:0]  io_mem_cluster_7_addr,
  input  [63:0] io_mem_cluster_7_data,
  output        io_mem_cluster_8_en,
  output [7:0]  io_mem_cluster_8_addr,
  input  [63:0] io_mem_cluster_8_data,
  output        io_mem_cluster_9_en,
  output [7:0]  io_mem_cluster_9_addr,
  input  [63:0] io_mem_cluster_9_data,
  output        io_mem_cluster_10_en,
  output [7:0]  io_mem_cluster_10_addr,
  input  [63:0] io_mem_cluster_10_data,
  output        io_mem_cluster_11_en,
  output [7:0]  io_mem_cluster_11_addr,
  input  [63:0] io_mem_cluster_11_data,
  output        io_mem_cluster_12_en,
  output [7:0]  io_mem_cluster_12_addr,
  input  [63:0] io_mem_cluster_12_data,
  output        io_mem_cluster_13_en,
  output [7:0]  io_mem_cluster_13_addr,
  input  [63:0] io_mem_cluster_13_data,
  output        io_mem_cluster_14_en,
  output [7:0]  io_mem_cluster_14_addr,
  input  [63:0] io_mem_cluster_14_data,
  output        io_mem_cluster_15_en,
  output [7:0]  io_mem_cluster_15_addr,
  input  [63:0] io_mem_cluster_15_data
);
  wire  PAR_clock; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_0; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_1; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_2; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_3; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_4; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_5; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_6; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_7; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_8; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_9; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_10; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_11; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_12; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_13; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_14; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_15; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_16; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_17; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_18; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_19; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_20; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_21; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_22; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_23; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_24; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_25; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_26; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_27; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_28; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_29; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_30; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_31; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_32; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_33; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_34; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_35; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_36; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_37; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_38; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_39; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_40; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_41; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_42; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_43; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_44; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_45; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_46; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_47; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_48; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_49; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_50; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_51; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_52; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_53; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_54; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_55; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_56; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_57; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_58; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_59; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_60; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_61; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_62; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_63; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_64; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_65; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_66; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_67; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_68; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_69; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_70; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_71; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_72; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_73; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_74; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_75; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_76; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_77; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_78; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_79; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_80; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_81; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_82; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_83; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_84; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_85; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_86; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_87; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_88; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_89; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_90; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_91; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_92; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_93; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_94; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_95; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_96; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_97; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_98; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_99; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_100; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_101; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_102; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_103; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_104; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_105; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_106; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_107; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_108; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_109; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_110; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_111; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_112; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_113; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_114; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_115; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_116; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_117; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_118; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_119; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_120; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_121; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_122; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_123; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_124; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_125; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_126; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_127; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_128; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_129; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_130; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_131; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_132; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_133; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_134; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_135; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_136; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_137; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_138; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_139; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_140; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_141; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_142; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_143; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_144; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_145; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_146; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_147; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_148; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_149; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_150; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_151; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_152; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_153; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_154; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_155; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_156; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_157; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_158; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_159; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_160; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_161; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_162; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_163; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_164; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_165; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_166; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_167; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_168; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_169; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_170; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_171; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_172; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_173; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_174; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_175; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_176; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_177; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_178; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_179; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_180; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_181; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_182; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_183; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_184; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_185; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_186; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_187; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_188; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_189; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_190; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_191; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_192; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_193; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_194; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_195; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_196; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_197; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_198; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_199; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_200; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_201; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_202; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_203; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_204; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_205; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_206; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_207; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_208; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_209; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_210; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_211; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_212; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_213; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_214; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_215; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_216; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_217; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_218; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_219; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_220; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_221; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_222; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_223; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_224; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_225; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_226; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_227; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_228; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_229; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_230; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_231; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_232; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_233; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_234; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_235; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_236; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_237; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_238; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_239; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_240; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_241; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_242; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_243; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_244; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_245; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_246; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_247; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_248; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_249; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_250; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_251; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_252; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_253; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_254; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_255; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_256; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_257; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_258; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_259; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_260; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_261; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_262; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_263; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_264; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_265; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_266; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_267; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_268; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_269; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_270; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_271; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_272; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_273; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_274; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_275; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_276; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_277; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_278; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_279; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_280; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_281; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_282; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_283; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_284; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_285; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_286; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_287; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_288; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_289; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_290; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_291; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_292; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_293; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_294; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_295; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_296; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_297; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_298; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_299; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_300; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_301; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_302; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_303; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_304; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_305; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_306; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_307; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_308; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_309; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_310; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_311; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_312; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_313; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_314; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_315; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_316; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_317; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_318; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_319; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_320; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_321; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_322; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_323; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_324; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_325; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_326; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_327; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_328; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_329; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_330; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_331; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_332; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_333; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_334; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_335; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_336; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_337; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_338; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_339; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_340; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_341; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_342; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_343; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_344; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_345; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_346; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_347; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_348; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_349; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_350; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_351; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_352; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_353; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_354; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_355; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_356; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_357; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_358; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_359; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_360; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_361; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_362; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_363; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_364; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_365; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_366; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_367; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_368; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_369; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_370; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_371; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_372; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_373; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_374; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_375; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_376; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_377; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_378; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_379; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_380; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_381; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_382; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_383; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_384; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_385; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_386; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_387; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_388; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_389; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_390; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_391; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_392; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_393; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_394; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_395; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_396; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_397; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_398; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_399; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_400; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_401; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_402; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_403; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_404; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_405; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_406; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_407; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_408; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_409; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_410; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_411; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_412; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_413; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_414; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_415; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_416; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_417; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_418; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_419; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_420; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_421; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_422; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_423; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_424; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_425; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_426; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_427; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_428; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_429; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_430; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_431; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_432; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_433; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_434; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_435; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_436; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_437; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_438; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_439; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_440; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_441; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_442; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_443; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_444; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_445; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_446; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_447; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_448; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_449; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_450; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_451; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_452; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_453; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_454; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_455; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_456; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_457; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_458; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_459; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_460; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_461; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_462; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_463; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_464; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_465; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_466; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_467; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_468; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_469; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_470; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_471; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_472; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_473; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_474; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_475; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_476; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_477; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_478; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_479; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_480; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_481; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_482; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_483; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_484; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_485; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_486; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_487; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_488; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_489; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_490; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_491; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_492; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_493; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_494; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_495; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_496; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_497; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_498; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_499; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_500; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_501; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_502; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_503; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_504; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_505; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_506; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_507; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_508; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_509; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_510; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_511; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_0; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_1; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_2; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_3; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_4; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_5; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_6; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_7; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_8; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_9; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_10; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_11; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_12; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_13; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_14; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_15; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_parse_current_state; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_parse_current_offset; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_parse_transition_field; // @[processor.scala 13:21]
  wire [3:0] PAR_io_pipe_phv_in_next_processor_id; // @[processor.scala 13:21]
  wire  PAR_io_pipe_phv_in_next_config_id; // @[processor.scala 13:21]
  wire  PAR_io_pipe_phv_in_is_valid_processor; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_0; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_1; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_2; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_3; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_4; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_5; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_6; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_7; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_8; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_9; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_10; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_11; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_12; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_13; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_14; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_15; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_16; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_17; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_18; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_19; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_20; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_21; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_22; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_23; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_24; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_25; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_26; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_27; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_28; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_29; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_30; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_31; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_32; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_33; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_34; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_35; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_36; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_37; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_38; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_39; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_40; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_41; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_42; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_43; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_44; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_45; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_46; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_47; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_48; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_49; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_50; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_51; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_52; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_53; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_54; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_55; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_56; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_57; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_58; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_59; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_60; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_61; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_62; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_63; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_64; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_65; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_66; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_67; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_68; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_69; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_70; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_71; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_72; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_73; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_74; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_75; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_76; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_77; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_78; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_79; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_80; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_81; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_82; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_83; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_84; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_85; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_86; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_87; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_88; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_89; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_90; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_91; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_92; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_93; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_94; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_95; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_96; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_97; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_98; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_99; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_100; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_101; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_102; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_103; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_104; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_105; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_106; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_107; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_108; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_109; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_110; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_111; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_112; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_113; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_114; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_115; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_116; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_117; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_118; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_119; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_120; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_121; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_122; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_123; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_124; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_125; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_126; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_127; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_128; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_129; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_130; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_131; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_132; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_133; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_134; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_135; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_136; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_137; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_138; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_139; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_140; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_141; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_142; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_143; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_144; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_145; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_146; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_147; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_148; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_149; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_150; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_151; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_152; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_153; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_154; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_155; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_156; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_157; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_158; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_159; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_160; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_161; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_162; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_163; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_164; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_165; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_166; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_167; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_168; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_169; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_170; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_171; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_172; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_173; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_174; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_175; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_176; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_177; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_178; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_179; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_180; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_181; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_182; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_183; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_184; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_185; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_186; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_187; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_188; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_189; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_190; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_191; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_192; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_193; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_194; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_195; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_196; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_197; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_198; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_199; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_200; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_201; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_202; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_203; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_204; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_205; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_206; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_207; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_208; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_209; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_210; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_211; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_212; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_213; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_214; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_215; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_216; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_217; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_218; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_219; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_220; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_221; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_222; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_223; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_224; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_225; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_226; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_227; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_228; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_229; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_230; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_231; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_232; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_233; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_234; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_235; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_236; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_237; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_238; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_239; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_240; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_241; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_242; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_243; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_244; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_245; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_246; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_247; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_248; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_249; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_250; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_251; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_252; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_253; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_254; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_255; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_256; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_257; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_258; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_259; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_260; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_261; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_262; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_263; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_264; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_265; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_266; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_267; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_268; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_269; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_270; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_271; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_272; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_273; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_274; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_275; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_276; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_277; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_278; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_279; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_280; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_281; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_282; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_283; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_284; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_285; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_286; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_287; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_288; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_289; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_290; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_291; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_292; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_293; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_294; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_295; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_296; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_297; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_298; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_299; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_300; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_301; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_302; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_303; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_304; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_305; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_306; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_307; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_308; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_309; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_310; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_311; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_312; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_313; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_314; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_315; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_316; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_317; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_318; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_319; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_320; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_321; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_322; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_323; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_324; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_325; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_326; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_327; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_328; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_329; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_330; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_331; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_332; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_333; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_334; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_335; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_336; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_337; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_338; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_339; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_340; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_341; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_342; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_343; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_344; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_345; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_346; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_347; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_348; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_349; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_350; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_351; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_352; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_353; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_354; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_355; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_356; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_357; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_358; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_359; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_360; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_361; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_362; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_363; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_364; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_365; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_366; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_367; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_368; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_369; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_370; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_371; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_372; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_373; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_374; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_375; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_376; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_377; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_378; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_379; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_380; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_381; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_382; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_383; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_384; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_385; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_386; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_387; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_388; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_389; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_390; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_391; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_392; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_393; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_394; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_395; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_396; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_397; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_398; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_399; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_400; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_401; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_402; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_403; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_404; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_405; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_406; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_407; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_408; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_409; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_410; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_411; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_412; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_413; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_414; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_415; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_416; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_417; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_418; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_419; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_420; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_421; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_422; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_423; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_424; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_425; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_426; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_427; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_428; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_429; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_430; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_431; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_432; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_433; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_434; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_435; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_436; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_437; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_438; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_439; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_440; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_441; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_442; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_443; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_444; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_445; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_446; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_447; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_448; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_449; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_450; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_451; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_452; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_453; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_454; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_455; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_456; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_457; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_458; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_459; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_460; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_461; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_462; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_463; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_464; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_465; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_466; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_467; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_468; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_469; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_470; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_471; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_472; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_473; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_474; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_475; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_476; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_477; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_478; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_479; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_480; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_481; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_482; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_483; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_484; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_485; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_486; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_487; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_488; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_489; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_490; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_491; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_492; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_493; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_494; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_495; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_496; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_497; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_498; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_499; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_500; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_501; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_502; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_503; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_504; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_505; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_506; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_507; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_508; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_509; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_510; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_511; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_0; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_1; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_2; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_3; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_4; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_5; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_6; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_7; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_8; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_9; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_10; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_11; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_12; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_13; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_14; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_15; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_parse_current_state; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_parse_current_offset; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_parse_transition_field; // @[processor.scala 13:21]
  wire [3:0] PAR_io_pipe_phv_out_next_processor_id; // @[processor.scala 13:21]
  wire  PAR_io_pipe_phv_out_next_config_id; // @[processor.scala 13:21]
  wire  PAR_io_pipe_phv_out_is_valid_processor; // @[processor.scala 13:21]
  wire  PAR_io_mod_en; // @[processor.scala 13:21]
  wire  PAR_io_mod_last_mau_id_mod; // @[processor.scala 13:21]
  wire [1:0] PAR_io_mod_last_mau_id; // @[processor.scala 13:21]
  wire [1:0] PAR_io_mod_cs; // @[processor.scala 13:21]
  wire  PAR_io_mod_module_mod_state_id_mod; // @[processor.scala 13:21]
  wire [7:0] PAR_io_mod_module_mod_state_id; // @[processor.scala 13:21]
  wire  PAR_io_mod_module_mod_sram_w_cs; // @[processor.scala 13:21]
  wire  PAR_io_mod_module_mod_sram_w_en; // @[processor.scala 13:21]
  wire [7:0] PAR_io_mod_module_mod_sram_w_addr; // @[processor.scala 13:21]
  wire [63:0] PAR_io_mod_module_mod_sram_w_data; // @[processor.scala 13:21]
  wire  MAT_clock; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_0; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_1; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_2; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_3; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_4; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_5; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_6; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_7; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_8; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_9; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_10; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_11; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_12; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_13; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_14; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_15; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_16; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_17; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_18; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_19; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_20; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_21; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_22; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_23; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_24; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_25; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_26; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_27; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_28; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_29; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_30; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_31; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_32; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_33; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_34; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_35; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_36; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_37; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_38; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_39; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_40; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_41; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_42; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_43; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_44; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_45; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_46; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_47; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_48; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_49; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_50; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_51; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_52; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_53; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_54; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_55; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_56; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_57; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_58; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_59; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_60; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_61; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_62; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_63; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_64; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_65; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_66; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_67; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_68; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_69; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_70; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_71; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_72; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_73; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_74; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_75; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_76; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_77; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_78; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_79; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_80; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_81; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_82; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_83; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_84; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_85; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_86; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_87; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_88; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_89; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_90; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_91; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_92; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_93; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_94; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_95; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_96; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_97; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_98; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_99; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_100; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_101; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_102; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_103; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_104; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_105; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_106; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_107; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_108; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_109; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_110; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_111; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_112; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_113; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_114; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_115; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_116; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_117; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_118; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_119; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_120; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_121; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_122; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_123; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_124; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_125; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_126; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_127; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_128; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_129; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_130; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_131; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_132; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_133; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_134; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_135; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_136; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_137; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_138; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_139; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_140; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_141; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_142; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_143; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_144; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_145; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_146; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_147; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_148; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_149; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_150; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_151; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_152; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_153; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_154; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_155; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_156; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_157; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_158; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_159; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_160; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_161; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_162; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_163; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_164; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_165; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_166; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_167; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_168; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_169; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_170; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_171; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_172; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_173; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_174; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_175; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_176; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_177; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_178; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_179; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_180; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_181; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_182; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_183; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_184; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_185; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_186; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_187; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_188; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_189; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_190; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_191; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_192; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_193; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_194; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_195; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_196; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_197; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_198; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_199; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_200; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_201; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_202; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_203; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_204; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_205; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_206; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_207; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_208; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_209; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_210; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_211; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_212; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_213; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_214; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_215; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_216; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_217; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_218; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_219; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_220; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_221; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_222; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_223; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_224; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_225; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_226; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_227; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_228; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_229; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_230; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_231; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_232; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_233; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_234; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_235; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_236; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_237; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_238; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_239; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_240; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_241; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_242; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_243; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_244; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_245; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_246; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_247; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_248; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_249; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_250; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_251; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_252; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_253; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_254; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_255; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_256; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_257; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_258; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_259; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_260; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_261; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_262; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_263; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_264; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_265; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_266; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_267; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_268; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_269; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_270; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_271; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_272; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_273; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_274; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_275; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_276; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_277; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_278; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_279; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_280; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_281; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_282; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_283; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_284; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_285; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_286; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_287; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_288; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_289; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_290; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_291; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_292; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_293; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_294; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_295; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_296; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_297; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_298; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_299; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_300; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_301; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_302; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_303; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_304; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_305; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_306; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_307; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_308; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_309; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_310; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_311; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_312; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_313; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_314; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_315; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_316; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_317; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_318; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_319; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_320; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_321; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_322; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_323; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_324; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_325; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_326; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_327; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_328; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_329; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_330; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_331; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_332; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_333; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_334; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_335; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_336; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_337; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_338; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_339; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_340; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_341; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_342; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_343; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_344; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_345; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_346; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_347; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_348; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_349; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_350; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_351; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_352; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_353; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_354; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_355; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_356; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_357; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_358; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_359; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_360; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_361; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_362; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_363; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_364; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_365; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_366; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_367; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_368; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_369; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_370; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_371; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_372; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_373; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_374; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_375; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_376; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_377; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_378; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_379; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_380; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_381; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_382; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_383; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_384; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_385; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_386; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_387; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_388; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_389; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_390; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_391; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_392; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_393; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_394; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_395; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_396; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_397; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_398; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_399; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_400; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_401; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_402; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_403; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_404; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_405; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_406; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_407; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_408; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_409; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_410; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_411; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_412; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_413; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_414; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_415; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_416; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_417; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_418; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_419; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_420; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_421; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_422; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_423; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_424; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_425; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_426; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_427; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_428; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_429; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_430; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_431; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_432; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_433; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_434; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_435; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_436; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_437; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_438; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_439; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_440; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_441; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_442; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_443; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_444; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_445; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_446; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_447; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_448; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_449; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_450; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_451; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_452; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_453; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_454; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_455; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_456; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_457; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_458; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_459; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_460; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_461; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_462; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_463; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_464; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_465; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_466; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_467; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_468; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_469; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_470; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_471; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_472; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_473; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_474; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_475; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_476; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_477; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_478; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_479; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_480; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_481; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_482; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_483; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_484; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_485; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_486; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_487; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_488; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_489; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_490; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_491; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_492; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_493; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_494; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_495; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_496; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_497; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_498; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_499; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_500; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_501; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_502; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_503; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_504; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_505; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_506; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_507; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_508; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_509; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_510; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_511; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_0; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_1; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_2; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_3; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_4; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_5; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_6; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_7; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_8; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_9; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_10; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_11; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_12; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_13; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_14; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_15; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_parse_current_state; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_parse_current_offset; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_parse_transition_field; // @[processor.scala 14:21]
  wire [3:0] MAT_io_pipe_phv_in_next_processor_id; // @[processor.scala 14:21]
  wire  MAT_io_pipe_phv_in_next_config_id; // @[processor.scala 14:21]
  wire  MAT_io_pipe_phv_in_is_valid_processor; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_0; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_1; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_2; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_3; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_4; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_5; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_6; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_7; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_8; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_9; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_10; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_11; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_12; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_13; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_14; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_15; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_16; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_17; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_18; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_19; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_20; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_21; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_22; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_23; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_24; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_25; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_26; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_27; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_28; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_29; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_30; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_31; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_32; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_33; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_34; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_35; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_36; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_37; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_38; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_39; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_40; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_41; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_42; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_43; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_44; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_45; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_46; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_47; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_48; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_49; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_50; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_51; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_52; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_53; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_54; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_55; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_56; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_57; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_58; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_59; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_60; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_61; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_62; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_63; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_64; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_65; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_66; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_67; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_68; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_69; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_70; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_71; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_72; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_73; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_74; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_75; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_76; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_77; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_78; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_79; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_80; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_81; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_82; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_83; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_84; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_85; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_86; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_87; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_88; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_89; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_90; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_91; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_92; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_93; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_94; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_95; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_96; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_97; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_98; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_99; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_100; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_101; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_102; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_103; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_104; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_105; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_106; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_107; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_108; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_109; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_110; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_111; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_112; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_113; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_114; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_115; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_116; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_117; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_118; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_119; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_120; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_121; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_122; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_123; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_124; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_125; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_126; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_127; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_128; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_129; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_130; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_131; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_132; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_133; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_134; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_135; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_136; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_137; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_138; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_139; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_140; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_141; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_142; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_143; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_144; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_145; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_146; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_147; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_148; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_149; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_150; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_151; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_152; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_153; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_154; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_155; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_156; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_157; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_158; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_159; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_160; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_161; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_162; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_163; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_164; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_165; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_166; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_167; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_168; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_169; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_170; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_171; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_172; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_173; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_174; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_175; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_176; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_177; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_178; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_179; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_180; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_181; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_182; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_183; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_184; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_185; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_186; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_187; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_188; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_189; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_190; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_191; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_192; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_193; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_194; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_195; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_196; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_197; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_198; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_199; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_200; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_201; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_202; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_203; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_204; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_205; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_206; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_207; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_208; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_209; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_210; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_211; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_212; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_213; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_214; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_215; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_216; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_217; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_218; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_219; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_220; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_221; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_222; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_223; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_224; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_225; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_226; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_227; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_228; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_229; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_230; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_231; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_232; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_233; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_234; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_235; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_236; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_237; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_238; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_239; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_240; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_241; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_242; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_243; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_244; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_245; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_246; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_247; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_248; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_249; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_250; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_251; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_252; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_253; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_254; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_255; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_256; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_257; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_258; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_259; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_260; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_261; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_262; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_263; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_264; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_265; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_266; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_267; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_268; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_269; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_270; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_271; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_272; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_273; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_274; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_275; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_276; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_277; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_278; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_279; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_280; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_281; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_282; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_283; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_284; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_285; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_286; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_287; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_288; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_289; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_290; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_291; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_292; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_293; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_294; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_295; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_296; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_297; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_298; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_299; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_300; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_301; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_302; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_303; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_304; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_305; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_306; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_307; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_308; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_309; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_310; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_311; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_312; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_313; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_314; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_315; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_316; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_317; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_318; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_319; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_320; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_321; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_322; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_323; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_324; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_325; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_326; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_327; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_328; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_329; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_330; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_331; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_332; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_333; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_334; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_335; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_336; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_337; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_338; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_339; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_340; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_341; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_342; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_343; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_344; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_345; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_346; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_347; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_348; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_349; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_350; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_351; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_352; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_353; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_354; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_355; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_356; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_357; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_358; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_359; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_360; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_361; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_362; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_363; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_364; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_365; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_366; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_367; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_368; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_369; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_370; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_371; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_372; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_373; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_374; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_375; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_376; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_377; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_378; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_379; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_380; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_381; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_382; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_383; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_384; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_385; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_386; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_387; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_388; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_389; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_390; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_391; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_392; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_393; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_394; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_395; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_396; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_397; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_398; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_399; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_400; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_401; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_402; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_403; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_404; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_405; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_406; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_407; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_408; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_409; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_410; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_411; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_412; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_413; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_414; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_415; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_416; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_417; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_418; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_419; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_420; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_421; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_422; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_423; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_424; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_425; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_426; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_427; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_428; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_429; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_430; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_431; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_432; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_433; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_434; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_435; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_436; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_437; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_438; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_439; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_440; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_441; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_442; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_443; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_444; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_445; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_446; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_447; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_448; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_449; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_450; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_451; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_452; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_453; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_454; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_455; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_456; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_457; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_458; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_459; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_460; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_461; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_462; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_463; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_464; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_465; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_466; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_467; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_468; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_469; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_470; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_471; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_472; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_473; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_474; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_475; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_476; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_477; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_478; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_479; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_480; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_481; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_482; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_483; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_484; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_485; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_486; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_487; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_488; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_489; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_490; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_491; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_492; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_493; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_494; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_495; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_496; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_497; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_498; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_499; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_500; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_501; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_502; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_503; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_504; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_505; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_506; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_507; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_508; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_509; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_510; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_511; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_0; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_1; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_2; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_3; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_4; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_5; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_6; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_7; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_8; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_9; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_10; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_11; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_12; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_13; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_14; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_15; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_parse_current_state; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_parse_current_offset; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_parse_transition_field; // @[processor.scala 14:21]
  wire [3:0] MAT_io_pipe_phv_out_next_processor_id; // @[processor.scala 14:21]
  wire  MAT_io_pipe_phv_out_next_config_id; // @[processor.scala 14:21]
  wire  MAT_io_pipe_phv_out_is_valid_processor; // @[processor.scala 14:21]
  wire  MAT_io_mod_en; // @[processor.scala 14:21]
  wire  MAT_io_mod_config_id; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mod_key_mod_header_id; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mod_key_mod_internal_offset; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mod_key_mod_key_length; // @[processor.scala 14:21]
  wire [4:0] MAT_io_mod_table_mod_table_width; // @[processor.scala 14:21]
  wire [4:0] MAT_io_mod_table_mod_table_depth; // @[processor.scala 14:21]
  wire  MAT_io_hit; // @[processor.scala 14:21]
  wire [63:0] MAT_io_match_value; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_0_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_0_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_0_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_1_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_1_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_1_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_2_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_2_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_2_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_3_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_3_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_3_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_4_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_4_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_4_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_5_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_5_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_5_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_6_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_6_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_6_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_7_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_7_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_7_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_8_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_8_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_8_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_9_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_9_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_9_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_10_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_10_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_10_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_11_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_11_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_11_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_12_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_12_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_12_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_13_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_13_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_13_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_14_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_14_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_14_data; // @[processor.scala 14:21]
  wire  MAT_io_mem_cluster_15_en; // @[processor.scala 14:21]
  wire [7:0] MAT_io_mem_cluster_15_addr; // @[processor.scala 14:21]
  wire [63:0] MAT_io_mem_cluster_15_data; // @[processor.scala 14:21]
  wire  EXE_clock; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_0; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_1; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_2; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_3; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_4; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_5; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_6; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_7; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_8; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_9; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_10; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_11; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_12; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_13; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_14; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_15; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_16; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_17; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_18; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_19; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_20; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_21; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_22; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_23; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_24; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_25; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_26; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_27; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_28; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_29; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_30; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_31; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_32; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_33; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_34; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_35; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_36; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_37; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_38; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_39; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_40; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_41; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_42; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_43; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_44; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_45; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_46; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_47; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_48; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_49; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_50; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_51; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_52; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_53; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_54; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_55; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_56; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_57; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_58; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_59; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_60; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_61; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_62; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_63; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_64; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_65; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_66; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_67; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_68; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_69; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_70; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_71; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_72; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_73; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_74; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_75; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_76; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_77; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_78; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_79; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_80; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_81; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_82; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_83; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_84; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_85; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_86; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_87; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_88; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_89; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_90; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_91; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_92; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_93; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_94; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_95; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_96; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_97; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_98; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_99; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_100; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_101; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_102; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_103; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_104; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_105; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_106; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_107; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_108; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_109; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_110; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_111; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_112; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_113; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_114; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_115; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_116; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_117; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_118; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_119; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_120; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_121; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_122; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_123; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_124; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_125; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_126; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_127; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_128; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_129; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_130; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_131; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_132; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_133; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_134; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_135; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_136; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_137; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_138; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_139; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_140; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_141; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_142; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_143; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_144; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_145; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_146; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_147; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_148; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_149; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_150; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_151; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_152; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_153; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_154; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_155; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_156; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_157; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_158; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_159; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_160; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_161; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_162; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_163; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_164; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_165; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_166; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_167; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_168; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_169; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_170; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_171; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_172; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_173; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_174; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_175; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_176; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_177; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_178; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_179; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_180; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_181; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_182; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_183; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_184; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_185; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_186; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_187; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_188; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_189; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_190; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_191; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_192; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_193; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_194; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_195; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_196; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_197; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_198; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_199; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_200; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_201; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_202; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_203; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_204; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_205; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_206; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_207; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_208; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_209; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_210; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_211; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_212; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_213; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_214; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_215; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_216; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_217; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_218; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_219; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_220; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_221; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_222; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_223; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_224; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_225; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_226; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_227; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_228; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_229; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_230; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_231; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_232; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_233; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_234; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_235; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_236; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_237; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_238; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_239; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_240; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_241; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_242; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_243; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_244; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_245; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_246; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_247; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_248; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_249; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_250; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_251; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_252; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_253; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_254; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_255; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_256; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_257; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_258; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_259; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_260; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_261; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_262; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_263; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_264; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_265; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_266; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_267; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_268; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_269; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_270; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_271; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_272; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_273; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_274; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_275; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_276; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_277; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_278; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_279; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_280; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_281; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_282; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_283; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_284; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_285; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_286; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_287; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_288; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_289; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_290; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_291; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_292; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_293; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_294; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_295; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_296; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_297; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_298; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_299; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_300; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_301; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_302; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_303; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_304; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_305; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_306; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_307; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_308; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_309; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_310; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_311; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_312; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_313; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_314; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_315; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_316; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_317; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_318; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_319; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_320; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_321; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_322; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_323; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_324; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_325; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_326; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_327; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_328; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_329; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_330; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_331; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_332; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_333; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_334; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_335; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_336; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_337; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_338; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_339; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_340; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_341; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_342; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_343; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_344; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_345; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_346; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_347; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_348; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_349; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_350; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_351; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_352; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_353; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_354; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_355; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_356; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_357; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_358; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_359; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_360; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_361; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_362; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_363; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_364; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_365; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_366; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_367; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_368; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_369; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_370; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_371; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_372; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_373; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_374; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_375; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_376; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_377; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_378; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_379; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_380; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_381; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_382; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_383; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_384; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_385; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_386; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_387; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_388; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_389; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_390; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_391; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_392; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_393; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_394; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_395; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_396; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_397; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_398; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_399; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_400; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_401; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_402; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_403; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_404; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_405; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_406; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_407; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_408; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_409; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_410; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_411; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_412; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_413; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_414; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_415; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_416; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_417; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_418; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_419; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_420; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_421; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_422; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_423; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_424; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_425; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_426; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_427; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_428; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_429; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_430; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_431; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_432; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_433; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_434; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_435; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_436; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_437; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_438; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_439; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_440; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_441; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_442; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_443; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_444; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_445; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_446; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_447; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_448; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_449; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_450; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_451; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_452; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_453; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_454; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_455; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_456; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_457; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_458; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_459; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_460; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_461; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_462; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_463; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_464; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_465; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_466; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_467; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_468; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_469; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_470; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_471; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_472; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_473; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_474; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_475; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_476; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_477; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_478; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_479; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_480; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_481; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_482; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_483; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_484; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_485; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_486; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_487; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_488; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_489; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_490; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_491; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_492; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_493; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_494; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_495; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_496; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_497; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_498; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_499; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_500; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_501; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_502; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_503; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_504; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_505; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_506; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_507; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_508; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_509; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_510; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_511; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_0; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_1; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_2; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_3; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_4; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_5; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_6; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_7; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_8; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_9; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_10; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_11; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_12; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_13; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_14; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_15; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_parse_current_state; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_parse_current_offset; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_parse_transition_field; // @[processor.scala 15:21]
  wire [3:0] EXE_io_pipe_phv_in_next_processor_id; // @[processor.scala 15:21]
  wire  EXE_io_pipe_phv_in_next_config_id; // @[processor.scala 15:21]
  wire  EXE_io_pipe_phv_in_is_valid_processor; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_0; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_1; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_2; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_3; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_4; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_5; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_6; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_7; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_8; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_9; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_10; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_11; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_12; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_13; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_14; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_15; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_16; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_17; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_18; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_19; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_20; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_21; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_22; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_23; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_24; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_25; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_26; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_27; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_28; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_29; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_30; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_31; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_32; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_33; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_34; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_35; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_36; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_37; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_38; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_39; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_40; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_41; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_42; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_43; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_44; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_45; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_46; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_47; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_48; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_49; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_50; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_51; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_52; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_53; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_54; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_55; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_56; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_57; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_58; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_59; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_60; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_61; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_62; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_63; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_64; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_65; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_66; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_67; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_68; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_69; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_70; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_71; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_72; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_73; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_74; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_75; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_76; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_77; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_78; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_79; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_80; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_81; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_82; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_83; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_84; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_85; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_86; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_87; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_88; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_89; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_90; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_91; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_92; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_93; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_94; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_95; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_96; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_97; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_98; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_99; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_100; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_101; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_102; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_103; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_104; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_105; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_106; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_107; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_108; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_109; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_110; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_111; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_112; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_113; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_114; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_115; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_116; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_117; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_118; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_119; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_120; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_121; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_122; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_123; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_124; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_125; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_126; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_127; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_128; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_129; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_130; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_131; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_132; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_133; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_134; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_135; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_136; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_137; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_138; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_139; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_140; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_141; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_142; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_143; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_144; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_145; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_146; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_147; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_148; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_149; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_150; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_151; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_152; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_153; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_154; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_155; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_156; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_157; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_158; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_159; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_160; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_161; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_162; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_163; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_164; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_165; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_166; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_167; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_168; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_169; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_170; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_171; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_172; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_173; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_174; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_175; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_176; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_177; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_178; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_179; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_180; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_181; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_182; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_183; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_184; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_185; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_186; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_187; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_188; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_189; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_190; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_191; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_192; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_193; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_194; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_195; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_196; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_197; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_198; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_199; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_200; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_201; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_202; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_203; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_204; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_205; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_206; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_207; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_208; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_209; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_210; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_211; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_212; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_213; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_214; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_215; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_216; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_217; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_218; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_219; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_220; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_221; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_222; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_223; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_224; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_225; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_226; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_227; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_228; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_229; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_230; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_231; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_232; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_233; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_234; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_235; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_236; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_237; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_238; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_239; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_240; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_241; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_242; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_243; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_244; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_245; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_246; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_247; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_248; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_249; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_250; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_251; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_252; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_253; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_254; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_255; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_256; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_257; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_258; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_259; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_260; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_261; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_262; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_263; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_264; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_265; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_266; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_267; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_268; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_269; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_270; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_271; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_272; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_273; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_274; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_275; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_276; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_277; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_278; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_279; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_280; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_281; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_282; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_283; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_284; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_285; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_286; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_287; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_288; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_289; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_290; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_291; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_292; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_293; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_294; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_295; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_296; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_297; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_298; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_299; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_300; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_301; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_302; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_303; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_304; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_305; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_306; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_307; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_308; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_309; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_310; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_311; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_312; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_313; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_314; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_315; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_316; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_317; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_318; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_319; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_320; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_321; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_322; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_323; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_324; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_325; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_326; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_327; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_328; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_329; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_330; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_331; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_332; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_333; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_334; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_335; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_336; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_337; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_338; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_339; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_340; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_341; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_342; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_343; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_344; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_345; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_346; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_347; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_348; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_349; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_350; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_351; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_352; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_353; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_354; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_355; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_356; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_357; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_358; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_359; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_360; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_361; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_362; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_363; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_364; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_365; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_366; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_367; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_368; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_369; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_370; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_371; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_372; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_373; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_374; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_375; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_376; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_377; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_378; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_379; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_380; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_381; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_382; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_383; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_384; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_385; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_386; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_387; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_388; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_389; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_390; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_391; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_392; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_393; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_394; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_395; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_396; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_397; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_398; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_399; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_400; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_401; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_402; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_403; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_404; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_405; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_406; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_407; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_408; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_409; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_410; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_411; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_412; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_413; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_414; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_415; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_416; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_417; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_418; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_419; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_420; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_421; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_422; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_423; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_424; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_425; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_426; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_427; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_428; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_429; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_430; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_431; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_432; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_433; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_434; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_435; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_436; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_437; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_438; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_439; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_440; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_441; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_442; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_443; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_444; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_445; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_446; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_447; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_448; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_449; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_450; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_451; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_452; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_453; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_454; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_455; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_456; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_457; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_458; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_459; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_460; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_461; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_462; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_463; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_464; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_465; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_466; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_467; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_468; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_469; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_470; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_471; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_472; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_473; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_474; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_475; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_476; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_477; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_478; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_479; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_480; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_481; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_482; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_483; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_484; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_485; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_486; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_487; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_488; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_489; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_490; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_491; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_492; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_493; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_494; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_495; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_496; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_497; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_498; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_499; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_500; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_501; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_502; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_503; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_504; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_505; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_506; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_507; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_508; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_509; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_510; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_511; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_0; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_1; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_2; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_3; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_4; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_5; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_6; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_7; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_8; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_9; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_10; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_11; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_12; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_13; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_14; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_15; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_parse_current_state; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_parse_current_offset; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_parse_transition_field; // @[processor.scala 15:21]
  wire [3:0] EXE_io_pipe_phv_out_next_processor_id; // @[processor.scala 15:21]
  wire  EXE_io_pipe_phv_out_next_config_id; // @[processor.scala 15:21]
  wire  EXE_io_hit; // @[processor.scala 15:21]
  wire [63:0] EXE_io_match_value; // @[processor.scala 15:21]
  wire  EXE_io_action_mod_en_0; // @[processor.scala 15:21]
  wire  EXE_io_action_mod_en_1; // @[processor.scala 15:21]
  wire [7:0] EXE_io_action_mod_addr; // @[processor.scala 15:21]
  wire [63:0] EXE_io_action_mod_data_0; // @[processor.scala 15:21]
  wire [63:0] EXE_io_action_mod_data_1; // @[processor.scala 15:21]
  Parser PAR ( // @[processor.scala 13:21]
    .clock(PAR_clock),
    .io_pipe_phv_in_data_0(PAR_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(PAR_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(PAR_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(PAR_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(PAR_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(PAR_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(PAR_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(PAR_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(PAR_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(PAR_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(PAR_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(PAR_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(PAR_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(PAR_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(PAR_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(PAR_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(PAR_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(PAR_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(PAR_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(PAR_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(PAR_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(PAR_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(PAR_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(PAR_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(PAR_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(PAR_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(PAR_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(PAR_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(PAR_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(PAR_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(PAR_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(PAR_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(PAR_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(PAR_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(PAR_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(PAR_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(PAR_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(PAR_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(PAR_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(PAR_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(PAR_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(PAR_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(PAR_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(PAR_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(PAR_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(PAR_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(PAR_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(PAR_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(PAR_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(PAR_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(PAR_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(PAR_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(PAR_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(PAR_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(PAR_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(PAR_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(PAR_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(PAR_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(PAR_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(PAR_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(PAR_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(PAR_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(PAR_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(PAR_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(PAR_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(PAR_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(PAR_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(PAR_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(PAR_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(PAR_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(PAR_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(PAR_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(PAR_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(PAR_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(PAR_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(PAR_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(PAR_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(PAR_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(PAR_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(PAR_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(PAR_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(PAR_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(PAR_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(PAR_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(PAR_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(PAR_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(PAR_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(PAR_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(PAR_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(PAR_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(PAR_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(PAR_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(PAR_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(PAR_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(PAR_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(PAR_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(PAR_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(PAR_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(PAR_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(PAR_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(PAR_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(PAR_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(PAR_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(PAR_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(PAR_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(PAR_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(PAR_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(PAR_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(PAR_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(PAR_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(PAR_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(PAR_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(PAR_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(PAR_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(PAR_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(PAR_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(PAR_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(PAR_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(PAR_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(PAR_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(PAR_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(PAR_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(PAR_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(PAR_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(PAR_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(PAR_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(PAR_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(PAR_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(PAR_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(PAR_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(PAR_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(PAR_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(PAR_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(PAR_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(PAR_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(PAR_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(PAR_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(PAR_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(PAR_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(PAR_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(PAR_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(PAR_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(PAR_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(PAR_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(PAR_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(PAR_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(PAR_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(PAR_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(PAR_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(PAR_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(PAR_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(PAR_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(PAR_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(PAR_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(PAR_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(PAR_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(PAR_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(PAR_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(PAR_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(PAR_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(PAR_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(PAR_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(PAR_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(PAR_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(PAR_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(PAR_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(PAR_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(PAR_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(PAR_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(PAR_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(PAR_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(PAR_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(PAR_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(PAR_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(PAR_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(PAR_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(PAR_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(PAR_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(PAR_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(PAR_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(PAR_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(PAR_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(PAR_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(PAR_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(PAR_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(PAR_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(PAR_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(PAR_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(PAR_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(PAR_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(PAR_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(PAR_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(PAR_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(PAR_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(PAR_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(PAR_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(PAR_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(PAR_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(PAR_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(PAR_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(PAR_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(PAR_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(PAR_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(PAR_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(PAR_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(PAR_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(PAR_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(PAR_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(PAR_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(PAR_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(PAR_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(PAR_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(PAR_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(PAR_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(PAR_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(PAR_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(PAR_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(PAR_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(PAR_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(PAR_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(PAR_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(PAR_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(PAR_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(PAR_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(PAR_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(PAR_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(PAR_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(PAR_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(PAR_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(PAR_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(PAR_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(PAR_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(PAR_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(PAR_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(PAR_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(PAR_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(PAR_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(PAR_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(PAR_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(PAR_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(PAR_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(PAR_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(PAR_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(PAR_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(PAR_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(PAR_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(PAR_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(PAR_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(PAR_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(PAR_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(PAR_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(PAR_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(PAR_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(PAR_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(PAR_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(PAR_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(PAR_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(PAR_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(PAR_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(PAR_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(PAR_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(PAR_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(PAR_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(PAR_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(PAR_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(PAR_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(PAR_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(PAR_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(PAR_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(PAR_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(PAR_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(PAR_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(PAR_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(PAR_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(PAR_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(PAR_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(PAR_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(PAR_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(PAR_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(PAR_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(PAR_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(PAR_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(PAR_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(PAR_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(PAR_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(PAR_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(PAR_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(PAR_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(PAR_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(PAR_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(PAR_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(PAR_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(PAR_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(PAR_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(PAR_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(PAR_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(PAR_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(PAR_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(PAR_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(PAR_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(PAR_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(PAR_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(PAR_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(PAR_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(PAR_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(PAR_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(PAR_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(PAR_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(PAR_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(PAR_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(PAR_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(PAR_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(PAR_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(PAR_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(PAR_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(PAR_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(PAR_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(PAR_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(PAR_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(PAR_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(PAR_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(PAR_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(PAR_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(PAR_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(PAR_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(PAR_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(PAR_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(PAR_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(PAR_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(PAR_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(PAR_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(PAR_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(PAR_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(PAR_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(PAR_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(PAR_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(PAR_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(PAR_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(PAR_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(PAR_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(PAR_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(PAR_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(PAR_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(PAR_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(PAR_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(PAR_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(PAR_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(PAR_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(PAR_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(PAR_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(PAR_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(PAR_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(PAR_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(PAR_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(PAR_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(PAR_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(PAR_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(PAR_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(PAR_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(PAR_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(PAR_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(PAR_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(PAR_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(PAR_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(PAR_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(PAR_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(PAR_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(PAR_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(PAR_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(PAR_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(PAR_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(PAR_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(PAR_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(PAR_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(PAR_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(PAR_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(PAR_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(PAR_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(PAR_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(PAR_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(PAR_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(PAR_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(PAR_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(PAR_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(PAR_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(PAR_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(PAR_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(PAR_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(PAR_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(PAR_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(PAR_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(PAR_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(PAR_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(PAR_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(PAR_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(PAR_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(PAR_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(PAR_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(PAR_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(PAR_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(PAR_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(PAR_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(PAR_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(PAR_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(PAR_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(PAR_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(PAR_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(PAR_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(PAR_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(PAR_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(PAR_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(PAR_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(PAR_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(PAR_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(PAR_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(PAR_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(PAR_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(PAR_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(PAR_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(PAR_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(PAR_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(PAR_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(PAR_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(PAR_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(PAR_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(PAR_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(PAR_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(PAR_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(PAR_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(PAR_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(PAR_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(PAR_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(PAR_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(PAR_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(PAR_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(PAR_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(PAR_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(PAR_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(PAR_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(PAR_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(PAR_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(PAR_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(PAR_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(PAR_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(PAR_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(PAR_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(PAR_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(PAR_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(PAR_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(PAR_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(PAR_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(PAR_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(PAR_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(PAR_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(PAR_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(PAR_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(PAR_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(PAR_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(PAR_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(PAR_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(PAR_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(PAR_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(PAR_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(PAR_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(PAR_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(PAR_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(PAR_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(PAR_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(PAR_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(PAR_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(PAR_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(PAR_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(PAR_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(PAR_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(PAR_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(PAR_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(PAR_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(PAR_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(PAR_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(PAR_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(PAR_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(PAR_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(PAR_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(PAR_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(PAR_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(PAR_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(PAR_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(PAR_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(PAR_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(PAR_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(PAR_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(PAR_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(PAR_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(PAR_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(PAR_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(PAR_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(PAR_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(PAR_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(PAR_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(PAR_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(PAR_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(PAR_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(PAR_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(PAR_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(PAR_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(PAR_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(PAR_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(PAR_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(PAR_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(PAR_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(PAR_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(PAR_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(PAR_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(PAR_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(PAR_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(PAR_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(PAR_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(PAR_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(PAR_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(PAR_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(PAR_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(PAR_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(PAR_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(PAR_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(PAR_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(PAR_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(PAR_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(PAR_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(PAR_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(PAR_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(PAR_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(PAR_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(PAR_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(PAR_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(PAR_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(PAR_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(PAR_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(PAR_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(PAR_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(PAR_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(PAR_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(PAR_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(PAR_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(PAR_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(PAR_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(PAR_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(PAR_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(PAR_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(PAR_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(PAR_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(PAR_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(PAR_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(PAR_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(PAR_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(PAR_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(PAR_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(PAR_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(PAR_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(PAR_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(PAR_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(PAR_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(PAR_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(PAR_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(PAR_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(PAR_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(PAR_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(PAR_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(PAR_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(PAR_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(PAR_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(PAR_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(PAR_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(PAR_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(PAR_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(PAR_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(PAR_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(PAR_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(PAR_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(PAR_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(PAR_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(PAR_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(PAR_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(PAR_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(PAR_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(PAR_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(PAR_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(PAR_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(PAR_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(PAR_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(PAR_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(PAR_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(PAR_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(PAR_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(PAR_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(PAR_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(PAR_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(PAR_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(PAR_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(PAR_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(PAR_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(PAR_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(PAR_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(PAR_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(PAR_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(PAR_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(PAR_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(PAR_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(PAR_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(PAR_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(PAR_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(PAR_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(PAR_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(PAR_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(PAR_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(PAR_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(PAR_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(PAR_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(PAR_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(PAR_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(PAR_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(PAR_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(PAR_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(PAR_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(PAR_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(PAR_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(PAR_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(PAR_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(PAR_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(PAR_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(PAR_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(PAR_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(PAR_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(PAR_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(PAR_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(PAR_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(PAR_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(PAR_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(PAR_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(PAR_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(PAR_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(PAR_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(PAR_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(PAR_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(PAR_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(PAR_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(PAR_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(PAR_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(PAR_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(PAR_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(PAR_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(PAR_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(PAR_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(PAR_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(PAR_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(PAR_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(PAR_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(PAR_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(PAR_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(PAR_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(PAR_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(PAR_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(PAR_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(PAR_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(PAR_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(PAR_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(PAR_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(PAR_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(PAR_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(PAR_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(PAR_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(PAR_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(PAR_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(PAR_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(PAR_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(PAR_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(PAR_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(PAR_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(PAR_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(PAR_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(PAR_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(PAR_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(PAR_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(PAR_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(PAR_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(PAR_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(PAR_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(PAR_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(PAR_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(PAR_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(PAR_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(PAR_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(PAR_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(PAR_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(PAR_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(PAR_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(PAR_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(PAR_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(PAR_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(PAR_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(PAR_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(PAR_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(PAR_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(PAR_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(PAR_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(PAR_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(PAR_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(PAR_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(PAR_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(PAR_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(PAR_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(PAR_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(PAR_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(PAR_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(PAR_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(PAR_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(PAR_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(PAR_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(PAR_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(PAR_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(PAR_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(PAR_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(PAR_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(PAR_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(PAR_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(PAR_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(PAR_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(PAR_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(PAR_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(PAR_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(PAR_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(PAR_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(PAR_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(PAR_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(PAR_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(PAR_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(PAR_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(PAR_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(PAR_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(PAR_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(PAR_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(PAR_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(PAR_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(PAR_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(PAR_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(PAR_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(PAR_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(PAR_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(PAR_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(PAR_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(PAR_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(PAR_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(PAR_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(PAR_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(PAR_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(PAR_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(PAR_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(PAR_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(PAR_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(PAR_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(PAR_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(PAR_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(PAR_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(PAR_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(PAR_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(PAR_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(PAR_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(PAR_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(PAR_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(PAR_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(PAR_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(PAR_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(PAR_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(PAR_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(PAR_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(PAR_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(PAR_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(PAR_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(PAR_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(PAR_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(PAR_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(PAR_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(PAR_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(PAR_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(PAR_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(PAR_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(PAR_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(PAR_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(PAR_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(PAR_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(PAR_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(PAR_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(PAR_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(PAR_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(PAR_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(PAR_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(PAR_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(PAR_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(PAR_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(PAR_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(PAR_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(PAR_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(PAR_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(PAR_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(PAR_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(PAR_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(PAR_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(PAR_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(PAR_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(PAR_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(PAR_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(PAR_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(PAR_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(PAR_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(PAR_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(PAR_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(PAR_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(PAR_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(PAR_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(PAR_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(PAR_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(PAR_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(PAR_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(PAR_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(PAR_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(PAR_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(PAR_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(PAR_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(PAR_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(PAR_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(PAR_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(PAR_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(PAR_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(PAR_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(PAR_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(PAR_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(PAR_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(PAR_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(PAR_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(PAR_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(PAR_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(PAR_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(PAR_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(PAR_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(PAR_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(PAR_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(PAR_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(PAR_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(PAR_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(PAR_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(PAR_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(PAR_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(PAR_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(PAR_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(PAR_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(PAR_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(PAR_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(PAR_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(PAR_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(PAR_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(PAR_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(PAR_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(PAR_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(PAR_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(PAR_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(PAR_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(PAR_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(PAR_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(PAR_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(PAR_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(PAR_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(PAR_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(PAR_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(PAR_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(PAR_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(PAR_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(PAR_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(PAR_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(PAR_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(PAR_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(PAR_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(PAR_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(PAR_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(PAR_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(PAR_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(PAR_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(PAR_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(PAR_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(PAR_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(PAR_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(PAR_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(PAR_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(PAR_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(PAR_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(PAR_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(PAR_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(PAR_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(PAR_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(PAR_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(PAR_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(PAR_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(PAR_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(PAR_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(PAR_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(PAR_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(PAR_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(PAR_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(PAR_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(PAR_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(PAR_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(PAR_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(PAR_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(PAR_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(PAR_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(PAR_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(PAR_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(PAR_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(PAR_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(PAR_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(PAR_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(PAR_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(PAR_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(PAR_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(PAR_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(PAR_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(PAR_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(PAR_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(PAR_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(PAR_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(PAR_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(PAR_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(PAR_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(PAR_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(PAR_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(PAR_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(PAR_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(PAR_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(PAR_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(PAR_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(PAR_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(PAR_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(PAR_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(PAR_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(PAR_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(PAR_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(PAR_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(PAR_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(PAR_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(PAR_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(PAR_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(PAR_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(PAR_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(PAR_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(PAR_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(PAR_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(PAR_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(PAR_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(PAR_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(PAR_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(PAR_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(PAR_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(PAR_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(PAR_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(PAR_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(PAR_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(PAR_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(PAR_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(PAR_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(PAR_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(PAR_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(PAR_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(PAR_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(PAR_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(PAR_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(PAR_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(PAR_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(PAR_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(PAR_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(PAR_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(PAR_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(PAR_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(PAR_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(PAR_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(PAR_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(PAR_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(PAR_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(PAR_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(PAR_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(PAR_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(PAR_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(PAR_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(PAR_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(PAR_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(PAR_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(PAR_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(PAR_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(PAR_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(PAR_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(PAR_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(PAR_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(PAR_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(PAR_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(PAR_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(PAR_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(PAR_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(PAR_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(PAR_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(PAR_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(PAR_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(PAR_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(PAR_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(PAR_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(PAR_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(PAR_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(PAR_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(PAR_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(PAR_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(PAR_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(PAR_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(PAR_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(PAR_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(PAR_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(PAR_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(PAR_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(PAR_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(PAR_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(PAR_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(PAR_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(PAR_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(PAR_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(PAR_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(PAR_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(PAR_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(PAR_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(PAR_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(PAR_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(PAR_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(PAR_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(PAR_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(PAR_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(PAR_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(PAR_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(PAR_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(PAR_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(PAR_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(PAR_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(PAR_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(PAR_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(PAR_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(PAR_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(PAR_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(PAR_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(PAR_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(PAR_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(PAR_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(PAR_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(PAR_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(PAR_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(PAR_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(PAR_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(PAR_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(PAR_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(PAR_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(PAR_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(PAR_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(PAR_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(PAR_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(PAR_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(PAR_io_pipe_phv_out_is_valid_processor),
    .io_mod_en(PAR_io_mod_en),
    .io_mod_last_mau_id_mod(PAR_io_mod_last_mau_id_mod),
    .io_mod_last_mau_id(PAR_io_mod_last_mau_id),
    .io_mod_cs(PAR_io_mod_cs),
    .io_mod_module_mod_state_id_mod(PAR_io_mod_module_mod_state_id_mod),
    .io_mod_module_mod_state_id(PAR_io_mod_module_mod_state_id),
    .io_mod_module_mod_sram_w_cs(PAR_io_mod_module_mod_sram_w_cs),
    .io_mod_module_mod_sram_w_en(PAR_io_mod_module_mod_sram_w_en),
    .io_mod_module_mod_sram_w_addr(PAR_io_mod_module_mod_sram_w_addr),
    .io_mod_module_mod_sram_w_data(PAR_io_mod_module_mod_sram_w_data)
  );
  Matcher MAT ( // @[processor.scala 14:21]
    .clock(MAT_clock),
    .io_pipe_phv_in_data_0(MAT_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(MAT_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(MAT_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(MAT_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(MAT_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(MAT_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(MAT_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(MAT_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(MAT_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(MAT_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(MAT_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(MAT_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(MAT_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(MAT_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(MAT_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(MAT_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(MAT_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(MAT_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(MAT_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(MAT_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(MAT_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(MAT_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(MAT_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(MAT_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(MAT_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(MAT_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(MAT_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(MAT_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(MAT_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(MAT_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(MAT_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(MAT_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(MAT_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(MAT_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(MAT_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(MAT_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(MAT_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(MAT_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(MAT_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(MAT_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(MAT_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(MAT_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(MAT_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(MAT_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(MAT_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(MAT_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(MAT_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(MAT_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(MAT_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(MAT_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(MAT_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(MAT_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(MAT_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(MAT_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(MAT_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(MAT_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(MAT_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(MAT_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(MAT_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(MAT_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(MAT_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(MAT_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(MAT_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(MAT_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(MAT_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(MAT_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(MAT_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(MAT_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(MAT_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(MAT_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(MAT_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(MAT_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(MAT_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(MAT_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(MAT_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(MAT_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(MAT_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(MAT_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(MAT_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(MAT_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(MAT_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(MAT_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(MAT_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(MAT_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(MAT_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(MAT_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(MAT_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(MAT_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(MAT_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(MAT_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(MAT_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(MAT_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(MAT_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(MAT_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(MAT_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(MAT_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(MAT_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(MAT_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(MAT_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(MAT_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(MAT_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(MAT_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(MAT_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(MAT_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(MAT_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(MAT_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(MAT_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(MAT_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(MAT_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(MAT_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(MAT_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(MAT_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(MAT_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(MAT_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(MAT_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(MAT_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(MAT_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(MAT_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(MAT_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(MAT_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(MAT_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(MAT_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(MAT_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(MAT_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(MAT_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(MAT_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(MAT_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(MAT_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(MAT_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(MAT_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(MAT_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(MAT_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(MAT_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(MAT_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(MAT_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(MAT_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(MAT_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(MAT_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(MAT_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(MAT_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(MAT_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(MAT_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(MAT_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(MAT_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(MAT_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(MAT_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(MAT_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(MAT_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(MAT_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(MAT_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(MAT_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(MAT_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(MAT_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(MAT_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(MAT_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(MAT_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(MAT_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(MAT_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(MAT_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(MAT_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(MAT_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(MAT_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(MAT_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(MAT_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(MAT_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(MAT_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(MAT_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(MAT_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(MAT_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(MAT_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(MAT_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(MAT_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(MAT_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(MAT_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(MAT_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(MAT_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(MAT_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(MAT_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(MAT_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(MAT_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(MAT_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(MAT_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(MAT_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(MAT_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(MAT_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(MAT_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(MAT_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(MAT_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(MAT_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(MAT_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(MAT_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(MAT_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(MAT_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(MAT_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(MAT_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(MAT_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(MAT_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(MAT_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(MAT_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(MAT_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(MAT_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(MAT_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(MAT_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(MAT_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(MAT_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(MAT_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(MAT_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(MAT_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(MAT_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(MAT_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(MAT_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(MAT_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(MAT_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(MAT_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(MAT_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(MAT_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(MAT_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(MAT_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(MAT_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(MAT_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(MAT_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(MAT_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(MAT_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(MAT_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(MAT_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(MAT_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(MAT_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(MAT_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(MAT_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(MAT_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(MAT_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(MAT_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(MAT_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(MAT_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(MAT_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(MAT_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(MAT_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(MAT_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(MAT_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(MAT_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(MAT_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(MAT_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(MAT_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(MAT_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(MAT_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(MAT_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(MAT_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(MAT_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(MAT_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(MAT_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(MAT_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(MAT_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(MAT_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(MAT_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(MAT_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(MAT_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(MAT_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(MAT_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(MAT_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(MAT_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(MAT_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(MAT_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(MAT_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(MAT_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(MAT_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(MAT_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(MAT_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(MAT_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(MAT_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(MAT_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(MAT_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(MAT_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(MAT_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(MAT_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(MAT_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(MAT_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(MAT_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(MAT_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(MAT_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(MAT_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(MAT_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(MAT_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(MAT_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(MAT_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(MAT_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(MAT_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(MAT_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(MAT_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(MAT_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(MAT_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(MAT_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(MAT_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(MAT_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(MAT_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(MAT_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(MAT_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(MAT_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(MAT_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(MAT_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(MAT_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(MAT_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(MAT_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(MAT_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(MAT_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(MAT_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(MAT_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(MAT_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(MAT_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(MAT_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(MAT_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(MAT_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(MAT_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(MAT_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(MAT_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(MAT_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(MAT_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(MAT_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(MAT_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(MAT_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(MAT_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(MAT_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(MAT_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(MAT_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(MAT_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(MAT_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(MAT_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(MAT_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(MAT_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(MAT_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(MAT_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(MAT_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(MAT_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(MAT_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(MAT_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(MAT_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(MAT_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(MAT_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(MAT_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(MAT_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(MAT_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(MAT_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(MAT_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(MAT_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(MAT_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(MAT_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(MAT_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(MAT_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(MAT_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(MAT_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(MAT_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(MAT_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(MAT_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(MAT_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(MAT_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(MAT_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(MAT_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(MAT_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(MAT_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(MAT_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(MAT_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(MAT_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(MAT_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(MAT_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(MAT_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(MAT_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(MAT_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(MAT_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(MAT_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(MAT_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(MAT_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(MAT_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(MAT_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(MAT_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(MAT_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(MAT_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(MAT_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(MAT_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(MAT_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(MAT_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(MAT_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(MAT_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(MAT_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(MAT_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(MAT_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(MAT_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(MAT_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(MAT_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(MAT_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(MAT_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(MAT_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(MAT_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(MAT_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(MAT_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(MAT_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(MAT_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(MAT_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(MAT_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(MAT_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(MAT_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(MAT_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(MAT_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(MAT_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(MAT_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(MAT_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(MAT_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(MAT_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(MAT_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(MAT_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(MAT_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(MAT_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(MAT_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(MAT_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(MAT_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(MAT_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(MAT_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(MAT_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(MAT_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(MAT_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(MAT_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(MAT_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(MAT_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(MAT_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(MAT_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(MAT_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(MAT_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(MAT_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(MAT_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(MAT_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(MAT_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(MAT_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(MAT_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(MAT_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(MAT_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(MAT_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(MAT_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(MAT_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(MAT_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(MAT_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(MAT_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(MAT_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(MAT_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(MAT_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(MAT_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(MAT_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(MAT_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(MAT_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(MAT_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(MAT_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(MAT_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(MAT_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(MAT_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(MAT_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(MAT_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(MAT_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(MAT_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(MAT_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(MAT_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(MAT_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(MAT_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(MAT_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(MAT_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(MAT_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(MAT_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(MAT_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(MAT_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(MAT_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(MAT_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(MAT_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(MAT_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(MAT_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(MAT_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(MAT_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(MAT_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(MAT_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(MAT_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(MAT_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(MAT_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(MAT_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(MAT_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(MAT_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(MAT_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(MAT_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(MAT_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(MAT_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(MAT_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(MAT_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(MAT_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(MAT_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(MAT_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(MAT_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(MAT_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(MAT_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(MAT_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(MAT_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(MAT_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(MAT_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(MAT_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(MAT_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(MAT_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(MAT_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(MAT_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(MAT_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(MAT_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(MAT_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(MAT_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(MAT_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(MAT_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(MAT_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(MAT_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(MAT_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(MAT_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(MAT_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(MAT_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(MAT_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(MAT_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(MAT_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(MAT_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(MAT_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(MAT_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(MAT_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(MAT_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(MAT_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(MAT_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(MAT_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(MAT_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(MAT_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(MAT_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(MAT_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(MAT_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(MAT_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(MAT_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(MAT_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(MAT_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(MAT_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(MAT_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(MAT_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(MAT_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(MAT_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(MAT_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(MAT_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(MAT_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(MAT_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(MAT_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(MAT_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(MAT_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(MAT_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(MAT_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(MAT_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(MAT_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(MAT_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(MAT_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(MAT_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(MAT_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(MAT_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(MAT_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(MAT_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(MAT_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(MAT_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(MAT_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(MAT_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(MAT_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(MAT_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(MAT_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(MAT_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(MAT_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(MAT_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(MAT_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(MAT_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(MAT_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(MAT_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(MAT_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(MAT_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(MAT_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(MAT_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(MAT_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(MAT_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(MAT_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(MAT_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(MAT_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(MAT_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(MAT_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(MAT_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(MAT_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(MAT_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(MAT_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(MAT_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(MAT_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(MAT_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(MAT_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(MAT_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(MAT_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(MAT_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(MAT_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(MAT_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(MAT_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(MAT_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(MAT_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(MAT_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(MAT_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(MAT_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(MAT_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(MAT_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(MAT_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(MAT_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(MAT_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(MAT_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(MAT_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(MAT_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(MAT_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(MAT_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(MAT_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(MAT_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(MAT_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(MAT_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(MAT_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(MAT_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(MAT_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(MAT_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(MAT_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(MAT_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(MAT_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(MAT_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(MAT_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(MAT_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(MAT_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(MAT_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(MAT_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(MAT_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(MAT_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(MAT_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(MAT_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(MAT_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(MAT_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(MAT_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(MAT_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(MAT_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(MAT_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(MAT_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(MAT_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(MAT_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(MAT_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(MAT_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(MAT_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(MAT_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(MAT_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(MAT_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(MAT_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(MAT_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(MAT_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(MAT_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(MAT_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(MAT_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(MAT_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(MAT_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(MAT_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(MAT_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(MAT_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(MAT_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(MAT_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(MAT_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(MAT_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(MAT_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(MAT_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(MAT_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(MAT_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(MAT_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(MAT_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(MAT_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(MAT_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(MAT_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(MAT_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(MAT_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(MAT_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(MAT_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(MAT_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(MAT_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(MAT_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(MAT_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(MAT_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(MAT_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(MAT_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(MAT_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(MAT_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(MAT_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(MAT_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(MAT_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(MAT_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(MAT_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(MAT_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(MAT_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(MAT_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(MAT_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(MAT_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(MAT_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(MAT_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(MAT_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(MAT_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(MAT_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(MAT_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(MAT_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(MAT_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(MAT_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(MAT_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(MAT_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(MAT_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(MAT_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(MAT_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(MAT_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(MAT_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(MAT_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(MAT_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(MAT_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(MAT_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(MAT_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(MAT_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(MAT_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(MAT_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(MAT_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(MAT_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(MAT_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(MAT_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(MAT_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(MAT_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(MAT_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(MAT_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(MAT_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(MAT_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(MAT_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(MAT_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(MAT_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(MAT_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(MAT_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(MAT_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(MAT_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(MAT_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(MAT_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(MAT_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(MAT_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(MAT_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(MAT_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(MAT_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(MAT_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(MAT_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(MAT_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(MAT_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(MAT_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(MAT_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(MAT_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(MAT_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(MAT_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(MAT_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(MAT_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(MAT_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(MAT_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(MAT_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(MAT_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(MAT_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(MAT_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(MAT_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(MAT_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(MAT_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(MAT_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(MAT_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(MAT_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(MAT_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(MAT_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(MAT_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(MAT_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(MAT_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(MAT_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(MAT_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(MAT_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(MAT_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(MAT_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(MAT_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(MAT_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(MAT_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(MAT_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(MAT_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(MAT_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(MAT_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(MAT_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(MAT_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(MAT_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(MAT_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(MAT_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(MAT_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(MAT_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(MAT_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(MAT_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(MAT_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(MAT_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(MAT_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(MAT_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(MAT_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(MAT_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(MAT_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(MAT_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(MAT_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(MAT_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(MAT_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(MAT_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(MAT_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(MAT_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(MAT_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(MAT_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(MAT_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(MAT_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(MAT_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(MAT_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(MAT_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(MAT_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(MAT_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(MAT_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(MAT_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(MAT_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(MAT_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(MAT_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(MAT_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(MAT_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(MAT_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(MAT_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(MAT_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(MAT_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(MAT_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(MAT_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(MAT_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(MAT_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(MAT_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(MAT_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(MAT_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(MAT_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(MAT_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(MAT_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(MAT_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(MAT_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(MAT_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(MAT_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(MAT_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(MAT_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(MAT_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(MAT_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(MAT_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(MAT_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(MAT_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(MAT_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(MAT_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(MAT_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(MAT_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(MAT_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(MAT_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(MAT_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(MAT_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(MAT_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(MAT_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(MAT_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(MAT_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(MAT_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(MAT_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(MAT_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(MAT_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(MAT_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(MAT_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(MAT_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(MAT_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(MAT_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(MAT_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(MAT_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(MAT_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(MAT_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(MAT_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(MAT_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(MAT_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(MAT_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(MAT_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(MAT_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(MAT_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(MAT_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(MAT_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(MAT_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(MAT_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(MAT_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(MAT_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(MAT_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(MAT_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(MAT_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(MAT_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(MAT_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(MAT_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(MAT_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(MAT_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(MAT_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(MAT_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(MAT_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(MAT_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(MAT_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(MAT_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(MAT_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(MAT_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(MAT_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(MAT_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(MAT_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(MAT_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(MAT_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(MAT_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(MAT_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(MAT_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(MAT_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(MAT_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(MAT_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(MAT_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(MAT_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(MAT_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(MAT_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(MAT_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(MAT_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(MAT_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(MAT_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(MAT_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(MAT_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(MAT_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(MAT_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(MAT_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(MAT_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(MAT_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(MAT_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(MAT_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(MAT_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(MAT_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(MAT_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(MAT_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(MAT_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(MAT_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(MAT_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(MAT_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(MAT_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(MAT_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(MAT_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(MAT_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(MAT_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(MAT_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(MAT_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(MAT_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(MAT_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(MAT_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(MAT_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(MAT_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(MAT_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(MAT_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(MAT_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(MAT_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(MAT_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(MAT_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(MAT_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(MAT_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(MAT_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(MAT_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(MAT_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(MAT_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(MAT_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(MAT_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(MAT_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(MAT_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(MAT_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(MAT_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(MAT_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(MAT_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(MAT_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(MAT_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(MAT_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(MAT_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(MAT_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(MAT_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(MAT_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(MAT_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(MAT_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(MAT_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(MAT_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(MAT_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(MAT_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(MAT_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(MAT_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(MAT_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(MAT_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(MAT_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(MAT_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(MAT_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(MAT_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(MAT_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(MAT_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(MAT_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(MAT_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(MAT_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(MAT_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(MAT_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(MAT_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(MAT_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(MAT_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(MAT_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(MAT_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(MAT_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(MAT_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(MAT_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(MAT_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(MAT_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(MAT_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(MAT_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(MAT_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(MAT_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(MAT_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(MAT_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(MAT_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(MAT_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(MAT_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(MAT_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(MAT_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(MAT_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(MAT_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(MAT_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(MAT_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(MAT_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(MAT_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(MAT_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(MAT_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(MAT_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(MAT_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(MAT_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(MAT_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(MAT_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(MAT_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(MAT_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(MAT_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(MAT_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(MAT_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(MAT_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(MAT_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(MAT_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(MAT_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(MAT_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(MAT_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(MAT_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(MAT_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(MAT_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(MAT_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(MAT_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(MAT_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(MAT_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(MAT_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(MAT_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(MAT_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(MAT_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(MAT_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(MAT_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(MAT_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(MAT_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(MAT_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(MAT_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(MAT_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(MAT_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(MAT_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(MAT_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(MAT_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(MAT_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(MAT_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(MAT_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(MAT_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(MAT_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(MAT_io_pipe_phv_out_is_valid_processor),
    .io_mod_en(MAT_io_mod_en),
    .io_mod_config_id(MAT_io_mod_config_id),
    .io_mod_key_mod_header_id(MAT_io_mod_key_mod_header_id),
    .io_mod_key_mod_internal_offset(MAT_io_mod_key_mod_internal_offset),
    .io_mod_key_mod_key_length(MAT_io_mod_key_mod_key_length),
    .io_mod_table_mod_table_width(MAT_io_mod_table_mod_table_width),
    .io_mod_table_mod_table_depth(MAT_io_mod_table_mod_table_depth),
    .io_hit(MAT_io_hit),
    .io_match_value(MAT_io_match_value),
    .io_mem_cluster_0_en(MAT_io_mem_cluster_0_en),
    .io_mem_cluster_0_addr(MAT_io_mem_cluster_0_addr),
    .io_mem_cluster_0_data(MAT_io_mem_cluster_0_data),
    .io_mem_cluster_1_en(MAT_io_mem_cluster_1_en),
    .io_mem_cluster_1_addr(MAT_io_mem_cluster_1_addr),
    .io_mem_cluster_1_data(MAT_io_mem_cluster_1_data),
    .io_mem_cluster_2_en(MAT_io_mem_cluster_2_en),
    .io_mem_cluster_2_addr(MAT_io_mem_cluster_2_addr),
    .io_mem_cluster_2_data(MAT_io_mem_cluster_2_data),
    .io_mem_cluster_3_en(MAT_io_mem_cluster_3_en),
    .io_mem_cluster_3_addr(MAT_io_mem_cluster_3_addr),
    .io_mem_cluster_3_data(MAT_io_mem_cluster_3_data),
    .io_mem_cluster_4_en(MAT_io_mem_cluster_4_en),
    .io_mem_cluster_4_addr(MAT_io_mem_cluster_4_addr),
    .io_mem_cluster_4_data(MAT_io_mem_cluster_4_data),
    .io_mem_cluster_5_en(MAT_io_mem_cluster_5_en),
    .io_mem_cluster_5_addr(MAT_io_mem_cluster_5_addr),
    .io_mem_cluster_5_data(MAT_io_mem_cluster_5_data),
    .io_mem_cluster_6_en(MAT_io_mem_cluster_6_en),
    .io_mem_cluster_6_addr(MAT_io_mem_cluster_6_addr),
    .io_mem_cluster_6_data(MAT_io_mem_cluster_6_data),
    .io_mem_cluster_7_en(MAT_io_mem_cluster_7_en),
    .io_mem_cluster_7_addr(MAT_io_mem_cluster_7_addr),
    .io_mem_cluster_7_data(MAT_io_mem_cluster_7_data),
    .io_mem_cluster_8_en(MAT_io_mem_cluster_8_en),
    .io_mem_cluster_8_addr(MAT_io_mem_cluster_8_addr),
    .io_mem_cluster_8_data(MAT_io_mem_cluster_8_data),
    .io_mem_cluster_9_en(MAT_io_mem_cluster_9_en),
    .io_mem_cluster_9_addr(MAT_io_mem_cluster_9_addr),
    .io_mem_cluster_9_data(MAT_io_mem_cluster_9_data),
    .io_mem_cluster_10_en(MAT_io_mem_cluster_10_en),
    .io_mem_cluster_10_addr(MAT_io_mem_cluster_10_addr),
    .io_mem_cluster_10_data(MAT_io_mem_cluster_10_data),
    .io_mem_cluster_11_en(MAT_io_mem_cluster_11_en),
    .io_mem_cluster_11_addr(MAT_io_mem_cluster_11_addr),
    .io_mem_cluster_11_data(MAT_io_mem_cluster_11_data),
    .io_mem_cluster_12_en(MAT_io_mem_cluster_12_en),
    .io_mem_cluster_12_addr(MAT_io_mem_cluster_12_addr),
    .io_mem_cluster_12_data(MAT_io_mem_cluster_12_data),
    .io_mem_cluster_13_en(MAT_io_mem_cluster_13_en),
    .io_mem_cluster_13_addr(MAT_io_mem_cluster_13_addr),
    .io_mem_cluster_13_data(MAT_io_mem_cluster_13_data),
    .io_mem_cluster_14_en(MAT_io_mem_cluster_14_en),
    .io_mem_cluster_14_addr(MAT_io_mem_cluster_14_addr),
    .io_mem_cluster_14_data(MAT_io_mem_cluster_14_data),
    .io_mem_cluster_15_en(MAT_io_mem_cluster_15_en),
    .io_mem_cluster_15_addr(MAT_io_mem_cluster_15_addr),
    .io_mem_cluster_15_data(MAT_io_mem_cluster_15_data)
  );
  Executor EXE ( // @[processor.scala 15:21]
    .clock(EXE_clock),
    .io_pipe_phv_in_data_0(EXE_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(EXE_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(EXE_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(EXE_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(EXE_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(EXE_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(EXE_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(EXE_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(EXE_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(EXE_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(EXE_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(EXE_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(EXE_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(EXE_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(EXE_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(EXE_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(EXE_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(EXE_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(EXE_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(EXE_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(EXE_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(EXE_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(EXE_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(EXE_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(EXE_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(EXE_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(EXE_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(EXE_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(EXE_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(EXE_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(EXE_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(EXE_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(EXE_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(EXE_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(EXE_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(EXE_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(EXE_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(EXE_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(EXE_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(EXE_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(EXE_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(EXE_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(EXE_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(EXE_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(EXE_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(EXE_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(EXE_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(EXE_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(EXE_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(EXE_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(EXE_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(EXE_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(EXE_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(EXE_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(EXE_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(EXE_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(EXE_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(EXE_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(EXE_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(EXE_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(EXE_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(EXE_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(EXE_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(EXE_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(EXE_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(EXE_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(EXE_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(EXE_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(EXE_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(EXE_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(EXE_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(EXE_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(EXE_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(EXE_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(EXE_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(EXE_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(EXE_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(EXE_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(EXE_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(EXE_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(EXE_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(EXE_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(EXE_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(EXE_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(EXE_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(EXE_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(EXE_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(EXE_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(EXE_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(EXE_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(EXE_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(EXE_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(EXE_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(EXE_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(EXE_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(EXE_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(EXE_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(EXE_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(EXE_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(EXE_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(EXE_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(EXE_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(EXE_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(EXE_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(EXE_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(EXE_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(EXE_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(EXE_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(EXE_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(EXE_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(EXE_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(EXE_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(EXE_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(EXE_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(EXE_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(EXE_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(EXE_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(EXE_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(EXE_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(EXE_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(EXE_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(EXE_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(EXE_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(EXE_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(EXE_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(EXE_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(EXE_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(EXE_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(EXE_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(EXE_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(EXE_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(EXE_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(EXE_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(EXE_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(EXE_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(EXE_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(EXE_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(EXE_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(EXE_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(EXE_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(EXE_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(EXE_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(EXE_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(EXE_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(EXE_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(EXE_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(EXE_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(EXE_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(EXE_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(EXE_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(EXE_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(EXE_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(EXE_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(EXE_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(EXE_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(EXE_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(EXE_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(EXE_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(EXE_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(EXE_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(EXE_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(EXE_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(EXE_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(EXE_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(EXE_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(EXE_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(EXE_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(EXE_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(EXE_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(EXE_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(EXE_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(EXE_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(EXE_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(EXE_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(EXE_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(EXE_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(EXE_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(EXE_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(EXE_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(EXE_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(EXE_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(EXE_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(EXE_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(EXE_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(EXE_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(EXE_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(EXE_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(EXE_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(EXE_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(EXE_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(EXE_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(EXE_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(EXE_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(EXE_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(EXE_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(EXE_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(EXE_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(EXE_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(EXE_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(EXE_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(EXE_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(EXE_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(EXE_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(EXE_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(EXE_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(EXE_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(EXE_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(EXE_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(EXE_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(EXE_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(EXE_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(EXE_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(EXE_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(EXE_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(EXE_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(EXE_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(EXE_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(EXE_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(EXE_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(EXE_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(EXE_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(EXE_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(EXE_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(EXE_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(EXE_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(EXE_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(EXE_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(EXE_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(EXE_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(EXE_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(EXE_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(EXE_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(EXE_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(EXE_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(EXE_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(EXE_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(EXE_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(EXE_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(EXE_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(EXE_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(EXE_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(EXE_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(EXE_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(EXE_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(EXE_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(EXE_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(EXE_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(EXE_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(EXE_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(EXE_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(EXE_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(EXE_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(EXE_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(EXE_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(EXE_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(EXE_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(EXE_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(EXE_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(EXE_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(EXE_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(EXE_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(EXE_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(EXE_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(EXE_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(EXE_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(EXE_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(EXE_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(EXE_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(EXE_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(EXE_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(EXE_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(EXE_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(EXE_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(EXE_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(EXE_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(EXE_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(EXE_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(EXE_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(EXE_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(EXE_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(EXE_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(EXE_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(EXE_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(EXE_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(EXE_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(EXE_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(EXE_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(EXE_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(EXE_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(EXE_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(EXE_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(EXE_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(EXE_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(EXE_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(EXE_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(EXE_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(EXE_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(EXE_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(EXE_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(EXE_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(EXE_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(EXE_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(EXE_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(EXE_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(EXE_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(EXE_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(EXE_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(EXE_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(EXE_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(EXE_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(EXE_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(EXE_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(EXE_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(EXE_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(EXE_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(EXE_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(EXE_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(EXE_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(EXE_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(EXE_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(EXE_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(EXE_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(EXE_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(EXE_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(EXE_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(EXE_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(EXE_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(EXE_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(EXE_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(EXE_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(EXE_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(EXE_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(EXE_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(EXE_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(EXE_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(EXE_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(EXE_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(EXE_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(EXE_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(EXE_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(EXE_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(EXE_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(EXE_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(EXE_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(EXE_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(EXE_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(EXE_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(EXE_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(EXE_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(EXE_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(EXE_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(EXE_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(EXE_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(EXE_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(EXE_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(EXE_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(EXE_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(EXE_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(EXE_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(EXE_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(EXE_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(EXE_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(EXE_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(EXE_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(EXE_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(EXE_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(EXE_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(EXE_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(EXE_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(EXE_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(EXE_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(EXE_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(EXE_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(EXE_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(EXE_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(EXE_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(EXE_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(EXE_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(EXE_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(EXE_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(EXE_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(EXE_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(EXE_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(EXE_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(EXE_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(EXE_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(EXE_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(EXE_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(EXE_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(EXE_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(EXE_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(EXE_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(EXE_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(EXE_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(EXE_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(EXE_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(EXE_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(EXE_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(EXE_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(EXE_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(EXE_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(EXE_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(EXE_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(EXE_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(EXE_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(EXE_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(EXE_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(EXE_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(EXE_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(EXE_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(EXE_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(EXE_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(EXE_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(EXE_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(EXE_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(EXE_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(EXE_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(EXE_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(EXE_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(EXE_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(EXE_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(EXE_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(EXE_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(EXE_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(EXE_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(EXE_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(EXE_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(EXE_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(EXE_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(EXE_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(EXE_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(EXE_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(EXE_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(EXE_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(EXE_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(EXE_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(EXE_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(EXE_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(EXE_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(EXE_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(EXE_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(EXE_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(EXE_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(EXE_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(EXE_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(EXE_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(EXE_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(EXE_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(EXE_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(EXE_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(EXE_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(EXE_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(EXE_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(EXE_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(EXE_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(EXE_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(EXE_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(EXE_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(EXE_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(EXE_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(EXE_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(EXE_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(EXE_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(EXE_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(EXE_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(EXE_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(EXE_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(EXE_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(EXE_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(EXE_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(EXE_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(EXE_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(EXE_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(EXE_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(EXE_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(EXE_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(EXE_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(EXE_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(EXE_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(EXE_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(EXE_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(EXE_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(EXE_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(EXE_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(EXE_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(EXE_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(EXE_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(EXE_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(EXE_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(EXE_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(EXE_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(EXE_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(EXE_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(EXE_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(EXE_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(EXE_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(EXE_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(EXE_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(EXE_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(EXE_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(EXE_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(EXE_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(EXE_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(EXE_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(EXE_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(EXE_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(EXE_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(EXE_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(EXE_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(EXE_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(EXE_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(EXE_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(EXE_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(EXE_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(EXE_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(EXE_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(EXE_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(EXE_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(EXE_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(EXE_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(EXE_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(EXE_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(EXE_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(EXE_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(EXE_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(EXE_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(EXE_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(EXE_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(EXE_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(EXE_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(EXE_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(EXE_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(EXE_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(EXE_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(EXE_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(EXE_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(EXE_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(EXE_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(EXE_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(EXE_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(EXE_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(EXE_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(EXE_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(EXE_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(EXE_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(EXE_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(EXE_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(EXE_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(EXE_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(EXE_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(EXE_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(EXE_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(EXE_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(EXE_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(EXE_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(EXE_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(EXE_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(EXE_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(EXE_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(EXE_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(EXE_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(EXE_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(EXE_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(EXE_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(EXE_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(EXE_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(EXE_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(EXE_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(EXE_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(EXE_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(EXE_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(EXE_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(EXE_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(EXE_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(EXE_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(EXE_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(EXE_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(EXE_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(EXE_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(EXE_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(EXE_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(EXE_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(EXE_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(EXE_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(EXE_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(EXE_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(EXE_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(EXE_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(EXE_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(EXE_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(EXE_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(EXE_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(EXE_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(EXE_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(EXE_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(EXE_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(EXE_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(EXE_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(EXE_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(EXE_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(EXE_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(EXE_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(EXE_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(EXE_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(EXE_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(EXE_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(EXE_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(EXE_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(EXE_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(EXE_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(EXE_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(EXE_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(EXE_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(EXE_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(EXE_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(EXE_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(EXE_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(EXE_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(EXE_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(EXE_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(EXE_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(EXE_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(EXE_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(EXE_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(EXE_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(EXE_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(EXE_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(EXE_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(EXE_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(EXE_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(EXE_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(EXE_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(EXE_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(EXE_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(EXE_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(EXE_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(EXE_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(EXE_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(EXE_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(EXE_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(EXE_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(EXE_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(EXE_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(EXE_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(EXE_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(EXE_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(EXE_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(EXE_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(EXE_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(EXE_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(EXE_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(EXE_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(EXE_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(EXE_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(EXE_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(EXE_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(EXE_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(EXE_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(EXE_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(EXE_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(EXE_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(EXE_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(EXE_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(EXE_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(EXE_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(EXE_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(EXE_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(EXE_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(EXE_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(EXE_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(EXE_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(EXE_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(EXE_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(EXE_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(EXE_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(EXE_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(EXE_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(EXE_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(EXE_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(EXE_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(EXE_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(EXE_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(EXE_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(EXE_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(EXE_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(EXE_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(EXE_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(EXE_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(EXE_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(EXE_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(EXE_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(EXE_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(EXE_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(EXE_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(EXE_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(EXE_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(EXE_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(EXE_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(EXE_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(EXE_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(EXE_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(EXE_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(EXE_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(EXE_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(EXE_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(EXE_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(EXE_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(EXE_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(EXE_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(EXE_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(EXE_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(EXE_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(EXE_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(EXE_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(EXE_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(EXE_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(EXE_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(EXE_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(EXE_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(EXE_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(EXE_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(EXE_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(EXE_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(EXE_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(EXE_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(EXE_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(EXE_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(EXE_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(EXE_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(EXE_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(EXE_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(EXE_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(EXE_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(EXE_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(EXE_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(EXE_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(EXE_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(EXE_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(EXE_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(EXE_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(EXE_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(EXE_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(EXE_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(EXE_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(EXE_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(EXE_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(EXE_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(EXE_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(EXE_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(EXE_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(EXE_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(EXE_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(EXE_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(EXE_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(EXE_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(EXE_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(EXE_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(EXE_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(EXE_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(EXE_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(EXE_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(EXE_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(EXE_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(EXE_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(EXE_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(EXE_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(EXE_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(EXE_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(EXE_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(EXE_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(EXE_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(EXE_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(EXE_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(EXE_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(EXE_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(EXE_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(EXE_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(EXE_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(EXE_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(EXE_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(EXE_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(EXE_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(EXE_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(EXE_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(EXE_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(EXE_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(EXE_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(EXE_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(EXE_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(EXE_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(EXE_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(EXE_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(EXE_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(EXE_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(EXE_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(EXE_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(EXE_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(EXE_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(EXE_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(EXE_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(EXE_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(EXE_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(EXE_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(EXE_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(EXE_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(EXE_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(EXE_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(EXE_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(EXE_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(EXE_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(EXE_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(EXE_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(EXE_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(EXE_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(EXE_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(EXE_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(EXE_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(EXE_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(EXE_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(EXE_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(EXE_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(EXE_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(EXE_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(EXE_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(EXE_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(EXE_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(EXE_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(EXE_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(EXE_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(EXE_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(EXE_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(EXE_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(EXE_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(EXE_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(EXE_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(EXE_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(EXE_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(EXE_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(EXE_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(EXE_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(EXE_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(EXE_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(EXE_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(EXE_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(EXE_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(EXE_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(EXE_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(EXE_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(EXE_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(EXE_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(EXE_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(EXE_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(EXE_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(EXE_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(EXE_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(EXE_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(EXE_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(EXE_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(EXE_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(EXE_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(EXE_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(EXE_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(EXE_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(EXE_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(EXE_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(EXE_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(EXE_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(EXE_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(EXE_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(EXE_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(EXE_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(EXE_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(EXE_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(EXE_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(EXE_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(EXE_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(EXE_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(EXE_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(EXE_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(EXE_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(EXE_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(EXE_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(EXE_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(EXE_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(EXE_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(EXE_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(EXE_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(EXE_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(EXE_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(EXE_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(EXE_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(EXE_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(EXE_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(EXE_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(EXE_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(EXE_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(EXE_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(EXE_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(EXE_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(EXE_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(EXE_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(EXE_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(EXE_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(EXE_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(EXE_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(EXE_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(EXE_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(EXE_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(EXE_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(EXE_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(EXE_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(EXE_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(EXE_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(EXE_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(EXE_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(EXE_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(EXE_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(EXE_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(EXE_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(EXE_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(EXE_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(EXE_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(EXE_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(EXE_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(EXE_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(EXE_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(EXE_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(EXE_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(EXE_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(EXE_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(EXE_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(EXE_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(EXE_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(EXE_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(EXE_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(EXE_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(EXE_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(EXE_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(EXE_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(EXE_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(EXE_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(EXE_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(EXE_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(EXE_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(EXE_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(EXE_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(EXE_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(EXE_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(EXE_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(EXE_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(EXE_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(EXE_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(EXE_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(EXE_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(EXE_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(EXE_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(EXE_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(EXE_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(EXE_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(EXE_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(EXE_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(EXE_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(EXE_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(EXE_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(EXE_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(EXE_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(EXE_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(EXE_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(EXE_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(EXE_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(EXE_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(EXE_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(EXE_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(EXE_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(EXE_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(EXE_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(EXE_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(EXE_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(EXE_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(EXE_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(EXE_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(EXE_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(EXE_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(EXE_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(EXE_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(EXE_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(EXE_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(EXE_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(EXE_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(EXE_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(EXE_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(EXE_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(EXE_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(EXE_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(EXE_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(EXE_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(EXE_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(EXE_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(EXE_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(EXE_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(EXE_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(EXE_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(EXE_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(EXE_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(EXE_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(EXE_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(EXE_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(EXE_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(EXE_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(EXE_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(EXE_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(EXE_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(EXE_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(EXE_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(EXE_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(EXE_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(EXE_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(EXE_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(EXE_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(EXE_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(EXE_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(EXE_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(EXE_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(EXE_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(EXE_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(EXE_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(EXE_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(EXE_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(EXE_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(EXE_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(EXE_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(EXE_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(EXE_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(EXE_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(EXE_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(EXE_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(EXE_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(EXE_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(EXE_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(EXE_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(EXE_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(EXE_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(EXE_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(EXE_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(EXE_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(EXE_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(EXE_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(EXE_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(EXE_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(EXE_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(EXE_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(EXE_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(EXE_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(EXE_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(EXE_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(EXE_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(EXE_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(EXE_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(EXE_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(EXE_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(EXE_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(EXE_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(EXE_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(EXE_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(EXE_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(EXE_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(EXE_io_pipe_phv_out_next_config_id),
    .io_hit(EXE_io_hit),
    .io_match_value(EXE_io_match_value),
    .io_action_mod_en_0(EXE_io_action_mod_en_0),
    .io_action_mod_en_1(EXE_io_action_mod_en_1),
    .io_action_mod_addr(EXE_io_action_mod_addr),
    .io_action_mod_data_0(EXE_io_action_mod_data_0),
    .io_action_mod_data_1(EXE_io_action_mod_data_1)
  );
  assign io_pipe_phv_out_data_0 = EXE_io_pipe_phv_out_data_0; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_1 = EXE_io_pipe_phv_out_data_1; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_2 = EXE_io_pipe_phv_out_data_2; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_3 = EXE_io_pipe_phv_out_data_3; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_4 = EXE_io_pipe_phv_out_data_4; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_5 = EXE_io_pipe_phv_out_data_5; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_6 = EXE_io_pipe_phv_out_data_6; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_7 = EXE_io_pipe_phv_out_data_7; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_8 = EXE_io_pipe_phv_out_data_8; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_9 = EXE_io_pipe_phv_out_data_9; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_10 = EXE_io_pipe_phv_out_data_10; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_11 = EXE_io_pipe_phv_out_data_11; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_12 = EXE_io_pipe_phv_out_data_12; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_13 = EXE_io_pipe_phv_out_data_13; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_14 = EXE_io_pipe_phv_out_data_14; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_15 = EXE_io_pipe_phv_out_data_15; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_16 = EXE_io_pipe_phv_out_data_16; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_17 = EXE_io_pipe_phv_out_data_17; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_18 = EXE_io_pipe_phv_out_data_18; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_19 = EXE_io_pipe_phv_out_data_19; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_20 = EXE_io_pipe_phv_out_data_20; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_21 = EXE_io_pipe_phv_out_data_21; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_22 = EXE_io_pipe_phv_out_data_22; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_23 = EXE_io_pipe_phv_out_data_23; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_24 = EXE_io_pipe_phv_out_data_24; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_25 = EXE_io_pipe_phv_out_data_25; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_26 = EXE_io_pipe_phv_out_data_26; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_27 = EXE_io_pipe_phv_out_data_27; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_28 = EXE_io_pipe_phv_out_data_28; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_29 = EXE_io_pipe_phv_out_data_29; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_30 = EXE_io_pipe_phv_out_data_30; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_31 = EXE_io_pipe_phv_out_data_31; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_32 = EXE_io_pipe_phv_out_data_32; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_33 = EXE_io_pipe_phv_out_data_33; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_34 = EXE_io_pipe_phv_out_data_34; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_35 = EXE_io_pipe_phv_out_data_35; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_36 = EXE_io_pipe_phv_out_data_36; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_37 = EXE_io_pipe_phv_out_data_37; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_38 = EXE_io_pipe_phv_out_data_38; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_39 = EXE_io_pipe_phv_out_data_39; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_40 = EXE_io_pipe_phv_out_data_40; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_41 = EXE_io_pipe_phv_out_data_41; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_42 = EXE_io_pipe_phv_out_data_42; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_43 = EXE_io_pipe_phv_out_data_43; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_44 = EXE_io_pipe_phv_out_data_44; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_45 = EXE_io_pipe_phv_out_data_45; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_46 = EXE_io_pipe_phv_out_data_46; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_47 = EXE_io_pipe_phv_out_data_47; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_48 = EXE_io_pipe_phv_out_data_48; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_49 = EXE_io_pipe_phv_out_data_49; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_50 = EXE_io_pipe_phv_out_data_50; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_51 = EXE_io_pipe_phv_out_data_51; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_52 = EXE_io_pipe_phv_out_data_52; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_53 = EXE_io_pipe_phv_out_data_53; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_54 = EXE_io_pipe_phv_out_data_54; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_55 = EXE_io_pipe_phv_out_data_55; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_56 = EXE_io_pipe_phv_out_data_56; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_57 = EXE_io_pipe_phv_out_data_57; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_58 = EXE_io_pipe_phv_out_data_58; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_59 = EXE_io_pipe_phv_out_data_59; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_60 = EXE_io_pipe_phv_out_data_60; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_61 = EXE_io_pipe_phv_out_data_61; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_62 = EXE_io_pipe_phv_out_data_62; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_63 = EXE_io_pipe_phv_out_data_63; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_64 = EXE_io_pipe_phv_out_data_64; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_65 = EXE_io_pipe_phv_out_data_65; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_66 = EXE_io_pipe_phv_out_data_66; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_67 = EXE_io_pipe_phv_out_data_67; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_68 = EXE_io_pipe_phv_out_data_68; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_69 = EXE_io_pipe_phv_out_data_69; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_70 = EXE_io_pipe_phv_out_data_70; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_71 = EXE_io_pipe_phv_out_data_71; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_72 = EXE_io_pipe_phv_out_data_72; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_73 = EXE_io_pipe_phv_out_data_73; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_74 = EXE_io_pipe_phv_out_data_74; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_75 = EXE_io_pipe_phv_out_data_75; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_76 = EXE_io_pipe_phv_out_data_76; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_77 = EXE_io_pipe_phv_out_data_77; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_78 = EXE_io_pipe_phv_out_data_78; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_79 = EXE_io_pipe_phv_out_data_79; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_80 = EXE_io_pipe_phv_out_data_80; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_81 = EXE_io_pipe_phv_out_data_81; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_82 = EXE_io_pipe_phv_out_data_82; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_83 = EXE_io_pipe_phv_out_data_83; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_84 = EXE_io_pipe_phv_out_data_84; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_85 = EXE_io_pipe_phv_out_data_85; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_86 = EXE_io_pipe_phv_out_data_86; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_87 = EXE_io_pipe_phv_out_data_87; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_88 = EXE_io_pipe_phv_out_data_88; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_89 = EXE_io_pipe_phv_out_data_89; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_90 = EXE_io_pipe_phv_out_data_90; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_91 = EXE_io_pipe_phv_out_data_91; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_92 = EXE_io_pipe_phv_out_data_92; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_93 = EXE_io_pipe_phv_out_data_93; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_94 = EXE_io_pipe_phv_out_data_94; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_95 = EXE_io_pipe_phv_out_data_95; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_96 = EXE_io_pipe_phv_out_data_96; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_97 = EXE_io_pipe_phv_out_data_97; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_98 = EXE_io_pipe_phv_out_data_98; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_99 = EXE_io_pipe_phv_out_data_99; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_100 = EXE_io_pipe_phv_out_data_100; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_101 = EXE_io_pipe_phv_out_data_101; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_102 = EXE_io_pipe_phv_out_data_102; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_103 = EXE_io_pipe_phv_out_data_103; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_104 = EXE_io_pipe_phv_out_data_104; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_105 = EXE_io_pipe_phv_out_data_105; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_106 = EXE_io_pipe_phv_out_data_106; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_107 = EXE_io_pipe_phv_out_data_107; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_108 = EXE_io_pipe_phv_out_data_108; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_109 = EXE_io_pipe_phv_out_data_109; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_110 = EXE_io_pipe_phv_out_data_110; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_111 = EXE_io_pipe_phv_out_data_111; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_112 = EXE_io_pipe_phv_out_data_112; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_113 = EXE_io_pipe_phv_out_data_113; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_114 = EXE_io_pipe_phv_out_data_114; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_115 = EXE_io_pipe_phv_out_data_115; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_116 = EXE_io_pipe_phv_out_data_116; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_117 = EXE_io_pipe_phv_out_data_117; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_118 = EXE_io_pipe_phv_out_data_118; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_119 = EXE_io_pipe_phv_out_data_119; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_120 = EXE_io_pipe_phv_out_data_120; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_121 = EXE_io_pipe_phv_out_data_121; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_122 = EXE_io_pipe_phv_out_data_122; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_123 = EXE_io_pipe_phv_out_data_123; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_124 = EXE_io_pipe_phv_out_data_124; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_125 = EXE_io_pipe_phv_out_data_125; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_126 = EXE_io_pipe_phv_out_data_126; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_127 = EXE_io_pipe_phv_out_data_127; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_128 = EXE_io_pipe_phv_out_data_128; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_129 = EXE_io_pipe_phv_out_data_129; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_130 = EXE_io_pipe_phv_out_data_130; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_131 = EXE_io_pipe_phv_out_data_131; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_132 = EXE_io_pipe_phv_out_data_132; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_133 = EXE_io_pipe_phv_out_data_133; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_134 = EXE_io_pipe_phv_out_data_134; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_135 = EXE_io_pipe_phv_out_data_135; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_136 = EXE_io_pipe_phv_out_data_136; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_137 = EXE_io_pipe_phv_out_data_137; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_138 = EXE_io_pipe_phv_out_data_138; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_139 = EXE_io_pipe_phv_out_data_139; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_140 = EXE_io_pipe_phv_out_data_140; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_141 = EXE_io_pipe_phv_out_data_141; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_142 = EXE_io_pipe_phv_out_data_142; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_143 = EXE_io_pipe_phv_out_data_143; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_144 = EXE_io_pipe_phv_out_data_144; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_145 = EXE_io_pipe_phv_out_data_145; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_146 = EXE_io_pipe_phv_out_data_146; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_147 = EXE_io_pipe_phv_out_data_147; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_148 = EXE_io_pipe_phv_out_data_148; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_149 = EXE_io_pipe_phv_out_data_149; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_150 = EXE_io_pipe_phv_out_data_150; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_151 = EXE_io_pipe_phv_out_data_151; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_152 = EXE_io_pipe_phv_out_data_152; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_153 = EXE_io_pipe_phv_out_data_153; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_154 = EXE_io_pipe_phv_out_data_154; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_155 = EXE_io_pipe_phv_out_data_155; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_156 = EXE_io_pipe_phv_out_data_156; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_157 = EXE_io_pipe_phv_out_data_157; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_158 = EXE_io_pipe_phv_out_data_158; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_159 = EXE_io_pipe_phv_out_data_159; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_160 = EXE_io_pipe_phv_out_data_160; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_161 = EXE_io_pipe_phv_out_data_161; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_162 = EXE_io_pipe_phv_out_data_162; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_163 = EXE_io_pipe_phv_out_data_163; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_164 = EXE_io_pipe_phv_out_data_164; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_165 = EXE_io_pipe_phv_out_data_165; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_166 = EXE_io_pipe_phv_out_data_166; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_167 = EXE_io_pipe_phv_out_data_167; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_168 = EXE_io_pipe_phv_out_data_168; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_169 = EXE_io_pipe_phv_out_data_169; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_170 = EXE_io_pipe_phv_out_data_170; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_171 = EXE_io_pipe_phv_out_data_171; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_172 = EXE_io_pipe_phv_out_data_172; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_173 = EXE_io_pipe_phv_out_data_173; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_174 = EXE_io_pipe_phv_out_data_174; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_175 = EXE_io_pipe_phv_out_data_175; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_176 = EXE_io_pipe_phv_out_data_176; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_177 = EXE_io_pipe_phv_out_data_177; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_178 = EXE_io_pipe_phv_out_data_178; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_179 = EXE_io_pipe_phv_out_data_179; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_180 = EXE_io_pipe_phv_out_data_180; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_181 = EXE_io_pipe_phv_out_data_181; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_182 = EXE_io_pipe_phv_out_data_182; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_183 = EXE_io_pipe_phv_out_data_183; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_184 = EXE_io_pipe_phv_out_data_184; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_185 = EXE_io_pipe_phv_out_data_185; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_186 = EXE_io_pipe_phv_out_data_186; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_187 = EXE_io_pipe_phv_out_data_187; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_188 = EXE_io_pipe_phv_out_data_188; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_189 = EXE_io_pipe_phv_out_data_189; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_190 = EXE_io_pipe_phv_out_data_190; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_191 = EXE_io_pipe_phv_out_data_191; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_192 = EXE_io_pipe_phv_out_data_192; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_193 = EXE_io_pipe_phv_out_data_193; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_194 = EXE_io_pipe_phv_out_data_194; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_195 = EXE_io_pipe_phv_out_data_195; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_196 = EXE_io_pipe_phv_out_data_196; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_197 = EXE_io_pipe_phv_out_data_197; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_198 = EXE_io_pipe_phv_out_data_198; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_199 = EXE_io_pipe_phv_out_data_199; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_200 = EXE_io_pipe_phv_out_data_200; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_201 = EXE_io_pipe_phv_out_data_201; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_202 = EXE_io_pipe_phv_out_data_202; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_203 = EXE_io_pipe_phv_out_data_203; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_204 = EXE_io_pipe_phv_out_data_204; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_205 = EXE_io_pipe_phv_out_data_205; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_206 = EXE_io_pipe_phv_out_data_206; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_207 = EXE_io_pipe_phv_out_data_207; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_208 = EXE_io_pipe_phv_out_data_208; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_209 = EXE_io_pipe_phv_out_data_209; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_210 = EXE_io_pipe_phv_out_data_210; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_211 = EXE_io_pipe_phv_out_data_211; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_212 = EXE_io_pipe_phv_out_data_212; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_213 = EXE_io_pipe_phv_out_data_213; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_214 = EXE_io_pipe_phv_out_data_214; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_215 = EXE_io_pipe_phv_out_data_215; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_216 = EXE_io_pipe_phv_out_data_216; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_217 = EXE_io_pipe_phv_out_data_217; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_218 = EXE_io_pipe_phv_out_data_218; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_219 = EXE_io_pipe_phv_out_data_219; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_220 = EXE_io_pipe_phv_out_data_220; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_221 = EXE_io_pipe_phv_out_data_221; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_222 = EXE_io_pipe_phv_out_data_222; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_223 = EXE_io_pipe_phv_out_data_223; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_224 = EXE_io_pipe_phv_out_data_224; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_225 = EXE_io_pipe_phv_out_data_225; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_226 = EXE_io_pipe_phv_out_data_226; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_227 = EXE_io_pipe_phv_out_data_227; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_228 = EXE_io_pipe_phv_out_data_228; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_229 = EXE_io_pipe_phv_out_data_229; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_230 = EXE_io_pipe_phv_out_data_230; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_231 = EXE_io_pipe_phv_out_data_231; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_232 = EXE_io_pipe_phv_out_data_232; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_233 = EXE_io_pipe_phv_out_data_233; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_234 = EXE_io_pipe_phv_out_data_234; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_235 = EXE_io_pipe_phv_out_data_235; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_236 = EXE_io_pipe_phv_out_data_236; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_237 = EXE_io_pipe_phv_out_data_237; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_238 = EXE_io_pipe_phv_out_data_238; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_239 = EXE_io_pipe_phv_out_data_239; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_240 = EXE_io_pipe_phv_out_data_240; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_241 = EXE_io_pipe_phv_out_data_241; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_242 = EXE_io_pipe_phv_out_data_242; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_243 = EXE_io_pipe_phv_out_data_243; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_244 = EXE_io_pipe_phv_out_data_244; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_245 = EXE_io_pipe_phv_out_data_245; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_246 = EXE_io_pipe_phv_out_data_246; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_247 = EXE_io_pipe_phv_out_data_247; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_248 = EXE_io_pipe_phv_out_data_248; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_249 = EXE_io_pipe_phv_out_data_249; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_250 = EXE_io_pipe_phv_out_data_250; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_251 = EXE_io_pipe_phv_out_data_251; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_252 = EXE_io_pipe_phv_out_data_252; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_253 = EXE_io_pipe_phv_out_data_253; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_254 = EXE_io_pipe_phv_out_data_254; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_255 = EXE_io_pipe_phv_out_data_255; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_256 = EXE_io_pipe_phv_out_data_256; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_257 = EXE_io_pipe_phv_out_data_257; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_258 = EXE_io_pipe_phv_out_data_258; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_259 = EXE_io_pipe_phv_out_data_259; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_260 = EXE_io_pipe_phv_out_data_260; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_261 = EXE_io_pipe_phv_out_data_261; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_262 = EXE_io_pipe_phv_out_data_262; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_263 = EXE_io_pipe_phv_out_data_263; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_264 = EXE_io_pipe_phv_out_data_264; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_265 = EXE_io_pipe_phv_out_data_265; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_266 = EXE_io_pipe_phv_out_data_266; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_267 = EXE_io_pipe_phv_out_data_267; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_268 = EXE_io_pipe_phv_out_data_268; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_269 = EXE_io_pipe_phv_out_data_269; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_270 = EXE_io_pipe_phv_out_data_270; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_271 = EXE_io_pipe_phv_out_data_271; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_272 = EXE_io_pipe_phv_out_data_272; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_273 = EXE_io_pipe_phv_out_data_273; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_274 = EXE_io_pipe_phv_out_data_274; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_275 = EXE_io_pipe_phv_out_data_275; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_276 = EXE_io_pipe_phv_out_data_276; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_277 = EXE_io_pipe_phv_out_data_277; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_278 = EXE_io_pipe_phv_out_data_278; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_279 = EXE_io_pipe_phv_out_data_279; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_280 = EXE_io_pipe_phv_out_data_280; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_281 = EXE_io_pipe_phv_out_data_281; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_282 = EXE_io_pipe_phv_out_data_282; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_283 = EXE_io_pipe_phv_out_data_283; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_284 = EXE_io_pipe_phv_out_data_284; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_285 = EXE_io_pipe_phv_out_data_285; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_286 = EXE_io_pipe_phv_out_data_286; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_287 = EXE_io_pipe_phv_out_data_287; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_288 = EXE_io_pipe_phv_out_data_288; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_289 = EXE_io_pipe_phv_out_data_289; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_290 = EXE_io_pipe_phv_out_data_290; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_291 = EXE_io_pipe_phv_out_data_291; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_292 = EXE_io_pipe_phv_out_data_292; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_293 = EXE_io_pipe_phv_out_data_293; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_294 = EXE_io_pipe_phv_out_data_294; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_295 = EXE_io_pipe_phv_out_data_295; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_296 = EXE_io_pipe_phv_out_data_296; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_297 = EXE_io_pipe_phv_out_data_297; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_298 = EXE_io_pipe_phv_out_data_298; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_299 = EXE_io_pipe_phv_out_data_299; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_300 = EXE_io_pipe_phv_out_data_300; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_301 = EXE_io_pipe_phv_out_data_301; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_302 = EXE_io_pipe_phv_out_data_302; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_303 = EXE_io_pipe_phv_out_data_303; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_304 = EXE_io_pipe_phv_out_data_304; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_305 = EXE_io_pipe_phv_out_data_305; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_306 = EXE_io_pipe_phv_out_data_306; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_307 = EXE_io_pipe_phv_out_data_307; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_308 = EXE_io_pipe_phv_out_data_308; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_309 = EXE_io_pipe_phv_out_data_309; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_310 = EXE_io_pipe_phv_out_data_310; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_311 = EXE_io_pipe_phv_out_data_311; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_312 = EXE_io_pipe_phv_out_data_312; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_313 = EXE_io_pipe_phv_out_data_313; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_314 = EXE_io_pipe_phv_out_data_314; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_315 = EXE_io_pipe_phv_out_data_315; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_316 = EXE_io_pipe_phv_out_data_316; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_317 = EXE_io_pipe_phv_out_data_317; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_318 = EXE_io_pipe_phv_out_data_318; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_319 = EXE_io_pipe_phv_out_data_319; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_320 = EXE_io_pipe_phv_out_data_320; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_321 = EXE_io_pipe_phv_out_data_321; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_322 = EXE_io_pipe_phv_out_data_322; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_323 = EXE_io_pipe_phv_out_data_323; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_324 = EXE_io_pipe_phv_out_data_324; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_325 = EXE_io_pipe_phv_out_data_325; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_326 = EXE_io_pipe_phv_out_data_326; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_327 = EXE_io_pipe_phv_out_data_327; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_328 = EXE_io_pipe_phv_out_data_328; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_329 = EXE_io_pipe_phv_out_data_329; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_330 = EXE_io_pipe_phv_out_data_330; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_331 = EXE_io_pipe_phv_out_data_331; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_332 = EXE_io_pipe_phv_out_data_332; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_333 = EXE_io_pipe_phv_out_data_333; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_334 = EXE_io_pipe_phv_out_data_334; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_335 = EXE_io_pipe_phv_out_data_335; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_336 = EXE_io_pipe_phv_out_data_336; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_337 = EXE_io_pipe_phv_out_data_337; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_338 = EXE_io_pipe_phv_out_data_338; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_339 = EXE_io_pipe_phv_out_data_339; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_340 = EXE_io_pipe_phv_out_data_340; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_341 = EXE_io_pipe_phv_out_data_341; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_342 = EXE_io_pipe_phv_out_data_342; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_343 = EXE_io_pipe_phv_out_data_343; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_344 = EXE_io_pipe_phv_out_data_344; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_345 = EXE_io_pipe_phv_out_data_345; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_346 = EXE_io_pipe_phv_out_data_346; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_347 = EXE_io_pipe_phv_out_data_347; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_348 = EXE_io_pipe_phv_out_data_348; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_349 = EXE_io_pipe_phv_out_data_349; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_350 = EXE_io_pipe_phv_out_data_350; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_351 = EXE_io_pipe_phv_out_data_351; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_352 = EXE_io_pipe_phv_out_data_352; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_353 = EXE_io_pipe_phv_out_data_353; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_354 = EXE_io_pipe_phv_out_data_354; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_355 = EXE_io_pipe_phv_out_data_355; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_356 = EXE_io_pipe_phv_out_data_356; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_357 = EXE_io_pipe_phv_out_data_357; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_358 = EXE_io_pipe_phv_out_data_358; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_359 = EXE_io_pipe_phv_out_data_359; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_360 = EXE_io_pipe_phv_out_data_360; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_361 = EXE_io_pipe_phv_out_data_361; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_362 = EXE_io_pipe_phv_out_data_362; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_363 = EXE_io_pipe_phv_out_data_363; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_364 = EXE_io_pipe_phv_out_data_364; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_365 = EXE_io_pipe_phv_out_data_365; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_366 = EXE_io_pipe_phv_out_data_366; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_367 = EXE_io_pipe_phv_out_data_367; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_368 = EXE_io_pipe_phv_out_data_368; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_369 = EXE_io_pipe_phv_out_data_369; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_370 = EXE_io_pipe_phv_out_data_370; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_371 = EXE_io_pipe_phv_out_data_371; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_372 = EXE_io_pipe_phv_out_data_372; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_373 = EXE_io_pipe_phv_out_data_373; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_374 = EXE_io_pipe_phv_out_data_374; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_375 = EXE_io_pipe_phv_out_data_375; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_376 = EXE_io_pipe_phv_out_data_376; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_377 = EXE_io_pipe_phv_out_data_377; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_378 = EXE_io_pipe_phv_out_data_378; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_379 = EXE_io_pipe_phv_out_data_379; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_380 = EXE_io_pipe_phv_out_data_380; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_381 = EXE_io_pipe_phv_out_data_381; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_382 = EXE_io_pipe_phv_out_data_382; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_383 = EXE_io_pipe_phv_out_data_383; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_384 = EXE_io_pipe_phv_out_data_384; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_385 = EXE_io_pipe_phv_out_data_385; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_386 = EXE_io_pipe_phv_out_data_386; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_387 = EXE_io_pipe_phv_out_data_387; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_388 = EXE_io_pipe_phv_out_data_388; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_389 = EXE_io_pipe_phv_out_data_389; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_390 = EXE_io_pipe_phv_out_data_390; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_391 = EXE_io_pipe_phv_out_data_391; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_392 = EXE_io_pipe_phv_out_data_392; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_393 = EXE_io_pipe_phv_out_data_393; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_394 = EXE_io_pipe_phv_out_data_394; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_395 = EXE_io_pipe_phv_out_data_395; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_396 = EXE_io_pipe_phv_out_data_396; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_397 = EXE_io_pipe_phv_out_data_397; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_398 = EXE_io_pipe_phv_out_data_398; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_399 = EXE_io_pipe_phv_out_data_399; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_400 = EXE_io_pipe_phv_out_data_400; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_401 = EXE_io_pipe_phv_out_data_401; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_402 = EXE_io_pipe_phv_out_data_402; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_403 = EXE_io_pipe_phv_out_data_403; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_404 = EXE_io_pipe_phv_out_data_404; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_405 = EXE_io_pipe_phv_out_data_405; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_406 = EXE_io_pipe_phv_out_data_406; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_407 = EXE_io_pipe_phv_out_data_407; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_408 = EXE_io_pipe_phv_out_data_408; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_409 = EXE_io_pipe_phv_out_data_409; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_410 = EXE_io_pipe_phv_out_data_410; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_411 = EXE_io_pipe_phv_out_data_411; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_412 = EXE_io_pipe_phv_out_data_412; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_413 = EXE_io_pipe_phv_out_data_413; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_414 = EXE_io_pipe_phv_out_data_414; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_415 = EXE_io_pipe_phv_out_data_415; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_416 = EXE_io_pipe_phv_out_data_416; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_417 = EXE_io_pipe_phv_out_data_417; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_418 = EXE_io_pipe_phv_out_data_418; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_419 = EXE_io_pipe_phv_out_data_419; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_420 = EXE_io_pipe_phv_out_data_420; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_421 = EXE_io_pipe_phv_out_data_421; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_422 = EXE_io_pipe_phv_out_data_422; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_423 = EXE_io_pipe_phv_out_data_423; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_424 = EXE_io_pipe_phv_out_data_424; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_425 = EXE_io_pipe_phv_out_data_425; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_426 = EXE_io_pipe_phv_out_data_426; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_427 = EXE_io_pipe_phv_out_data_427; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_428 = EXE_io_pipe_phv_out_data_428; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_429 = EXE_io_pipe_phv_out_data_429; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_430 = EXE_io_pipe_phv_out_data_430; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_431 = EXE_io_pipe_phv_out_data_431; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_432 = EXE_io_pipe_phv_out_data_432; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_433 = EXE_io_pipe_phv_out_data_433; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_434 = EXE_io_pipe_phv_out_data_434; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_435 = EXE_io_pipe_phv_out_data_435; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_436 = EXE_io_pipe_phv_out_data_436; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_437 = EXE_io_pipe_phv_out_data_437; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_438 = EXE_io_pipe_phv_out_data_438; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_439 = EXE_io_pipe_phv_out_data_439; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_440 = EXE_io_pipe_phv_out_data_440; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_441 = EXE_io_pipe_phv_out_data_441; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_442 = EXE_io_pipe_phv_out_data_442; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_443 = EXE_io_pipe_phv_out_data_443; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_444 = EXE_io_pipe_phv_out_data_444; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_445 = EXE_io_pipe_phv_out_data_445; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_446 = EXE_io_pipe_phv_out_data_446; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_447 = EXE_io_pipe_phv_out_data_447; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_448 = EXE_io_pipe_phv_out_data_448; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_449 = EXE_io_pipe_phv_out_data_449; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_450 = EXE_io_pipe_phv_out_data_450; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_451 = EXE_io_pipe_phv_out_data_451; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_452 = EXE_io_pipe_phv_out_data_452; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_453 = EXE_io_pipe_phv_out_data_453; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_454 = EXE_io_pipe_phv_out_data_454; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_455 = EXE_io_pipe_phv_out_data_455; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_456 = EXE_io_pipe_phv_out_data_456; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_457 = EXE_io_pipe_phv_out_data_457; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_458 = EXE_io_pipe_phv_out_data_458; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_459 = EXE_io_pipe_phv_out_data_459; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_460 = EXE_io_pipe_phv_out_data_460; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_461 = EXE_io_pipe_phv_out_data_461; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_462 = EXE_io_pipe_phv_out_data_462; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_463 = EXE_io_pipe_phv_out_data_463; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_464 = EXE_io_pipe_phv_out_data_464; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_465 = EXE_io_pipe_phv_out_data_465; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_466 = EXE_io_pipe_phv_out_data_466; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_467 = EXE_io_pipe_phv_out_data_467; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_468 = EXE_io_pipe_phv_out_data_468; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_469 = EXE_io_pipe_phv_out_data_469; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_470 = EXE_io_pipe_phv_out_data_470; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_471 = EXE_io_pipe_phv_out_data_471; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_472 = EXE_io_pipe_phv_out_data_472; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_473 = EXE_io_pipe_phv_out_data_473; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_474 = EXE_io_pipe_phv_out_data_474; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_475 = EXE_io_pipe_phv_out_data_475; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_476 = EXE_io_pipe_phv_out_data_476; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_477 = EXE_io_pipe_phv_out_data_477; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_478 = EXE_io_pipe_phv_out_data_478; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_479 = EXE_io_pipe_phv_out_data_479; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_480 = EXE_io_pipe_phv_out_data_480; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_481 = EXE_io_pipe_phv_out_data_481; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_482 = EXE_io_pipe_phv_out_data_482; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_483 = EXE_io_pipe_phv_out_data_483; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_484 = EXE_io_pipe_phv_out_data_484; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_485 = EXE_io_pipe_phv_out_data_485; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_486 = EXE_io_pipe_phv_out_data_486; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_487 = EXE_io_pipe_phv_out_data_487; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_488 = EXE_io_pipe_phv_out_data_488; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_489 = EXE_io_pipe_phv_out_data_489; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_490 = EXE_io_pipe_phv_out_data_490; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_491 = EXE_io_pipe_phv_out_data_491; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_492 = EXE_io_pipe_phv_out_data_492; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_493 = EXE_io_pipe_phv_out_data_493; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_494 = EXE_io_pipe_phv_out_data_494; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_495 = EXE_io_pipe_phv_out_data_495; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_496 = EXE_io_pipe_phv_out_data_496; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_497 = EXE_io_pipe_phv_out_data_497; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_498 = EXE_io_pipe_phv_out_data_498; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_499 = EXE_io_pipe_phv_out_data_499; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_500 = EXE_io_pipe_phv_out_data_500; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_501 = EXE_io_pipe_phv_out_data_501; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_502 = EXE_io_pipe_phv_out_data_502; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_503 = EXE_io_pipe_phv_out_data_503; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_504 = EXE_io_pipe_phv_out_data_504; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_505 = EXE_io_pipe_phv_out_data_505; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_506 = EXE_io_pipe_phv_out_data_506; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_507 = EXE_io_pipe_phv_out_data_507; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_508 = EXE_io_pipe_phv_out_data_508; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_509 = EXE_io_pipe_phv_out_data_509; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_510 = EXE_io_pipe_phv_out_data_510; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_511 = EXE_io_pipe_phv_out_data_511; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_0 = EXE_io_pipe_phv_out_header_0; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_1 = EXE_io_pipe_phv_out_header_1; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_2 = EXE_io_pipe_phv_out_header_2; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_3 = EXE_io_pipe_phv_out_header_3; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_4 = EXE_io_pipe_phv_out_header_4; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_5 = EXE_io_pipe_phv_out_header_5; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_6 = EXE_io_pipe_phv_out_header_6; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_7 = EXE_io_pipe_phv_out_header_7; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_8 = EXE_io_pipe_phv_out_header_8; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_9 = EXE_io_pipe_phv_out_header_9; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_10 = EXE_io_pipe_phv_out_header_10; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_11 = EXE_io_pipe_phv_out_header_11; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_12 = EXE_io_pipe_phv_out_header_12; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_13 = EXE_io_pipe_phv_out_header_13; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_14 = EXE_io_pipe_phv_out_header_14; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_15 = EXE_io_pipe_phv_out_header_15; // @[processor.scala 29:24]
  assign io_pipe_phv_out_parse_current_state = EXE_io_pipe_phv_out_parse_current_state; // @[processor.scala 29:24]
  assign io_pipe_phv_out_parse_current_offset = EXE_io_pipe_phv_out_parse_current_offset; // @[processor.scala 29:24]
  assign io_pipe_phv_out_parse_transition_field = EXE_io_pipe_phv_out_parse_transition_field; // @[processor.scala 29:24]
  assign io_pipe_phv_out_next_processor_id = EXE_io_pipe_phv_out_next_processor_id; // @[processor.scala 29:24]
  assign io_pipe_phv_out_next_config_id = EXE_io_pipe_phv_out_next_config_id; // @[processor.scala 29:24]
  assign io_mem_cluster_0_en = MAT_io_mem_cluster_0_en; // @[processor.scala 22:24]
  assign io_mem_cluster_0_addr = MAT_io_mem_cluster_0_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_1_en = MAT_io_mem_cluster_1_en; // @[processor.scala 22:24]
  assign io_mem_cluster_1_addr = MAT_io_mem_cluster_1_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_2_en = MAT_io_mem_cluster_2_en; // @[processor.scala 22:24]
  assign io_mem_cluster_2_addr = MAT_io_mem_cluster_2_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_3_en = MAT_io_mem_cluster_3_en; // @[processor.scala 22:24]
  assign io_mem_cluster_3_addr = MAT_io_mem_cluster_3_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_4_en = MAT_io_mem_cluster_4_en; // @[processor.scala 22:24]
  assign io_mem_cluster_4_addr = MAT_io_mem_cluster_4_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_5_en = MAT_io_mem_cluster_5_en; // @[processor.scala 22:24]
  assign io_mem_cluster_5_addr = MAT_io_mem_cluster_5_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_6_en = MAT_io_mem_cluster_6_en; // @[processor.scala 22:24]
  assign io_mem_cluster_6_addr = MAT_io_mem_cluster_6_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_7_en = MAT_io_mem_cluster_7_en; // @[processor.scala 22:24]
  assign io_mem_cluster_7_addr = MAT_io_mem_cluster_7_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_8_en = MAT_io_mem_cluster_8_en; // @[processor.scala 22:24]
  assign io_mem_cluster_8_addr = MAT_io_mem_cluster_8_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_9_en = MAT_io_mem_cluster_9_en; // @[processor.scala 22:24]
  assign io_mem_cluster_9_addr = MAT_io_mem_cluster_9_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_10_en = MAT_io_mem_cluster_10_en; // @[processor.scala 22:24]
  assign io_mem_cluster_10_addr = MAT_io_mem_cluster_10_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_11_en = MAT_io_mem_cluster_11_en; // @[processor.scala 22:24]
  assign io_mem_cluster_11_addr = MAT_io_mem_cluster_11_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_12_en = MAT_io_mem_cluster_12_en; // @[processor.scala 22:24]
  assign io_mem_cluster_12_addr = MAT_io_mem_cluster_12_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_13_en = MAT_io_mem_cluster_13_en; // @[processor.scala 22:24]
  assign io_mem_cluster_13_addr = MAT_io_mem_cluster_13_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_14_en = MAT_io_mem_cluster_14_en; // @[processor.scala 22:24]
  assign io_mem_cluster_14_addr = MAT_io_mem_cluster_14_addr; // @[processor.scala 22:24]
  assign io_mem_cluster_15_en = MAT_io_mem_cluster_15_en; // @[processor.scala 22:24]
  assign io_mem_cluster_15_addr = MAT_io_mem_cluster_15_addr; // @[processor.scala 22:24]
  assign PAR_clock = clock;
  assign PAR_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_160 = io_pipe_phv_in_data_160; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_161 = io_pipe_phv_in_data_161; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_162 = io_pipe_phv_in_data_162; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_163 = io_pipe_phv_in_data_163; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_164 = io_pipe_phv_in_data_164; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_165 = io_pipe_phv_in_data_165; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_166 = io_pipe_phv_in_data_166; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_167 = io_pipe_phv_in_data_167; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_168 = io_pipe_phv_in_data_168; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_169 = io_pipe_phv_in_data_169; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_170 = io_pipe_phv_in_data_170; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_171 = io_pipe_phv_in_data_171; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_172 = io_pipe_phv_in_data_172; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_173 = io_pipe_phv_in_data_173; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_174 = io_pipe_phv_in_data_174; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_175 = io_pipe_phv_in_data_175; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_176 = io_pipe_phv_in_data_176; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_177 = io_pipe_phv_in_data_177; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_178 = io_pipe_phv_in_data_178; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_179 = io_pipe_phv_in_data_179; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_180 = io_pipe_phv_in_data_180; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_181 = io_pipe_phv_in_data_181; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_182 = io_pipe_phv_in_data_182; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_183 = io_pipe_phv_in_data_183; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_184 = io_pipe_phv_in_data_184; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_185 = io_pipe_phv_in_data_185; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_186 = io_pipe_phv_in_data_186; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_187 = io_pipe_phv_in_data_187; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_188 = io_pipe_phv_in_data_188; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_189 = io_pipe_phv_in_data_189; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_190 = io_pipe_phv_in_data_190; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_191 = io_pipe_phv_in_data_191; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_192 = io_pipe_phv_in_data_192; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_193 = io_pipe_phv_in_data_193; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_194 = io_pipe_phv_in_data_194; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_195 = io_pipe_phv_in_data_195; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_196 = io_pipe_phv_in_data_196; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_197 = io_pipe_phv_in_data_197; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_198 = io_pipe_phv_in_data_198; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_199 = io_pipe_phv_in_data_199; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_200 = io_pipe_phv_in_data_200; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_201 = io_pipe_phv_in_data_201; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_202 = io_pipe_phv_in_data_202; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_203 = io_pipe_phv_in_data_203; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_204 = io_pipe_phv_in_data_204; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_205 = io_pipe_phv_in_data_205; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_206 = io_pipe_phv_in_data_206; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_207 = io_pipe_phv_in_data_207; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_208 = io_pipe_phv_in_data_208; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_209 = io_pipe_phv_in_data_209; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_210 = io_pipe_phv_in_data_210; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_211 = io_pipe_phv_in_data_211; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_212 = io_pipe_phv_in_data_212; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_213 = io_pipe_phv_in_data_213; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_214 = io_pipe_phv_in_data_214; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_215 = io_pipe_phv_in_data_215; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_216 = io_pipe_phv_in_data_216; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_217 = io_pipe_phv_in_data_217; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_218 = io_pipe_phv_in_data_218; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_219 = io_pipe_phv_in_data_219; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_220 = io_pipe_phv_in_data_220; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_221 = io_pipe_phv_in_data_221; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_222 = io_pipe_phv_in_data_222; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_223 = io_pipe_phv_in_data_223; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_224 = io_pipe_phv_in_data_224; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_225 = io_pipe_phv_in_data_225; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_226 = io_pipe_phv_in_data_226; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_227 = io_pipe_phv_in_data_227; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_228 = io_pipe_phv_in_data_228; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_229 = io_pipe_phv_in_data_229; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_230 = io_pipe_phv_in_data_230; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_231 = io_pipe_phv_in_data_231; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_232 = io_pipe_phv_in_data_232; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_233 = io_pipe_phv_in_data_233; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_234 = io_pipe_phv_in_data_234; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_235 = io_pipe_phv_in_data_235; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_236 = io_pipe_phv_in_data_236; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_237 = io_pipe_phv_in_data_237; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_238 = io_pipe_phv_in_data_238; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_239 = io_pipe_phv_in_data_239; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_240 = io_pipe_phv_in_data_240; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_241 = io_pipe_phv_in_data_241; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_242 = io_pipe_phv_in_data_242; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_243 = io_pipe_phv_in_data_243; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_244 = io_pipe_phv_in_data_244; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_245 = io_pipe_phv_in_data_245; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_246 = io_pipe_phv_in_data_246; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_247 = io_pipe_phv_in_data_247; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_248 = io_pipe_phv_in_data_248; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_249 = io_pipe_phv_in_data_249; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_250 = io_pipe_phv_in_data_250; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_251 = io_pipe_phv_in_data_251; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_252 = io_pipe_phv_in_data_252; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_253 = io_pipe_phv_in_data_253; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_254 = io_pipe_phv_in_data_254; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_255 = io_pipe_phv_in_data_255; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_256 = io_pipe_phv_in_data_256; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_257 = io_pipe_phv_in_data_257; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_258 = io_pipe_phv_in_data_258; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_259 = io_pipe_phv_in_data_259; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_260 = io_pipe_phv_in_data_260; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_261 = io_pipe_phv_in_data_261; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_262 = io_pipe_phv_in_data_262; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_263 = io_pipe_phv_in_data_263; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_264 = io_pipe_phv_in_data_264; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_265 = io_pipe_phv_in_data_265; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_266 = io_pipe_phv_in_data_266; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_267 = io_pipe_phv_in_data_267; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_268 = io_pipe_phv_in_data_268; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_269 = io_pipe_phv_in_data_269; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_270 = io_pipe_phv_in_data_270; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_271 = io_pipe_phv_in_data_271; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_272 = io_pipe_phv_in_data_272; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_273 = io_pipe_phv_in_data_273; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_274 = io_pipe_phv_in_data_274; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_275 = io_pipe_phv_in_data_275; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_276 = io_pipe_phv_in_data_276; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_277 = io_pipe_phv_in_data_277; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_278 = io_pipe_phv_in_data_278; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_279 = io_pipe_phv_in_data_279; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_280 = io_pipe_phv_in_data_280; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_281 = io_pipe_phv_in_data_281; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_282 = io_pipe_phv_in_data_282; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_283 = io_pipe_phv_in_data_283; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_284 = io_pipe_phv_in_data_284; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_285 = io_pipe_phv_in_data_285; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_286 = io_pipe_phv_in_data_286; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_287 = io_pipe_phv_in_data_287; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_288 = io_pipe_phv_in_data_288; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_289 = io_pipe_phv_in_data_289; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_290 = io_pipe_phv_in_data_290; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_291 = io_pipe_phv_in_data_291; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_292 = io_pipe_phv_in_data_292; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_293 = io_pipe_phv_in_data_293; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_294 = io_pipe_phv_in_data_294; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_295 = io_pipe_phv_in_data_295; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_296 = io_pipe_phv_in_data_296; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_297 = io_pipe_phv_in_data_297; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_298 = io_pipe_phv_in_data_298; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_299 = io_pipe_phv_in_data_299; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_300 = io_pipe_phv_in_data_300; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_301 = io_pipe_phv_in_data_301; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_302 = io_pipe_phv_in_data_302; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_303 = io_pipe_phv_in_data_303; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_304 = io_pipe_phv_in_data_304; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_305 = io_pipe_phv_in_data_305; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_306 = io_pipe_phv_in_data_306; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_307 = io_pipe_phv_in_data_307; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_308 = io_pipe_phv_in_data_308; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_309 = io_pipe_phv_in_data_309; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_310 = io_pipe_phv_in_data_310; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_311 = io_pipe_phv_in_data_311; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_312 = io_pipe_phv_in_data_312; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_313 = io_pipe_phv_in_data_313; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_314 = io_pipe_phv_in_data_314; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_315 = io_pipe_phv_in_data_315; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_316 = io_pipe_phv_in_data_316; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_317 = io_pipe_phv_in_data_317; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_318 = io_pipe_phv_in_data_318; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_319 = io_pipe_phv_in_data_319; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_320 = io_pipe_phv_in_data_320; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_321 = io_pipe_phv_in_data_321; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_322 = io_pipe_phv_in_data_322; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_323 = io_pipe_phv_in_data_323; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_324 = io_pipe_phv_in_data_324; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_325 = io_pipe_phv_in_data_325; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_326 = io_pipe_phv_in_data_326; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_327 = io_pipe_phv_in_data_327; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_328 = io_pipe_phv_in_data_328; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_329 = io_pipe_phv_in_data_329; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_330 = io_pipe_phv_in_data_330; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_331 = io_pipe_phv_in_data_331; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_332 = io_pipe_phv_in_data_332; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_333 = io_pipe_phv_in_data_333; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_334 = io_pipe_phv_in_data_334; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_335 = io_pipe_phv_in_data_335; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_336 = io_pipe_phv_in_data_336; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_337 = io_pipe_phv_in_data_337; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_338 = io_pipe_phv_in_data_338; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_339 = io_pipe_phv_in_data_339; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_340 = io_pipe_phv_in_data_340; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_341 = io_pipe_phv_in_data_341; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_342 = io_pipe_phv_in_data_342; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_343 = io_pipe_phv_in_data_343; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_344 = io_pipe_phv_in_data_344; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_345 = io_pipe_phv_in_data_345; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_346 = io_pipe_phv_in_data_346; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_347 = io_pipe_phv_in_data_347; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_348 = io_pipe_phv_in_data_348; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_349 = io_pipe_phv_in_data_349; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_350 = io_pipe_phv_in_data_350; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_351 = io_pipe_phv_in_data_351; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_352 = io_pipe_phv_in_data_352; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_353 = io_pipe_phv_in_data_353; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_354 = io_pipe_phv_in_data_354; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_355 = io_pipe_phv_in_data_355; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_356 = io_pipe_phv_in_data_356; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_357 = io_pipe_phv_in_data_357; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_358 = io_pipe_phv_in_data_358; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_359 = io_pipe_phv_in_data_359; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_360 = io_pipe_phv_in_data_360; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_361 = io_pipe_phv_in_data_361; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_362 = io_pipe_phv_in_data_362; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_363 = io_pipe_phv_in_data_363; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_364 = io_pipe_phv_in_data_364; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_365 = io_pipe_phv_in_data_365; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_366 = io_pipe_phv_in_data_366; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_367 = io_pipe_phv_in_data_367; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_368 = io_pipe_phv_in_data_368; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_369 = io_pipe_phv_in_data_369; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_370 = io_pipe_phv_in_data_370; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_371 = io_pipe_phv_in_data_371; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_372 = io_pipe_phv_in_data_372; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_373 = io_pipe_phv_in_data_373; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_374 = io_pipe_phv_in_data_374; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_375 = io_pipe_phv_in_data_375; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_376 = io_pipe_phv_in_data_376; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_377 = io_pipe_phv_in_data_377; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_378 = io_pipe_phv_in_data_378; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_379 = io_pipe_phv_in_data_379; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_380 = io_pipe_phv_in_data_380; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_381 = io_pipe_phv_in_data_381; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_382 = io_pipe_phv_in_data_382; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_383 = io_pipe_phv_in_data_383; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_384 = io_pipe_phv_in_data_384; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_385 = io_pipe_phv_in_data_385; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_386 = io_pipe_phv_in_data_386; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_387 = io_pipe_phv_in_data_387; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_388 = io_pipe_phv_in_data_388; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_389 = io_pipe_phv_in_data_389; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_390 = io_pipe_phv_in_data_390; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_391 = io_pipe_phv_in_data_391; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_392 = io_pipe_phv_in_data_392; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_393 = io_pipe_phv_in_data_393; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_394 = io_pipe_phv_in_data_394; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_395 = io_pipe_phv_in_data_395; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_396 = io_pipe_phv_in_data_396; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_397 = io_pipe_phv_in_data_397; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_398 = io_pipe_phv_in_data_398; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_399 = io_pipe_phv_in_data_399; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_400 = io_pipe_phv_in_data_400; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_401 = io_pipe_phv_in_data_401; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_402 = io_pipe_phv_in_data_402; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_403 = io_pipe_phv_in_data_403; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_404 = io_pipe_phv_in_data_404; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_405 = io_pipe_phv_in_data_405; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_406 = io_pipe_phv_in_data_406; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_407 = io_pipe_phv_in_data_407; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_408 = io_pipe_phv_in_data_408; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_409 = io_pipe_phv_in_data_409; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_410 = io_pipe_phv_in_data_410; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_411 = io_pipe_phv_in_data_411; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_412 = io_pipe_phv_in_data_412; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_413 = io_pipe_phv_in_data_413; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_414 = io_pipe_phv_in_data_414; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_415 = io_pipe_phv_in_data_415; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_416 = io_pipe_phv_in_data_416; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_417 = io_pipe_phv_in_data_417; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_418 = io_pipe_phv_in_data_418; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_419 = io_pipe_phv_in_data_419; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_420 = io_pipe_phv_in_data_420; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_421 = io_pipe_phv_in_data_421; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_422 = io_pipe_phv_in_data_422; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_423 = io_pipe_phv_in_data_423; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_424 = io_pipe_phv_in_data_424; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_425 = io_pipe_phv_in_data_425; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_426 = io_pipe_phv_in_data_426; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_427 = io_pipe_phv_in_data_427; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_428 = io_pipe_phv_in_data_428; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_429 = io_pipe_phv_in_data_429; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_430 = io_pipe_phv_in_data_430; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_431 = io_pipe_phv_in_data_431; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_432 = io_pipe_phv_in_data_432; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_433 = io_pipe_phv_in_data_433; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_434 = io_pipe_phv_in_data_434; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_435 = io_pipe_phv_in_data_435; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_436 = io_pipe_phv_in_data_436; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_437 = io_pipe_phv_in_data_437; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_438 = io_pipe_phv_in_data_438; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_439 = io_pipe_phv_in_data_439; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_440 = io_pipe_phv_in_data_440; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_441 = io_pipe_phv_in_data_441; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_442 = io_pipe_phv_in_data_442; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_443 = io_pipe_phv_in_data_443; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_444 = io_pipe_phv_in_data_444; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_445 = io_pipe_phv_in_data_445; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_446 = io_pipe_phv_in_data_446; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_447 = io_pipe_phv_in_data_447; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_448 = io_pipe_phv_in_data_448; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_449 = io_pipe_phv_in_data_449; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_450 = io_pipe_phv_in_data_450; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_451 = io_pipe_phv_in_data_451; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_452 = io_pipe_phv_in_data_452; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_453 = io_pipe_phv_in_data_453; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_454 = io_pipe_phv_in_data_454; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_455 = io_pipe_phv_in_data_455; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_456 = io_pipe_phv_in_data_456; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_457 = io_pipe_phv_in_data_457; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_458 = io_pipe_phv_in_data_458; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_459 = io_pipe_phv_in_data_459; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_460 = io_pipe_phv_in_data_460; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_461 = io_pipe_phv_in_data_461; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_462 = io_pipe_phv_in_data_462; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_463 = io_pipe_phv_in_data_463; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_464 = io_pipe_phv_in_data_464; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_465 = io_pipe_phv_in_data_465; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_466 = io_pipe_phv_in_data_466; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_467 = io_pipe_phv_in_data_467; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_468 = io_pipe_phv_in_data_468; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_469 = io_pipe_phv_in_data_469; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_470 = io_pipe_phv_in_data_470; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_471 = io_pipe_phv_in_data_471; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_472 = io_pipe_phv_in_data_472; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_473 = io_pipe_phv_in_data_473; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_474 = io_pipe_phv_in_data_474; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_475 = io_pipe_phv_in_data_475; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_476 = io_pipe_phv_in_data_476; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_477 = io_pipe_phv_in_data_477; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_478 = io_pipe_phv_in_data_478; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_479 = io_pipe_phv_in_data_479; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_480 = io_pipe_phv_in_data_480; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_481 = io_pipe_phv_in_data_481; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_482 = io_pipe_phv_in_data_482; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_483 = io_pipe_phv_in_data_483; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_484 = io_pipe_phv_in_data_484; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_485 = io_pipe_phv_in_data_485; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_486 = io_pipe_phv_in_data_486; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_487 = io_pipe_phv_in_data_487; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_488 = io_pipe_phv_in_data_488; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_489 = io_pipe_phv_in_data_489; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_490 = io_pipe_phv_in_data_490; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_491 = io_pipe_phv_in_data_491; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_492 = io_pipe_phv_in_data_492; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_493 = io_pipe_phv_in_data_493; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_494 = io_pipe_phv_in_data_494; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_495 = io_pipe_phv_in_data_495; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_496 = io_pipe_phv_in_data_496; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_497 = io_pipe_phv_in_data_497; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_498 = io_pipe_phv_in_data_498; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_499 = io_pipe_phv_in_data_499; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_500 = io_pipe_phv_in_data_500; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_501 = io_pipe_phv_in_data_501; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_502 = io_pipe_phv_in_data_502; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_503 = io_pipe_phv_in_data_503; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_504 = io_pipe_phv_in_data_504; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_505 = io_pipe_phv_in_data_505; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_506 = io_pipe_phv_in_data_506; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_507 = io_pipe_phv_in_data_507; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_508 = io_pipe_phv_in_data_508; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_509 = io_pipe_phv_in_data_509; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_510 = io_pipe_phv_in_data_510; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_511 = io_pipe_phv_in_data_511; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[processor.scala 17:24]
  assign PAR_io_mod_en = io_mod_par_mod_en; // @[processor.scala 18:24]
  assign PAR_io_mod_last_mau_id_mod = io_mod_par_mod_last_mau_id_mod; // @[processor.scala 18:24]
  assign PAR_io_mod_last_mau_id = io_mod_par_mod_last_mau_id; // @[processor.scala 18:24]
  assign PAR_io_mod_cs = io_mod_par_mod_cs; // @[processor.scala 18:24]
  assign PAR_io_mod_module_mod_state_id_mod = io_mod_par_mod_module_mod_state_id_mod; // @[processor.scala 18:24]
  assign PAR_io_mod_module_mod_state_id = io_mod_par_mod_module_mod_state_id; // @[processor.scala 18:24]
  assign PAR_io_mod_module_mod_sram_w_cs = io_mod_par_mod_module_mod_sram_w_cs; // @[processor.scala 18:24]
  assign PAR_io_mod_module_mod_sram_w_en = io_mod_par_mod_module_mod_sram_w_en; // @[processor.scala 18:24]
  assign PAR_io_mod_module_mod_sram_w_addr = io_mod_par_mod_module_mod_sram_w_addr; // @[processor.scala 18:24]
  assign PAR_io_mod_module_mod_sram_w_data = io_mod_par_mod_module_mod_sram_w_data; // @[processor.scala 18:24]
  assign MAT_clock = clock;
  assign MAT_io_pipe_phv_in_data_0 = PAR_io_pipe_phv_out_data_0; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_1 = PAR_io_pipe_phv_out_data_1; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_2 = PAR_io_pipe_phv_out_data_2; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_3 = PAR_io_pipe_phv_out_data_3; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_4 = PAR_io_pipe_phv_out_data_4; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_5 = PAR_io_pipe_phv_out_data_5; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_6 = PAR_io_pipe_phv_out_data_6; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_7 = PAR_io_pipe_phv_out_data_7; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_8 = PAR_io_pipe_phv_out_data_8; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_9 = PAR_io_pipe_phv_out_data_9; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_10 = PAR_io_pipe_phv_out_data_10; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_11 = PAR_io_pipe_phv_out_data_11; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_12 = PAR_io_pipe_phv_out_data_12; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_13 = PAR_io_pipe_phv_out_data_13; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_14 = PAR_io_pipe_phv_out_data_14; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_15 = PAR_io_pipe_phv_out_data_15; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_16 = PAR_io_pipe_phv_out_data_16; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_17 = PAR_io_pipe_phv_out_data_17; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_18 = PAR_io_pipe_phv_out_data_18; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_19 = PAR_io_pipe_phv_out_data_19; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_20 = PAR_io_pipe_phv_out_data_20; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_21 = PAR_io_pipe_phv_out_data_21; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_22 = PAR_io_pipe_phv_out_data_22; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_23 = PAR_io_pipe_phv_out_data_23; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_24 = PAR_io_pipe_phv_out_data_24; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_25 = PAR_io_pipe_phv_out_data_25; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_26 = PAR_io_pipe_phv_out_data_26; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_27 = PAR_io_pipe_phv_out_data_27; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_28 = PAR_io_pipe_phv_out_data_28; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_29 = PAR_io_pipe_phv_out_data_29; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_30 = PAR_io_pipe_phv_out_data_30; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_31 = PAR_io_pipe_phv_out_data_31; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_32 = PAR_io_pipe_phv_out_data_32; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_33 = PAR_io_pipe_phv_out_data_33; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_34 = PAR_io_pipe_phv_out_data_34; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_35 = PAR_io_pipe_phv_out_data_35; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_36 = PAR_io_pipe_phv_out_data_36; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_37 = PAR_io_pipe_phv_out_data_37; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_38 = PAR_io_pipe_phv_out_data_38; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_39 = PAR_io_pipe_phv_out_data_39; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_40 = PAR_io_pipe_phv_out_data_40; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_41 = PAR_io_pipe_phv_out_data_41; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_42 = PAR_io_pipe_phv_out_data_42; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_43 = PAR_io_pipe_phv_out_data_43; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_44 = PAR_io_pipe_phv_out_data_44; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_45 = PAR_io_pipe_phv_out_data_45; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_46 = PAR_io_pipe_phv_out_data_46; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_47 = PAR_io_pipe_phv_out_data_47; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_48 = PAR_io_pipe_phv_out_data_48; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_49 = PAR_io_pipe_phv_out_data_49; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_50 = PAR_io_pipe_phv_out_data_50; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_51 = PAR_io_pipe_phv_out_data_51; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_52 = PAR_io_pipe_phv_out_data_52; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_53 = PAR_io_pipe_phv_out_data_53; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_54 = PAR_io_pipe_phv_out_data_54; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_55 = PAR_io_pipe_phv_out_data_55; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_56 = PAR_io_pipe_phv_out_data_56; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_57 = PAR_io_pipe_phv_out_data_57; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_58 = PAR_io_pipe_phv_out_data_58; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_59 = PAR_io_pipe_phv_out_data_59; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_60 = PAR_io_pipe_phv_out_data_60; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_61 = PAR_io_pipe_phv_out_data_61; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_62 = PAR_io_pipe_phv_out_data_62; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_63 = PAR_io_pipe_phv_out_data_63; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_64 = PAR_io_pipe_phv_out_data_64; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_65 = PAR_io_pipe_phv_out_data_65; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_66 = PAR_io_pipe_phv_out_data_66; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_67 = PAR_io_pipe_phv_out_data_67; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_68 = PAR_io_pipe_phv_out_data_68; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_69 = PAR_io_pipe_phv_out_data_69; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_70 = PAR_io_pipe_phv_out_data_70; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_71 = PAR_io_pipe_phv_out_data_71; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_72 = PAR_io_pipe_phv_out_data_72; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_73 = PAR_io_pipe_phv_out_data_73; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_74 = PAR_io_pipe_phv_out_data_74; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_75 = PAR_io_pipe_phv_out_data_75; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_76 = PAR_io_pipe_phv_out_data_76; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_77 = PAR_io_pipe_phv_out_data_77; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_78 = PAR_io_pipe_phv_out_data_78; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_79 = PAR_io_pipe_phv_out_data_79; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_80 = PAR_io_pipe_phv_out_data_80; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_81 = PAR_io_pipe_phv_out_data_81; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_82 = PAR_io_pipe_phv_out_data_82; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_83 = PAR_io_pipe_phv_out_data_83; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_84 = PAR_io_pipe_phv_out_data_84; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_85 = PAR_io_pipe_phv_out_data_85; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_86 = PAR_io_pipe_phv_out_data_86; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_87 = PAR_io_pipe_phv_out_data_87; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_88 = PAR_io_pipe_phv_out_data_88; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_89 = PAR_io_pipe_phv_out_data_89; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_90 = PAR_io_pipe_phv_out_data_90; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_91 = PAR_io_pipe_phv_out_data_91; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_92 = PAR_io_pipe_phv_out_data_92; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_93 = PAR_io_pipe_phv_out_data_93; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_94 = PAR_io_pipe_phv_out_data_94; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_95 = PAR_io_pipe_phv_out_data_95; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_96 = PAR_io_pipe_phv_out_data_96; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_97 = PAR_io_pipe_phv_out_data_97; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_98 = PAR_io_pipe_phv_out_data_98; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_99 = PAR_io_pipe_phv_out_data_99; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_100 = PAR_io_pipe_phv_out_data_100; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_101 = PAR_io_pipe_phv_out_data_101; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_102 = PAR_io_pipe_phv_out_data_102; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_103 = PAR_io_pipe_phv_out_data_103; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_104 = PAR_io_pipe_phv_out_data_104; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_105 = PAR_io_pipe_phv_out_data_105; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_106 = PAR_io_pipe_phv_out_data_106; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_107 = PAR_io_pipe_phv_out_data_107; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_108 = PAR_io_pipe_phv_out_data_108; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_109 = PAR_io_pipe_phv_out_data_109; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_110 = PAR_io_pipe_phv_out_data_110; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_111 = PAR_io_pipe_phv_out_data_111; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_112 = PAR_io_pipe_phv_out_data_112; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_113 = PAR_io_pipe_phv_out_data_113; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_114 = PAR_io_pipe_phv_out_data_114; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_115 = PAR_io_pipe_phv_out_data_115; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_116 = PAR_io_pipe_phv_out_data_116; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_117 = PAR_io_pipe_phv_out_data_117; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_118 = PAR_io_pipe_phv_out_data_118; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_119 = PAR_io_pipe_phv_out_data_119; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_120 = PAR_io_pipe_phv_out_data_120; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_121 = PAR_io_pipe_phv_out_data_121; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_122 = PAR_io_pipe_phv_out_data_122; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_123 = PAR_io_pipe_phv_out_data_123; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_124 = PAR_io_pipe_phv_out_data_124; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_125 = PAR_io_pipe_phv_out_data_125; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_126 = PAR_io_pipe_phv_out_data_126; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_127 = PAR_io_pipe_phv_out_data_127; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_128 = PAR_io_pipe_phv_out_data_128; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_129 = PAR_io_pipe_phv_out_data_129; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_130 = PAR_io_pipe_phv_out_data_130; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_131 = PAR_io_pipe_phv_out_data_131; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_132 = PAR_io_pipe_phv_out_data_132; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_133 = PAR_io_pipe_phv_out_data_133; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_134 = PAR_io_pipe_phv_out_data_134; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_135 = PAR_io_pipe_phv_out_data_135; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_136 = PAR_io_pipe_phv_out_data_136; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_137 = PAR_io_pipe_phv_out_data_137; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_138 = PAR_io_pipe_phv_out_data_138; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_139 = PAR_io_pipe_phv_out_data_139; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_140 = PAR_io_pipe_phv_out_data_140; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_141 = PAR_io_pipe_phv_out_data_141; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_142 = PAR_io_pipe_phv_out_data_142; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_143 = PAR_io_pipe_phv_out_data_143; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_144 = PAR_io_pipe_phv_out_data_144; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_145 = PAR_io_pipe_phv_out_data_145; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_146 = PAR_io_pipe_phv_out_data_146; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_147 = PAR_io_pipe_phv_out_data_147; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_148 = PAR_io_pipe_phv_out_data_148; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_149 = PAR_io_pipe_phv_out_data_149; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_150 = PAR_io_pipe_phv_out_data_150; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_151 = PAR_io_pipe_phv_out_data_151; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_152 = PAR_io_pipe_phv_out_data_152; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_153 = PAR_io_pipe_phv_out_data_153; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_154 = PAR_io_pipe_phv_out_data_154; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_155 = PAR_io_pipe_phv_out_data_155; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_156 = PAR_io_pipe_phv_out_data_156; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_157 = PAR_io_pipe_phv_out_data_157; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_158 = PAR_io_pipe_phv_out_data_158; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_159 = PAR_io_pipe_phv_out_data_159; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_160 = PAR_io_pipe_phv_out_data_160; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_161 = PAR_io_pipe_phv_out_data_161; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_162 = PAR_io_pipe_phv_out_data_162; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_163 = PAR_io_pipe_phv_out_data_163; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_164 = PAR_io_pipe_phv_out_data_164; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_165 = PAR_io_pipe_phv_out_data_165; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_166 = PAR_io_pipe_phv_out_data_166; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_167 = PAR_io_pipe_phv_out_data_167; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_168 = PAR_io_pipe_phv_out_data_168; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_169 = PAR_io_pipe_phv_out_data_169; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_170 = PAR_io_pipe_phv_out_data_170; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_171 = PAR_io_pipe_phv_out_data_171; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_172 = PAR_io_pipe_phv_out_data_172; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_173 = PAR_io_pipe_phv_out_data_173; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_174 = PAR_io_pipe_phv_out_data_174; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_175 = PAR_io_pipe_phv_out_data_175; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_176 = PAR_io_pipe_phv_out_data_176; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_177 = PAR_io_pipe_phv_out_data_177; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_178 = PAR_io_pipe_phv_out_data_178; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_179 = PAR_io_pipe_phv_out_data_179; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_180 = PAR_io_pipe_phv_out_data_180; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_181 = PAR_io_pipe_phv_out_data_181; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_182 = PAR_io_pipe_phv_out_data_182; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_183 = PAR_io_pipe_phv_out_data_183; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_184 = PAR_io_pipe_phv_out_data_184; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_185 = PAR_io_pipe_phv_out_data_185; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_186 = PAR_io_pipe_phv_out_data_186; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_187 = PAR_io_pipe_phv_out_data_187; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_188 = PAR_io_pipe_phv_out_data_188; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_189 = PAR_io_pipe_phv_out_data_189; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_190 = PAR_io_pipe_phv_out_data_190; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_191 = PAR_io_pipe_phv_out_data_191; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_192 = PAR_io_pipe_phv_out_data_192; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_193 = PAR_io_pipe_phv_out_data_193; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_194 = PAR_io_pipe_phv_out_data_194; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_195 = PAR_io_pipe_phv_out_data_195; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_196 = PAR_io_pipe_phv_out_data_196; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_197 = PAR_io_pipe_phv_out_data_197; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_198 = PAR_io_pipe_phv_out_data_198; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_199 = PAR_io_pipe_phv_out_data_199; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_200 = PAR_io_pipe_phv_out_data_200; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_201 = PAR_io_pipe_phv_out_data_201; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_202 = PAR_io_pipe_phv_out_data_202; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_203 = PAR_io_pipe_phv_out_data_203; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_204 = PAR_io_pipe_phv_out_data_204; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_205 = PAR_io_pipe_phv_out_data_205; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_206 = PAR_io_pipe_phv_out_data_206; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_207 = PAR_io_pipe_phv_out_data_207; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_208 = PAR_io_pipe_phv_out_data_208; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_209 = PAR_io_pipe_phv_out_data_209; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_210 = PAR_io_pipe_phv_out_data_210; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_211 = PAR_io_pipe_phv_out_data_211; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_212 = PAR_io_pipe_phv_out_data_212; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_213 = PAR_io_pipe_phv_out_data_213; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_214 = PAR_io_pipe_phv_out_data_214; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_215 = PAR_io_pipe_phv_out_data_215; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_216 = PAR_io_pipe_phv_out_data_216; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_217 = PAR_io_pipe_phv_out_data_217; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_218 = PAR_io_pipe_phv_out_data_218; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_219 = PAR_io_pipe_phv_out_data_219; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_220 = PAR_io_pipe_phv_out_data_220; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_221 = PAR_io_pipe_phv_out_data_221; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_222 = PAR_io_pipe_phv_out_data_222; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_223 = PAR_io_pipe_phv_out_data_223; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_224 = PAR_io_pipe_phv_out_data_224; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_225 = PAR_io_pipe_phv_out_data_225; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_226 = PAR_io_pipe_phv_out_data_226; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_227 = PAR_io_pipe_phv_out_data_227; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_228 = PAR_io_pipe_phv_out_data_228; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_229 = PAR_io_pipe_phv_out_data_229; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_230 = PAR_io_pipe_phv_out_data_230; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_231 = PAR_io_pipe_phv_out_data_231; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_232 = PAR_io_pipe_phv_out_data_232; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_233 = PAR_io_pipe_phv_out_data_233; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_234 = PAR_io_pipe_phv_out_data_234; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_235 = PAR_io_pipe_phv_out_data_235; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_236 = PAR_io_pipe_phv_out_data_236; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_237 = PAR_io_pipe_phv_out_data_237; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_238 = PAR_io_pipe_phv_out_data_238; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_239 = PAR_io_pipe_phv_out_data_239; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_240 = PAR_io_pipe_phv_out_data_240; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_241 = PAR_io_pipe_phv_out_data_241; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_242 = PAR_io_pipe_phv_out_data_242; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_243 = PAR_io_pipe_phv_out_data_243; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_244 = PAR_io_pipe_phv_out_data_244; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_245 = PAR_io_pipe_phv_out_data_245; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_246 = PAR_io_pipe_phv_out_data_246; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_247 = PAR_io_pipe_phv_out_data_247; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_248 = PAR_io_pipe_phv_out_data_248; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_249 = PAR_io_pipe_phv_out_data_249; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_250 = PAR_io_pipe_phv_out_data_250; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_251 = PAR_io_pipe_phv_out_data_251; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_252 = PAR_io_pipe_phv_out_data_252; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_253 = PAR_io_pipe_phv_out_data_253; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_254 = PAR_io_pipe_phv_out_data_254; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_255 = PAR_io_pipe_phv_out_data_255; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_256 = PAR_io_pipe_phv_out_data_256; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_257 = PAR_io_pipe_phv_out_data_257; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_258 = PAR_io_pipe_phv_out_data_258; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_259 = PAR_io_pipe_phv_out_data_259; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_260 = PAR_io_pipe_phv_out_data_260; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_261 = PAR_io_pipe_phv_out_data_261; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_262 = PAR_io_pipe_phv_out_data_262; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_263 = PAR_io_pipe_phv_out_data_263; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_264 = PAR_io_pipe_phv_out_data_264; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_265 = PAR_io_pipe_phv_out_data_265; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_266 = PAR_io_pipe_phv_out_data_266; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_267 = PAR_io_pipe_phv_out_data_267; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_268 = PAR_io_pipe_phv_out_data_268; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_269 = PAR_io_pipe_phv_out_data_269; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_270 = PAR_io_pipe_phv_out_data_270; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_271 = PAR_io_pipe_phv_out_data_271; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_272 = PAR_io_pipe_phv_out_data_272; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_273 = PAR_io_pipe_phv_out_data_273; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_274 = PAR_io_pipe_phv_out_data_274; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_275 = PAR_io_pipe_phv_out_data_275; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_276 = PAR_io_pipe_phv_out_data_276; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_277 = PAR_io_pipe_phv_out_data_277; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_278 = PAR_io_pipe_phv_out_data_278; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_279 = PAR_io_pipe_phv_out_data_279; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_280 = PAR_io_pipe_phv_out_data_280; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_281 = PAR_io_pipe_phv_out_data_281; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_282 = PAR_io_pipe_phv_out_data_282; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_283 = PAR_io_pipe_phv_out_data_283; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_284 = PAR_io_pipe_phv_out_data_284; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_285 = PAR_io_pipe_phv_out_data_285; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_286 = PAR_io_pipe_phv_out_data_286; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_287 = PAR_io_pipe_phv_out_data_287; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_288 = PAR_io_pipe_phv_out_data_288; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_289 = PAR_io_pipe_phv_out_data_289; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_290 = PAR_io_pipe_phv_out_data_290; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_291 = PAR_io_pipe_phv_out_data_291; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_292 = PAR_io_pipe_phv_out_data_292; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_293 = PAR_io_pipe_phv_out_data_293; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_294 = PAR_io_pipe_phv_out_data_294; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_295 = PAR_io_pipe_phv_out_data_295; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_296 = PAR_io_pipe_phv_out_data_296; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_297 = PAR_io_pipe_phv_out_data_297; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_298 = PAR_io_pipe_phv_out_data_298; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_299 = PAR_io_pipe_phv_out_data_299; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_300 = PAR_io_pipe_phv_out_data_300; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_301 = PAR_io_pipe_phv_out_data_301; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_302 = PAR_io_pipe_phv_out_data_302; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_303 = PAR_io_pipe_phv_out_data_303; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_304 = PAR_io_pipe_phv_out_data_304; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_305 = PAR_io_pipe_phv_out_data_305; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_306 = PAR_io_pipe_phv_out_data_306; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_307 = PAR_io_pipe_phv_out_data_307; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_308 = PAR_io_pipe_phv_out_data_308; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_309 = PAR_io_pipe_phv_out_data_309; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_310 = PAR_io_pipe_phv_out_data_310; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_311 = PAR_io_pipe_phv_out_data_311; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_312 = PAR_io_pipe_phv_out_data_312; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_313 = PAR_io_pipe_phv_out_data_313; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_314 = PAR_io_pipe_phv_out_data_314; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_315 = PAR_io_pipe_phv_out_data_315; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_316 = PAR_io_pipe_phv_out_data_316; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_317 = PAR_io_pipe_phv_out_data_317; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_318 = PAR_io_pipe_phv_out_data_318; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_319 = PAR_io_pipe_phv_out_data_319; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_320 = PAR_io_pipe_phv_out_data_320; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_321 = PAR_io_pipe_phv_out_data_321; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_322 = PAR_io_pipe_phv_out_data_322; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_323 = PAR_io_pipe_phv_out_data_323; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_324 = PAR_io_pipe_phv_out_data_324; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_325 = PAR_io_pipe_phv_out_data_325; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_326 = PAR_io_pipe_phv_out_data_326; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_327 = PAR_io_pipe_phv_out_data_327; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_328 = PAR_io_pipe_phv_out_data_328; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_329 = PAR_io_pipe_phv_out_data_329; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_330 = PAR_io_pipe_phv_out_data_330; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_331 = PAR_io_pipe_phv_out_data_331; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_332 = PAR_io_pipe_phv_out_data_332; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_333 = PAR_io_pipe_phv_out_data_333; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_334 = PAR_io_pipe_phv_out_data_334; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_335 = PAR_io_pipe_phv_out_data_335; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_336 = PAR_io_pipe_phv_out_data_336; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_337 = PAR_io_pipe_phv_out_data_337; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_338 = PAR_io_pipe_phv_out_data_338; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_339 = PAR_io_pipe_phv_out_data_339; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_340 = PAR_io_pipe_phv_out_data_340; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_341 = PAR_io_pipe_phv_out_data_341; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_342 = PAR_io_pipe_phv_out_data_342; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_343 = PAR_io_pipe_phv_out_data_343; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_344 = PAR_io_pipe_phv_out_data_344; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_345 = PAR_io_pipe_phv_out_data_345; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_346 = PAR_io_pipe_phv_out_data_346; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_347 = PAR_io_pipe_phv_out_data_347; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_348 = PAR_io_pipe_phv_out_data_348; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_349 = PAR_io_pipe_phv_out_data_349; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_350 = PAR_io_pipe_phv_out_data_350; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_351 = PAR_io_pipe_phv_out_data_351; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_352 = PAR_io_pipe_phv_out_data_352; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_353 = PAR_io_pipe_phv_out_data_353; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_354 = PAR_io_pipe_phv_out_data_354; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_355 = PAR_io_pipe_phv_out_data_355; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_356 = PAR_io_pipe_phv_out_data_356; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_357 = PAR_io_pipe_phv_out_data_357; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_358 = PAR_io_pipe_phv_out_data_358; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_359 = PAR_io_pipe_phv_out_data_359; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_360 = PAR_io_pipe_phv_out_data_360; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_361 = PAR_io_pipe_phv_out_data_361; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_362 = PAR_io_pipe_phv_out_data_362; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_363 = PAR_io_pipe_phv_out_data_363; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_364 = PAR_io_pipe_phv_out_data_364; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_365 = PAR_io_pipe_phv_out_data_365; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_366 = PAR_io_pipe_phv_out_data_366; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_367 = PAR_io_pipe_phv_out_data_367; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_368 = PAR_io_pipe_phv_out_data_368; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_369 = PAR_io_pipe_phv_out_data_369; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_370 = PAR_io_pipe_phv_out_data_370; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_371 = PAR_io_pipe_phv_out_data_371; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_372 = PAR_io_pipe_phv_out_data_372; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_373 = PAR_io_pipe_phv_out_data_373; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_374 = PAR_io_pipe_phv_out_data_374; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_375 = PAR_io_pipe_phv_out_data_375; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_376 = PAR_io_pipe_phv_out_data_376; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_377 = PAR_io_pipe_phv_out_data_377; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_378 = PAR_io_pipe_phv_out_data_378; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_379 = PAR_io_pipe_phv_out_data_379; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_380 = PAR_io_pipe_phv_out_data_380; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_381 = PAR_io_pipe_phv_out_data_381; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_382 = PAR_io_pipe_phv_out_data_382; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_383 = PAR_io_pipe_phv_out_data_383; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_384 = PAR_io_pipe_phv_out_data_384; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_385 = PAR_io_pipe_phv_out_data_385; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_386 = PAR_io_pipe_phv_out_data_386; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_387 = PAR_io_pipe_phv_out_data_387; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_388 = PAR_io_pipe_phv_out_data_388; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_389 = PAR_io_pipe_phv_out_data_389; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_390 = PAR_io_pipe_phv_out_data_390; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_391 = PAR_io_pipe_phv_out_data_391; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_392 = PAR_io_pipe_phv_out_data_392; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_393 = PAR_io_pipe_phv_out_data_393; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_394 = PAR_io_pipe_phv_out_data_394; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_395 = PAR_io_pipe_phv_out_data_395; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_396 = PAR_io_pipe_phv_out_data_396; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_397 = PAR_io_pipe_phv_out_data_397; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_398 = PAR_io_pipe_phv_out_data_398; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_399 = PAR_io_pipe_phv_out_data_399; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_400 = PAR_io_pipe_phv_out_data_400; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_401 = PAR_io_pipe_phv_out_data_401; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_402 = PAR_io_pipe_phv_out_data_402; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_403 = PAR_io_pipe_phv_out_data_403; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_404 = PAR_io_pipe_phv_out_data_404; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_405 = PAR_io_pipe_phv_out_data_405; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_406 = PAR_io_pipe_phv_out_data_406; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_407 = PAR_io_pipe_phv_out_data_407; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_408 = PAR_io_pipe_phv_out_data_408; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_409 = PAR_io_pipe_phv_out_data_409; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_410 = PAR_io_pipe_phv_out_data_410; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_411 = PAR_io_pipe_phv_out_data_411; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_412 = PAR_io_pipe_phv_out_data_412; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_413 = PAR_io_pipe_phv_out_data_413; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_414 = PAR_io_pipe_phv_out_data_414; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_415 = PAR_io_pipe_phv_out_data_415; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_416 = PAR_io_pipe_phv_out_data_416; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_417 = PAR_io_pipe_phv_out_data_417; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_418 = PAR_io_pipe_phv_out_data_418; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_419 = PAR_io_pipe_phv_out_data_419; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_420 = PAR_io_pipe_phv_out_data_420; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_421 = PAR_io_pipe_phv_out_data_421; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_422 = PAR_io_pipe_phv_out_data_422; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_423 = PAR_io_pipe_phv_out_data_423; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_424 = PAR_io_pipe_phv_out_data_424; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_425 = PAR_io_pipe_phv_out_data_425; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_426 = PAR_io_pipe_phv_out_data_426; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_427 = PAR_io_pipe_phv_out_data_427; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_428 = PAR_io_pipe_phv_out_data_428; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_429 = PAR_io_pipe_phv_out_data_429; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_430 = PAR_io_pipe_phv_out_data_430; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_431 = PAR_io_pipe_phv_out_data_431; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_432 = PAR_io_pipe_phv_out_data_432; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_433 = PAR_io_pipe_phv_out_data_433; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_434 = PAR_io_pipe_phv_out_data_434; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_435 = PAR_io_pipe_phv_out_data_435; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_436 = PAR_io_pipe_phv_out_data_436; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_437 = PAR_io_pipe_phv_out_data_437; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_438 = PAR_io_pipe_phv_out_data_438; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_439 = PAR_io_pipe_phv_out_data_439; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_440 = PAR_io_pipe_phv_out_data_440; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_441 = PAR_io_pipe_phv_out_data_441; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_442 = PAR_io_pipe_phv_out_data_442; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_443 = PAR_io_pipe_phv_out_data_443; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_444 = PAR_io_pipe_phv_out_data_444; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_445 = PAR_io_pipe_phv_out_data_445; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_446 = PAR_io_pipe_phv_out_data_446; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_447 = PAR_io_pipe_phv_out_data_447; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_448 = PAR_io_pipe_phv_out_data_448; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_449 = PAR_io_pipe_phv_out_data_449; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_450 = PAR_io_pipe_phv_out_data_450; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_451 = PAR_io_pipe_phv_out_data_451; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_452 = PAR_io_pipe_phv_out_data_452; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_453 = PAR_io_pipe_phv_out_data_453; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_454 = PAR_io_pipe_phv_out_data_454; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_455 = PAR_io_pipe_phv_out_data_455; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_456 = PAR_io_pipe_phv_out_data_456; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_457 = PAR_io_pipe_phv_out_data_457; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_458 = PAR_io_pipe_phv_out_data_458; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_459 = PAR_io_pipe_phv_out_data_459; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_460 = PAR_io_pipe_phv_out_data_460; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_461 = PAR_io_pipe_phv_out_data_461; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_462 = PAR_io_pipe_phv_out_data_462; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_463 = PAR_io_pipe_phv_out_data_463; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_464 = PAR_io_pipe_phv_out_data_464; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_465 = PAR_io_pipe_phv_out_data_465; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_466 = PAR_io_pipe_phv_out_data_466; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_467 = PAR_io_pipe_phv_out_data_467; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_468 = PAR_io_pipe_phv_out_data_468; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_469 = PAR_io_pipe_phv_out_data_469; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_470 = PAR_io_pipe_phv_out_data_470; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_471 = PAR_io_pipe_phv_out_data_471; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_472 = PAR_io_pipe_phv_out_data_472; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_473 = PAR_io_pipe_phv_out_data_473; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_474 = PAR_io_pipe_phv_out_data_474; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_475 = PAR_io_pipe_phv_out_data_475; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_476 = PAR_io_pipe_phv_out_data_476; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_477 = PAR_io_pipe_phv_out_data_477; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_478 = PAR_io_pipe_phv_out_data_478; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_479 = PAR_io_pipe_phv_out_data_479; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_480 = PAR_io_pipe_phv_out_data_480; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_481 = PAR_io_pipe_phv_out_data_481; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_482 = PAR_io_pipe_phv_out_data_482; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_483 = PAR_io_pipe_phv_out_data_483; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_484 = PAR_io_pipe_phv_out_data_484; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_485 = PAR_io_pipe_phv_out_data_485; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_486 = PAR_io_pipe_phv_out_data_486; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_487 = PAR_io_pipe_phv_out_data_487; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_488 = PAR_io_pipe_phv_out_data_488; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_489 = PAR_io_pipe_phv_out_data_489; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_490 = PAR_io_pipe_phv_out_data_490; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_491 = PAR_io_pipe_phv_out_data_491; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_492 = PAR_io_pipe_phv_out_data_492; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_493 = PAR_io_pipe_phv_out_data_493; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_494 = PAR_io_pipe_phv_out_data_494; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_495 = PAR_io_pipe_phv_out_data_495; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_496 = PAR_io_pipe_phv_out_data_496; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_497 = PAR_io_pipe_phv_out_data_497; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_498 = PAR_io_pipe_phv_out_data_498; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_499 = PAR_io_pipe_phv_out_data_499; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_500 = PAR_io_pipe_phv_out_data_500; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_501 = PAR_io_pipe_phv_out_data_501; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_502 = PAR_io_pipe_phv_out_data_502; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_503 = PAR_io_pipe_phv_out_data_503; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_504 = PAR_io_pipe_phv_out_data_504; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_505 = PAR_io_pipe_phv_out_data_505; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_506 = PAR_io_pipe_phv_out_data_506; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_507 = PAR_io_pipe_phv_out_data_507; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_508 = PAR_io_pipe_phv_out_data_508; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_509 = PAR_io_pipe_phv_out_data_509; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_510 = PAR_io_pipe_phv_out_data_510; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_511 = PAR_io_pipe_phv_out_data_511; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_0 = PAR_io_pipe_phv_out_header_0; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_1 = PAR_io_pipe_phv_out_header_1; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_2 = PAR_io_pipe_phv_out_header_2; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_3 = PAR_io_pipe_phv_out_header_3; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_4 = PAR_io_pipe_phv_out_header_4; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_5 = PAR_io_pipe_phv_out_header_5; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_6 = PAR_io_pipe_phv_out_header_6; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_7 = PAR_io_pipe_phv_out_header_7; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_8 = PAR_io_pipe_phv_out_header_8; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_9 = PAR_io_pipe_phv_out_header_9; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_10 = PAR_io_pipe_phv_out_header_10; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_11 = PAR_io_pipe_phv_out_header_11; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_12 = PAR_io_pipe_phv_out_header_12; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_13 = PAR_io_pipe_phv_out_header_13; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_14 = PAR_io_pipe_phv_out_header_14; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_15 = PAR_io_pipe_phv_out_header_15; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_parse_current_state = PAR_io_pipe_phv_out_parse_current_state; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_parse_current_offset = PAR_io_pipe_phv_out_parse_current_offset; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_parse_transition_field = PAR_io_pipe_phv_out_parse_transition_field; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_next_processor_id = PAR_io_pipe_phv_out_next_processor_id; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_next_config_id = PAR_io_pipe_phv_out_next_config_id; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_is_valid_processor = PAR_io_pipe_phv_out_is_valid_processor; // @[processor.scala 20:24]
  assign MAT_io_mod_en = io_mod_mat_mod_en; // @[processor.scala 21:24]
  assign MAT_io_mod_config_id = io_mod_mat_mod_config_id; // @[processor.scala 21:24]
  assign MAT_io_mod_key_mod_header_id = io_mod_mat_mod_key_mod_header_id; // @[processor.scala 21:24]
  assign MAT_io_mod_key_mod_internal_offset = io_mod_mat_mod_key_mod_internal_offset; // @[processor.scala 21:24]
  assign MAT_io_mod_key_mod_key_length = io_mod_mat_mod_key_mod_key_length; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_table_width = io_mod_mat_mod_table_mod_table_width; // @[processor.scala 21:24]
  assign MAT_io_mod_table_mod_table_depth = io_mod_mat_mod_table_mod_table_depth; // @[processor.scala 21:24]
  assign MAT_io_mem_cluster_0_data = io_mem_cluster_0_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_1_data = io_mem_cluster_1_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_2_data = io_mem_cluster_2_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_3_data = io_mem_cluster_3_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_4_data = io_mem_cluster_4_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_5_data = io_mem_cluster_5_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_6_data = io_mem_cluster_6_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_7_data = io_mem_cluster_7_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_8_data = io_mem_cluster_8_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_9_data = io_mem_cluster_9_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_10_data = io_mem_cluster_10_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_11_data = io_mem_cluster_11_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_12_data = io_mem_cluster_12_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_13_data = io_mem_cluster_13_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_14_data = io_mem_cluster_14_data; // @[processor.scala 22:24]
  assign MAT_io_mem_cluster_15_data = io_mem_cluster_15_data; // @[processor.scala 22:24]
  assign EXE_clock = clock;
  assign EXE_io_pipe_phv_in_data_0 = MAT_io_pipe_phv_out_data_0; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_1 = MAT_io_pipe_phv_out_data_1; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_2 = MAT_io_pipe_phv_out_data_2; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_3 = MAT_io_pipe_phv_out_data_3; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_4 = MAT_io_pipe_phv_out_data_4; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_5 = MAT_io_pipe_phv_out_data_5; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_6 = MAT_io_pipe_phv_out_data_6; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_7 = MAT_io_pipe_phv_out_data_7; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_8 = MAT_io_pipe_phv_out_data_8; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_9 = MAT_io_pipe_phv_out_data_9; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_10 = MAT_io_pipe_phv_out_data_10; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_11 = MAT_io_pipe_phv_out_data_11; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_12 = MAT_io_pipe_phv_out_data_12; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_13 = MAT_io_pipe_phv_out_data_13; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_14 = MAT_io_pipe_phv_out_data_14; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_15 = MAT_io_pipe_phv_out_data_15; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_16 = MAT_io_pipe_phv_out_data_16; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_17 = MAT_io_pipe_phv_out_data_17; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_18 = MAT_io_pipe_phv_out_data_18; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_19 = MAT_io_pipe_phv_out_data_19; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_20 = MAT_io_pipe_phv_out_data_20; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_21 = MAT_io_pipe_phv_out_data_21; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_22 = MAT_io_pipe_phv_out_data_22; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_23 = MAT_io_pipe_phv_out_data_23; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_24 = MAT_io_pipe_phv_out_data_24; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_25 = MAT_io_pipe_phv_out_data_25; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_26 = MAT_io_pipe_phv_out_data_26; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_27 = MAT_io_pipe_phv_out_data_27; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_28 = MAT_io_pipe_phv_out_data_28; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_29 = MAT_io_pipe_phv_out_data_29; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_30 = MAT_io_pipe_phv_out_data_30; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_31 = MAT_io_pipe_phv_out_data_31; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_32 = MAT_io_pipe_phv_out_data_32; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_33 = MAT_io_pipe_phv_out_data_33; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_34 = MAT_io_pipe_phv_out_data_34; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_35 = MAT_io_pipe_phv_out_data_35; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_36 = MAT_io_pipe_phv_out_data_36; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_37 = MAT_io_pipe_phv_out_data_37; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_38 = MAT_io_pipe_phv_out_data_38; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_39 = MAT_io_pipe_phv_out_data_39; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_40 = MAT_io_pipe_phv_out_data_40; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_41 = MAT_io_pipe_phv_out_data_41; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_42 = MAT_io_pipe_phv_out_data_42; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_43 = MAT_io_pipe_phv_out_data_43; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_44 = MAT_io_pipe_phv_out_data_44; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_45 = MAT_io_pipe_phv_out_data_45; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_46 = MAT_io_pipe_phv_out_data_46; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_47 = MAT_io_pipe_phv_out_data_47; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_48 = MAT_io_pipe_phv_out_data_48; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_49 = MAT_io_pipe_phv_out_data_49; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_50 = MAT_io_pipe_phv_out_data_50; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_51 = MAT_io_pipe_phv_out_data_51; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_52 = MAT_io_pipe_phv_out_data_52; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_53 = MAT_io_pipe_phv_out_data_53; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_54 = MAT_io_pipe_phv_out_data_54; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_55 = MAT_io_pipe_phv_out_data_55; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_56 = MAT_io_pipe_phv_out_data_56; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_57 = MAT_io_pipe_phv_out_data_57; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_58 = MAT_io_pipe_phv_out_data_58; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_59 = MAT_io_pipe_phv_out_data_59; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_60 = MAT_io_pipe_phv_out_data_60; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_61 = MAT_io_pipe_phv_out_data_61; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_62 = MAT_io_pipe_phv_out_data_62; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_63 = MAT_io_pipe_phv_out_data_63; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_64 = MAT_io_pipe_phv_out_data_64; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_65 = MAT_io_pipe_phv_out_data_65; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_66 = MAT_io_pipe_phv_out_data_66; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_67 = MAT_io_pipe_phv_out_data_67; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_68 = MAT_io_pipe_phv_out_data_68; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_69 = MAT_io_pipe_phv_out_data_69; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_70 = MAT_io_pipe_phv_out_data_70; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_71 = MAT_io_pipe_phv_out_data_71; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_72 = MAT_io_pipe_phv_out_data_72; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_73 = MAT_io_pipe_phv_out_data_73; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_74 = MAT_io_pipe_phv_out_data_74; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_75 = MAT_io_pipe_phv_out_data_75; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_76 = MAT_io_pipe_phv_out_data_76; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_77 = MAT_io_pipe_phv_out_data_77; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_78 = MAT_io_pipe_phv_out_data_78; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_79 = MAT_io_pipe_phv_out_data_79; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_80 = MAT_io_pipe_phv_out_data_80; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_81 = MAT_io_pipe_phv_out_data_81; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_82 = MAT_io_pipe_phv_out_data_82; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_83 = MAT_io_pipe_phv_out_data_83; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_84 = MAT_io_pipe_phv_out_data_84; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_85 = MAT_io_pipe_phv_out_data_85; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_86 = MAT_io_pipe_phv_out_data_86; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_87 = MAT_io_pipe_phv_out_data_87; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_88 = MAT_io_pipe_phv_out_data_88; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_89 = MAT_io_pipe_phv_out_data_89; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_90 = MAT_io_pipe_phv_out_data_90; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_91 = MAT_io_pipe_phv_out_data_91; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_92 = MAT_io_pipe_phv_out_data_92; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_93 = MAT_io_pipe_phv_out_data_93; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_94 = MAT_io_pipe_phv_out_data_94; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_95 = MAT_io_pipe_phv_out_data_95; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_96 = MAT_io_pipe_phv_out_data_96; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_97 = MAT_io_pipe_phv_out_data_97; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_98 = MAT_io_pipe_phv_out_data_98; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_99 = MAT_io_pipe_phv_out_data_99; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_100 = MAT_io_pipe_phv_out_data_100; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_101 = MAT_io_pipe_phv_out_data_101; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_102 = MAT_io_pipe_phv_out_data_102; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_103 = MAT_io_pipe_phv_out_data_103; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_104 = MAT_io_pipe_phv_out_data_104; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_105 = MAT_io_pipe_phv_out_data_105; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_106 = MAT_io_pipe_phv_out_data_106; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_107 = MAT_io_pipe_phv_out_data_107; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_108 = MAT_io_pipe_phv_out_data_108; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_109 = MAT_io_pipe_phv_out_data_109; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_110 = MAT_io_pipe_phv_out_data_110; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_111 = MAT_io_pipe_phv_out_data_111; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_112 = MAT_io_pipe_phv_out_data_112; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_113 = MAT_io_pipe_phv_out_data_113; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_114 = MAT_io_pipe_phv_out_data_114; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_115 = MAT_io_pipe_phv_out_data_115; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_116 = MAT_io_pipe_phv_out_data_116; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_117 = MAT_io_pipe_phv_out_data_117; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_118 = MAT_io_pipe_phv_out_data_118; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_119 = MAT_io_pipe_phv_out_data_119; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_120 = MAT_io_pipe_phv_out_data_120; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_121 = MAT_io_pipe_phv_out_data_121; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_122 = MAT_io_pipe_phv_out_data_122; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_123 = MAT_io_pipe_phv_out_data_123; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_124 = MAT_io_pipe_phv_out_data_124; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_125 = MAT_io_pipe_phv_out_data_125; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_126 = MAT_io_pipe_phv_out_data_126; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_127 = MAT_io_pipe_phv_out_data_127; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_128 = MAT_io_pipe_phv_out_data_128; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_129 = MAT_io_pipe_phv_out_data_129; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_130 = MAT_io_pipe_phv_out_data_130; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_131 = MAT_io_pipe_phv_out_data_131; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_132 = MAT_io_pipe_phv_out_data_132; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_133 = MAT_io_pipe_phv_out_data_133; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_134 = MAT_io_pipe_phv_out_data_134; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_135 = MAT_io_pipe_phv_out_data_135; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_136 = MAT_io_pipe_phv_out_data_136; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_137 = MAT_io_pipe_phv_out_data_137; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_138 = MAT_io_pipe_phv_out_data_138; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_139 = MAT_io_pipe_phv_out_data_139; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_140 = MAT_io_pipe_phv_out_data_140; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_141 = MAT_io_pipe_phv_out_data_141; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_142 = MAT_io_pipe_phv_out_data_142; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_143 = MAT_io_pipe_phv_out_data_143; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_144 = MAT_io_pipe_phv_out_data_144; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_145 = MAT_io_pipe_phv_out_data_145; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_146 = MAT_io_pipe_phv_out_data_146; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_147 = MAT_io_pipe_phv_out_data_147; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_148 = MAT_io_pipe_phv_out_data_148; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_149 = MAT_io_pipe_phv_out_data_149; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_150 = MAT_io_pipe_phv_out_data_150; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_151 = MAT_io_pipe_phv_out_data_151; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_152 = MAT_io_pipe_phv_out_data_152; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_153 = MAT_io_pipe_phv_out_data_153; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_154 = MAT_io_pipe_phv_out_data_154; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_155 = MAT_io_pipe_phv_out_data_155; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_156 = MAT_io_pipe_phv_out_data_156; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_157 = MAT_io_pipe_phv_out_data_157; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_158 = MAT_io_pipe_phv_out_data_158; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_159 = MAT_io_pipe_phv_out_data_159; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_160 = MAT_io_pipe_phv_out_data_160; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_161 = MAT_io_pipe_phv_out_data_161; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_162 = MAT_io_pipe_phv_out_data_162; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_163 = MAT_io_pipe_phv_out_data_163; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_164 = MAT_io_pipe_phv_out_data_164; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_165 = MAT_io_pipe_phv_out_data_165; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_166 = MAT_io_pipe_phv_out_data_166; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_167 = MAT_io_pipe_phv_out_data_167; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_168 = MAT_io_pipe_phv_out_data_168; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_169 = MAT_io_pipe_phv_out_data_169; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_170 = MAT_io_pipe_phv_out_data_170; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_171 = MAT_io_pipe_phv_out_data_171; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_172 = MAT_io_pipe_phv_out_data_172; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_173 = MAT_io_pipe_phv_out_data_173; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_174 = MAT_io_pipe_phv_out_data_174; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_175 = MAT_io_pipe_phv_out_data_175; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_176 = MAT_io_pipe_phv_out_data_176; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_177 = MAT_io_pipe_phv_out_data_177; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_178 = MAT_io_pipe_phv_out_data_178; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_179 = MAT_io_pipe_phv_out_data_179; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_180 = MAT_io_pipe_phv_out_data_180; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_181 = MAT_io_pipe_phv_out_data_181; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_182 = MAT_io_pipe_phv_out_data_182; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_183 = MAT_io_pipe_phv_out_data_183; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_184 = MAT_io_pipe_phv_out_data_184; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_185 = MAT_io_pipe_phv_out_data_185; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_186 = MAT_io_pipe_phv_out_data_186; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_187 = MAT_io_pipe_phv_out_data_187; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_188 = MAT_io_pipe_phv_out_data_188; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_189 = MAT_io_pipe_phv_out_data_189; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_190 = MAT_io_pipe_phv_out_data_190; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_191 = MAT_io_pipe_phv_out_data_191; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_192 = MAT_io_pipe_phv_out_data_192; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_193 = MAT_io_pipe_phv_out_data_193; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_194 = MAT_io_pipe_phv_out_data_194; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_195 = MAT_io_pipe_phv_out_data_195; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_196 = MAT_io_pipe_phv_out_data_196; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_197 = MAT_io_pipe_phv_out_data_197; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_198 = MAT_io_pipe_phv_out_data_198; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_199 = MAT_io_pipe_phv_out_data_199; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_200 = MAT_io_pipe_phv_out_data_200; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_201 = MAT_io_pipe_phv_out_data_201; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_202 = MAT_io_pipe_phv_out_data_202; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_203 = MAT_io_pipe_phv_out_data_203; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_204 = MAT_io_pipe_phv_out_data_204; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_205 = MAT_io_pipe_phv_out_data_205; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_206 = MAT_io_pipe_phv_out_data_206; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_207 = MAT_io_pipe_phv_out_data_207; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_208 = MAT_io_pipe_phv_out_data_208; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_209 = MAT_io_pipe_phv_out_data_209; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_210 = MAT_io_pipe_phv_out_data_210; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_211 = MAT_io_pipe_phv_out_data_211; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_212 = MAT_io_pipe_phv_out_data_212; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_213 = MAT_io_pipe_phv_out_data_213; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_214 = MAT_io_pipe_phv_out_data_214; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_215 = MAT_io_pipe_phv_out_data_215; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_216 = MAT_io_pipe_phv_out_data_216; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_217 = MAT_io_pipe_phv_out_data_217; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_218 = MAT_io_pipe_phv_out_data_218; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_219 = MAT_io_pipe_phv_out_data_219; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_220 = MAT_io_pipe_phv_out_data_220; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_221 = MAT_io_pipe_phv_out_data_221; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_222 = MAT_io_pipe_phv_out_data_222; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_223 = MAT_io_pipe_phv_out_data_223; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_224 = MAT_io_pipe_phv_out_data_224; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_225 = MAT_io_pipe_phv_out_data_225; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_226 = MAT_io_pipe_phv_out_data_226; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_227 = MAT_io_pipe_phv_out_data_227; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_228 = MAT_io_pipe_phv_out_data_228; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_229 = MAT_io_pipe_phv_out_data_229; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_230 = MAT_io_pipe_phv_out_data_230; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_231 = MAT_io_pipe_phv_out_data_231; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_232 = MAT_io_pipe_phv_out_data_232; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_233 = MAT_io_pipe_phv_out_data_233; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_234 = MAT_io_pipe_phv_out_data_234; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_235 = MAT_io_pipe_phv_out_data_235; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_236 = MAT_io_pipe_phv_out_data_236; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_237 = MAT_io_pipe_phv_out_data_237; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_238 = MAT_io_pipe_phv_out_data_238; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_239 = MAT_io_pipe_phv_out_data_239; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_240 = MAT_io_pipe_phv_out_data_240; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_241 = MAT_io_pipe_phv_out_data_241; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_242 = MAT_io_pipe_phv_out_data_242; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_243 = MAT_io_pipe_phv_out_data_243; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_244 = MAT_io_pipe_phv_out_data_244; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_245 = MAT_io_pipe_phv_out_data_245; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_246 = MAT_io_pipe_phv_out_data_246; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_247 = MAT_io_pipe_phv_out_data_247; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_248 = MAT_io_pipe_phv_out_data_248; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_249 = MAT_io_pipe_phv_out_data_249; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_250 = MAT_io_pipe_phv_out_data_250; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_251 = MAT_io_pipe_phv_out_data_251; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_252 = MAT_io_pipe_phv_out_data_252; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_253 = MAT_io_pipe_phv_out_data_253; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_254 = MAT_io_pipe_phv_out_data_254; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_255 = MAT_io_pipe_phv_out_data_255; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_256 = MAT_io_pipe_phv_out_data_256; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_257 = MAT_io_pipe_phv_out_data_257; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_258 = MAT_io_pipe_phv_out_data_258; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_259 = MAT_io_pipe_phv_out_data_259; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_260 = MAT_io_pipe_phv_out_data_260; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_261 = MAT_io_pipe_phv_out_data_261; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_262 = MAT_io_pipe_phv_out_data_262; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_263 = MAT_io_pipe_phv_out_data_263; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_264 = MAT_io_pipe_phv_out_data_264; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_265 = MAT_io_pipe_phv_out_data_265; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_266 = MAT_io_pipe_phv_out_data_266; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_267 = MAT_io_pipe_phv_out_data_267; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_268 = MAT_io_pipe_phv_out_data_268; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_269 = MAT_io_pipe_phv_out_data_269; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_270 = MAT_io_pipe_phv_out_data_270; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_271 = MAT_io_pipe_phv_out_data_271; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_272 = MAT_io_pipe_phv_out_data_272; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_273 = MAT_io_pipe_phv_out_data_273; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_274 = MAT_io_pipe_phv_out_data_274; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_275 = MAT_io_pipe_phv_out_data_275; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_276 = MAT_io_pipe_phv_out_data_276; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_277 = MAT_io_pipe_phv_out_data_277; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_278 = MAT_io_pipe_phv_out_data_278; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_279 = MAT_io_pipe_phv_out_data_279; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_280 = MAT_io_pipe_phv_out_data_280; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_281 = MAT_io_pipe_phv_out_data_281; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_282 = MAT_io_pipe_phv_out_data_282; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_283 = MAT_io_pipe_phv_out_data_283; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_284 = MAT_io_pipe_phv_out_data_284; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_285 = MAT_io_pipe_phv_out_data_285; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_286 = MAT_io_pipe_phv_out_data_286; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_287 = MAT_io_pipe_phv_out_data_287; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_288 = MAT_io_pipe_phv_out_data_288; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_289 = MAT_io_pipe_phv_out_data_289; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_290 = MAT_io_pipe_phv_out_data_290; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_291 = MAT_io_pipe_phv_out_data_291; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_292 = MAT_io_pipe_phv_out_data_292; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_293 = MAT_io_pipe_phv_out_data_293; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_294 = MAT_io_pipe_phv_out_data_294; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_295 = MAT_io_pipe_phv_out_data_295; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_296 = MAT_io_pipe_phv_out_data_296; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_297 = MAT_io_pipe_phv_out_data_297; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_298 = MAT_io_pipe_phv_out_data_298; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_299 = MAT_io_pipe_phv_out_data_299; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_300 = MAT_io_pipe_phv_out_data_300; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_301 = MAT_io_pipe_phv_out_data_301; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_302 = MAT_io_pipe_phv_out_data_302; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_303 = MAT_io_pipe_phv_out_data_303; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_304 = MAT_io_pipe_phv_out_data_304; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_305 = MAT_io_pipe_phv_out_data_305; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_306 = MAT_io_pipe_phv_out_data_306; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_307 = MAT_io_pipe_phv_out_data_307; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_308 = MAT_io_pipe_phv_out_data_308; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_309 = MAT_io_pipe_phv_out_data_309; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_310 = MAT_io_pipe_phv_out_data_310; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_311 = MAT_io_pipe_phv_out_data_311; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_312 = MAT_io_pipe_phv_out_data_312; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_313 = MAT_io_pipe_phv_out_data_313; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_314 = MAT_io_pipe_phv_out_data_314; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_315 = MAT_io_pipe_phv_out_data_315; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_316 = MAT_io_pipe_phv_out_data_316; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_317 = MAT_io_pipe_phv_out_data_317; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_318 = MAT_io_pipe_phv_out_data_318; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_319 = MAT_io_pipe_phv_out_data_319; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_320 = MAT_io_pipe_phv_out_data_320; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_321 = MAT_io_pipe_phv_out_data_321; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_322 = MAT_io_pipe_phv_out_data_322; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_323 = MAT_io_pipe_phv_out_data_323; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_324 = MAT_io_pipe_phv_out_data_324; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_325 = MAT_io_pipe_phv_out_data_325; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_326 = MAT_io_pipe_phv_out_data_326; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_327 = MAT_io_pipe_phv_out_data_327; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_328 = MAT_io_pipe_phv_out_data_328; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_329 = MAT_io_pipe_phv_out_data_329; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_330 = MAT_io_pipe_phv_out_data_330; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_331 = MAT_io_pipe_phv_out_data_331; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_332 = MAT_io_pipe_phv_out_data_332; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_333 = MAT_io_pipe_phv_out_data_333; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_334 = MAT_io_pipe_phv_out_data_334; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_335 = MAT_io_pipe_phv_out_data_335; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_336 = MAT_io_pipe_phv_out_data_336; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_337 = MAT_io_pipe_phv_out_data_337; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_338 = MAT_io_pipe_phv_out_data_338; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_339 = MAT_io_pipe_phv_out_data_339; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_340 = MAT_io_pipe_phv_out_data_340; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_341 = MAT_io_pipe_phv_out_data_341; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_342 = MAT_io_pipe_phv_out_data_342; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_343 = MAT_io_pipe_phv_out_data_343; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_344 = MAT_io_pipe_phv_out_data_344; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_345 = MAT_io_pipe_phv_out_data_345; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_346 = MAT_io_pipe_phv_out_data_346; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_347 = MAT_io_pipe_phv_out_data_347; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_348 = MAT_io_pipe_phv_out_data_348; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_349 = MAT_io_pipe_phv_out_data_349; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_350 = MAT_io_pipe_phv_out_data_350; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_351 = MAT_io_pipe_phv_out_data_351; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_352 = MAT_io_pipe_phv_out_data_352; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_353 = MAT_io_pipe_phv_out_data_353; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_354 = MAT_io_pipe_phv_out_data_354; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_355 = MAT_io_pipe_phv_out_data_355; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_356 = MAT_io_pipe_phv_out_data_356; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_357 = MAT_io_pipe_phv_out_data_357; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_358 = MAT_io_pipe_phv_out_data_358; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_359 = MAT_io_pipe_phv_out_data_359; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_360 = MAT_io_pipe_phv_out_data_360; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_361 = MAT_io_pipe_phv_out_data_361; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_362 = MAT_io_pipe_phv_out_data_362; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_363 = MAT_io_pipe_phv_out_data_363; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_364 = MAT_io_pipe_phv_out_data_364; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_365 = MAT_io_pipe_phv_out_data_365; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_366 = MAT_io_pipe_phv_out_data_366; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_367 = MAT_io_pipe_phv_out_data_367; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_368 = MAT_io_pipe_phv_out_data_368; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_369 = MAT_io_pipe_phv_out_data_369; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_370 = MAT_io_pipe_phv_out_data_370; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_371 = MAT_io_pipe_phv_out_data_371; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_372 = MAT_io_pipe_phv_out_data_372; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_373 = MAT_io_pipe_phv_out_data_373; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_374 = MAT_io_pipe_phv_out_data_374; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_375 = MAT_io_pipe_phv_out_data_375; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_376 = MAT_io_pipe_phv_out_data_376; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_377 = MAT_io_pipe_phv_out_data_377; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_378 = MAT_io_pipe_phv_out_data_378; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_379 = MAT_io_pipe_phv_out_data_379; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_380 = MAT_io_pipe_phv_out_data_380; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_381 = MAT_io_pipe_phv_out_data_381; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_382 = MAT_io_pipe_phv_out_data_382; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_383 = MAT_io_pipe_phv_out_data_383; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_384 = MAT_io_pipe_phv_out_data_384; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_385 = MAT_io_pipe_phv_out_data_385; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_386 = MAT_io_pipe_phv_out_data_386; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_387 = MAT_io_pipe_phv_out_data_387; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_388 = MAT_io_pipe_phv_out_data_388; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_389 = MAT_io_pipe_phv_out_data_389; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_390 = MAT_io_pipe_phv_out_data_390; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_391 = MAT_io_pipe_phv_out_data_391; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_392 = MAT_io_pipe_phv_out_data_392; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_393 = MAT_io_pipe_phv_out_data_393; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_394 = MAT_io_pipe_phv_out_data_394; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_395 = MAT_io_pipe_phv_out_data_395; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_396 = MAT_io_pipe_phv_out_data_396; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_397 = MAT_io_pipe_phv_out_data_397; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_398 = MAT_io_pipe_phv_out_data_398; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_399 = MAT_io_pipe_phv_out_data_399; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_400 = MAT_io_pipe_phv_out_data_400; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_401 = MAT_io_pipe_phv_out_data_401; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_402 = MAT_io_pipe_phv_out_data_402; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_403 = MAT_io_pipe_phv_out_data_403; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_404 = MAT_io_pipe_phv_out_data_404; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_405 = MAT_io_pipe_phv_out_data_405; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_406 = MAT_io_pipe_phv_out_data_406; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_407 = MAT_io_pipe_phv_out_data_407; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_408 = MAT_io_pipe_phv_out_data_408; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_409 = MAT_io_pipe_phv_out_data_409; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_410 = MAT_io_pipe_phv_out_data_410; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_411 = MAT_io_pipe_phv_out_data_411; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_412 = MAT_io_pipe_phv_out_data_412; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_413 = MAT_io_pipe_phv_out_data_413; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_414 = MAT_io_pipe_phv_out_data_414; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_415 = MAT_io_pipe_phv_out_data_415; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_416 = MAT_io_pipe_phv_out_data_416; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_417 = MAT_io_pipe_phv_out_data_417; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_418 = MAT_io_pipe_phv_out_data_418; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_419 = MAT_io_pipe_phv_out_data_419; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_420 = MAT_io_pipe_phv_out_data_420; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_421 = MAT_io_pipe_phv_out_data_421; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_422 = MAT_io_pipe_phv_out_data_422; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_423 = MAT_io_pipe_phv_out_data_423; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_424 = MAT_io_pipe_phv_out_data_424; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_425 = MAT_io_pipe_phv_out_data_425; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_426 = MAT_io_pipe_phv_out_data_426; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_427 = MAT_io_pipe_phv_out_data_427; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_428 = MAT_io_pipe_phv_out_data_428; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_429 = MAT_io_pipe_phv_out_data_429; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_430 = MAT_io_pipe_phv_out_data_430; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_431 = MAT_io_pipe_phv_out_data_431; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_432 = MAT_io_pipe_phv_out_data_432; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_433 = MAT_io_pipe_phv_out_data_433; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_434 = MAT_io_pipe_phv_out_data_434; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_435 = MAT_io_pipe_phv_out_data_435; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_436 = MAT_io_pipe_phv_out_data_436; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_437 = MAT_io_pipe_phv_out_data_437; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_438 = MAT_io_pipe_phv_out_data_438; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_439 = MAT_io_pipe_phv_out_data_439; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_440 = MAT_io_pipe_phv_out_data_440; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_441 = MAT_io_pipe_phv_out_data_441; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_442 = MAT_io_pipe_phv_out_data_442; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_443 = MAT_io_pipe_phv_out_data_443; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_444 = MAT_io_pipe_phv_out_data_444; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_445 = MAT_io_pipe_phv_out_data_445; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_446 = MAT_io_pipe_phv_out_data_446; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_447 = MAT_io_pipe_phv_out_data_447; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_448 = MAT_io_pipe_phv_out_data_448; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_449 = MAT_io_pipe_phv_out_data_449; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_450 = MAT_io_pipe_phv_out_data_450; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_451 = MAT_io_pipe_phv_out_data_451; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_452 = MAT_io_pipe_phv_out_data_452; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_453 = MAT_io_pipe_phv_out_data_453; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_454 = MAT_io_pipe_phv_out_data_454; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_455 = MAT_io_pipe_phv_out_data_455; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_456 = MAT_io_pipe_phv_out_data_456; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_457 = MAT_io_pipe_phv_out_data_457; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_458 = MAT_io_pipe_phv_out_data_458; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_459 = MAT_io_pipe_phv_out_data_459; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_460 = MAT_io_pipe_phv_out_data_460; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_461 = MAT_io_pipe_phv_out_data_461; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_462 = MAT_io_pipe_phv_out_data_462; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_463 = MAT_io_pipe_phv_out_data_463; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_464 = MAT_io_pipe_phv_out_data_464; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_465 = MAT_io_pipe_phv_out_data_465; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_466 = MAT_io_pipe_phv_out_data_466; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_467 = MAT_io_pipe_phv_out_data_467; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_468 = MAT_io_pipe_phv_out_data_468; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_469 = MAT_io_pipe_phv_out_data_469; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_470 = MAT_io_pipe_phv_out_data_470; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_471 = MAT_io_pipe_phv_out_data_471; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_472 = MAT_io_pipe_phv_out_data_472; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_473 = MAT_io_pipe_phv_out_data_473; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_474 = MAT_io_pipe_phv_out_data_474; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_475 = MAT_io_pipe_phv_out_data_475; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_476 = MAT_io_pipe_phv_out_data_476; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_477 = MAT_io_pipe_phv_out_data_477; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_478 = MAT_io_pipe_phv_out_data_478; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_479 = MAT_io_pipe_phv_out_data_479; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_480 = MAT_io_pipe_phv_out_data_480; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_481 = MAT_io_pipe_phv_out_data_481; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_482 = MAT_io_pipe_phv_out_data_482; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_483 = MAT_io_pipe_phv_out_data_483; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_484 = MAT_io_pipe_phv_out_data_484; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_485 = MAT_io_pipe_phv_out_data_485; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_486 = MAT_io_pipe_phv_out_data_486; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_487 = MAT_io_pipe_phv_out_data_487; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_488 = MAT_io_pipe_phv_out_data_488; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_489 = MAT_io_pipe_phv_out_data_489; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_490 = MAT_io_pipe_phv_out_data_490; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_491 = MAT_io_pipe_phv_out_data_491; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_492 = MAT_io_pipe_phv_out_data_492; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_493 = MAT_io_pipe_phv_out_data_493; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_494 = MAT_io_pipe_phv_out_data_494; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_495 = MAT_io_pipe_phv_out_data_495; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_496 = MAT_io_pipe_phv_out_data_496; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_497 = MAT_io_pipe_phv_out_data_497; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_498 = MAT_io_pipe_phv_out_data_498; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_499 = MAT_io_pipe_phv_out_data_499; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_500 = MAT_io_pipe_phv_out_data_500; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_501 = MAT_io_pipe_phv_out_data_501; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_502 = MAT_io_pipe_phv_out_data_502; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_503 = MAT_io_pipe_phv_out_data_503; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_504 = MAT_io_pipe_phv_out_data_504; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_505 = MAT_io_pipe_phv_out_data_505; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_506 = MAT_io_pipe_phv_out_data_506; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_507 = MAT_io_pipe_phv_out_data_507; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_508 = MAT_io_pipe_phv_out_data_508; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_509 = MAT_io_pipe_phv_out_data_509; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_510 = MAT_io_pipe_phv_out_data_510; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_511 = MAT_io_pipe_phv_out_data_511; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_0 = MAT_io_pipe_phv_out_header_0; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_1 = MAT_io_pipe_phv_out_header_1; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_2 = MAT_io_pipe_phv_out_header_2; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_3 = MAT_io_pipe_phv_out_header_3; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_4 = MAT_io_pipe_phv_out_header_4; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_5 = MAT_io_pipe_phv_out_header_5; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_6 = MAT_io_pipe_phv_out_header_6; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_7 = MAT_io_pipe_phv_out_header_7; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_8 = MAT_io_pipe_phv_out_header_8; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_9 = MAT_io_pipe_phv_out_header_9; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_10 = MAT_io_pipe_phv_out_header_10; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_11 = MAT_io_pipe_phv_out_header_11; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_12 = MAT_io_pipe_phv_out_header_12; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_13 = MAT_io_pipe_phv_out_header_13; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_14 = MAT_io_pipe_phv_out_header_14; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_15 = MAT_io_pipe_phv_out_header_15; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_parse_current_state = MAT_io_pipe_phv_out_parse_current_state; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_parse_current_offset = MAT_io_pipe_phv_out_parse_current_offset; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_parse_transition_field = MAT_io_pipe_phv_out_parse_transition_field; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_next_processor_id = MAT_io_pipe_phv_out_next_processor_id; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_next_config_id = MAT_io_pipe_phv_out_next_config_id; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_is_valid_processor = MAT_io_pipe_phv_out_is_valid_processor; // @[processor.scala 24:24]
  assign EXE_io_hit = MAT_io_hit; // @[processor.scala 25:24]
  assign EXE_io_match_value = MAT_io_match_value; // @[processor.scala 26:24]
  assign EXE_io_action_mod_en_0 = io_mod_act_mod_en_0; // @[processor.scala 27:24]
  assign EXE_io_action_mod_en_1 = io_mod_act_mod_en_1; // @[processor.scala 27:24]
  assign EXE_io_action_mod_addr = io_mod_act_mod_addr; // @[processor.scala 27:24]
  assign EXE_io_action_mod_data_0 = io_mod_act_mod_data_0; // @[processor.scala 27:24]
  assign EXE_io_action_mod_data_1 = io_mod_act_mod_data_1; // @[processor.scala 27:24]
endmodule
