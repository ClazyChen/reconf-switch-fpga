module Matcher(
  input         clock,
  input         reset,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input         io_mod_en,
  input         io_mod_config_id,
  input  [7:0]  io_mod_key_mod_header_id,
  input  [7:0]  io_mod_key_mod_internal_offset,
  input  [3:0]  io_mod_key_mod_key_length,
  input  [3:0]  io_mod_key_mod_val_length,
  input  [2:0]  io_mod_table_mod_sram_id_table_0,
  input  [2:0]  io_mod_table_mod_sram_id_table_1,
  input  [2:0]  io_mod_table_mod_sram_id_table_2,
  input  [2:0]  io_mod_table_mod_sram_id_table_3,
  input  [2:0]  io_mod_table_mod_sram_id_table_4,
  input  [2:0]  io_mod_table_mod_sram_id_table_5,
  input  [2:0]  io_mod_table_mod_sram_id_table_6,
  input  [2:0]  io_mod_table_mod_sram_id_table_7,
  input  [3:0]  io_mod_table_mod_table_width,
  input  [3:0]  io_mod_table_mod_table_depth,
  output        io_hit,
  output [63:0] io_match_value,
  output        io_mem_cluster_0_en,
  output [7:0]  io_mem_cluster_0_addr,
  input  [63:0] io_mem_cluster_0_data,
  output        io_mem_cluster_1_en,
  output [7:0]  io_mem_cluster_1_addr,
  input  [63:0] io_mem_cluster_1_data,
  output        io_mem_cluster_2_en,
  output [7:0]  io_mem_cluster_2_addr,
  input  [63:0] io_mem_cluster_2_data,
  output        io_mem_cluster_3_en,
  output [7:0]  io_mem_cluster_3_addr,
  input  [63:0] io_mem_cluster_3_data,
  output        io_mem_cluster_4_en,
  output [7:0]  io_mem_cluster_4_addr,
  input  [63:0] io_mem_cluster_4_data,
  output        io_mem_cluster_5_en,
  output [7:0]  io_mem_cluster_5_addr,
  input  [63:0] io_mem_cluster_5_data,
  output        io_mem_cluster_6_en,
  output [7:0]  io_mem_cluster_6_addr,
  input  [63:0] io_mem_cluster_6_data,
  output        io_mem_cluster_7_en,
  output [7:0]  io_mem_cluster_7_addr,
  input  [63:0] io_mem_cluster_7_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  pipe1_clock; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_0; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_1; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_2; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_3; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_4; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_5; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_6; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_7; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_8; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_9; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_10; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_11; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_12; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_13; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_14; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_15; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_16; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_17; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_18; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_19; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_20; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_21; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_22; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_23; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_24; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_25; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_26; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_27; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_28; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_29; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_30; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_31; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_32; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_33; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_34; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_35; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_36; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_37; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_38; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_39; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_40; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_41; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_42; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_43; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_44; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_45; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_46; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_47; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_48; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_49; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_50; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_51; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_52; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_53; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_54; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_55; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_56; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_57; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_58; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_59; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_60; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_61; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_62; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_63; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_64; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_65; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_66; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_67; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_68; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_69; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_70; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_71; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_72; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_73; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_74; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_75; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_76; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_77; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_78; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_79; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_80; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_81; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_82; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_83; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_84; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_85; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_86; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_87; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_88; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_89; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_90; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_91; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_92; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_93; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_94; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_95; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_0; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_1; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_2; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_3; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_4; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_5; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_6; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_7; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_8; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_9; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_10; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_11; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_12; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_13; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_14; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_15; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_state; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 264:23]
  wire [1:0] pipe1_io_pipe_phv_in_next_processor_id; // @[matcher.scala 264:23]
  wire  pipe1_io_pipe_phv_in_next_config_id; // @[matcher.scala 264:23]
  wire  pipe1_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_0; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_1; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_2; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_3; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_4; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_5; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_6; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_7; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_8; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_9; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_10; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_11; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_12; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_13; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_14; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_15; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_16; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_17; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_18; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_19; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_20; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_21; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_22; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_23; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_24; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_25; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_26; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_27; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_28; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_29; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_30; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_31; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_32; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_33; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_34; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_35; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_36; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_37; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_38; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_39; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_40; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_41; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_42; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_43; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_44; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_45; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_46; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_47; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_48; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_49; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_50; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_51; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_52; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_53; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_54; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_55; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_56; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_57; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_58; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_59; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_60; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_61; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_62; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_63; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_64; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_65; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_66; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_67; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_68; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_69; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_70; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_71; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_72; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_73; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_74; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_75; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_76; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_77; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_78; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_79; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_80; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_81; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_82; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_83; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_84; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_85; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_86; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_87; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_88; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_89; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_90; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_91; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_92; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_93; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_94; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_95; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_0; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_1; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_2; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_3; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_4; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_5; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_6; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_7; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_8; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_9; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_10; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_11; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_12; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_13; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_14; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_15; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_state; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 264:23]
  wire [15:0] pipe1_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 264:23]
  wire [1:0] pipe1_io_pipe_phv_out_next_processor_id; // @[matcher.scala 264:23]
  wire  pipe1_io_pipe_phv_out_next_config_id; // @[matcher.scala 264:23]
  wire  pipe1_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_key_config_0_header_id; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_key_config_0_internal_offset; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_key_config_1_header_id; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_key_config_1_internal_offset; // @[matcher.scala 264:23]
  wire [7:0] pipe1_io_key_offset; // @[matcher.scala 264:23]
  wire  pipe2_clock; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_0; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_1; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_2; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_3; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_4; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_5; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_6; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_7; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_8; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_9; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_10; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_11; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_12; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_13; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_14; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_15; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_16; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_17; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_18; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_19; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_20; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_21; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_22; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_23; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_24; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_25; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_26; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_27; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_28; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_29; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_30; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_31; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_32; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_33; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_34; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_35; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_36; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_37; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_38; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_39; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_40; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_41; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_42; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_43; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_44; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_45; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_46; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_47; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_48; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_49; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_50; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_51; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_52; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_53; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_54; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_55; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_56; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_57; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_58; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_59; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_60; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_61; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_62; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_63; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_64; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_65; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_66; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_67; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_68; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_69; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_70; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_71; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_72; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_73; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_74; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_75; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_76; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_77; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_78; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_79; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_80; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_81; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_82; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_83; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_84; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_85; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_86; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_87; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_88; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_89; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_90; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_91; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_92; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_93; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_94; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_95; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_0; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_1; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_2; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_3; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_4; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_5; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_6; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_7; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_8; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_9; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_10; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_11; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_12; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_13; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_14; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_15; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_state; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 265:23]
  wire [1:0] pipe2_io_pipe_phv_in_next_processor_id; // @[matcher.scala 265:23]
  wire  pipe2_io_pipe_phv_in_next_config_id; // @[matcher.scala 265:23]
  wire  pipe2_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_0; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_1; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_2; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_3; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_4; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_5; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_6; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_7; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_8; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_9; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_10; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_11; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_12; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_13; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_14; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_15; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_16; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_17; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_18; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_19; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_20; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_21; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_22; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_23; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_24; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_25; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_26; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_27; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_28; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_29; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_30; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_31; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_32; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_33; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_34; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_35; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_36; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_37; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_38; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_39; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_40; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_41; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_42; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_43; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_44; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_45; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_46; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_47; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_48; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_49; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_50; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_51; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_52; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_53; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_54; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_55; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_56; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_57; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_58; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_59; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_60; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_61; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_62; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_63; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_64; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_65; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_66; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_67; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_68; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_69; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_70; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_71; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_72; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_73; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_74; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_75; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_76; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_77; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_78; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_79; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_80; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_81; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_82; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_83; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_84; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_85; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_86; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_87; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_88; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_89; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_90; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_91; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_92; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_93; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_94; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_95; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_0; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_1; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_2; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_3; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_4; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_5; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_6; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_7; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_8; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_9; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_10; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_11; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_12; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_13; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_14; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_15; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_state; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 265:23]
  wire [15:0] pipe2_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 265:23]
  wire [1:0] pipe2_io_pipe_phv_out_next_processor_id; // @[matcher.scala 265:23]
  wire  pipe2_io_pipe_phv_out_next_config_id; // @[matcher.scala 265:23]
  wire  pipe2_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 265:23]
  wire [3:0] pipe2_io_key_config_0_key_length; // @[matcher.scala 265:23]
  wire [3:0] pipe2_io_key_config_1_key_length; // @[matcher.scala 265:23]
  wire [7:0] pipe2_io_key_offset; // @[matcher.scala 265:23]
  wire [63:0] pipe2_io_match_key; // @[matcher.scala 265:23]
  wire  pipe3to8_clock; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_0; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_1; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_2; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_3; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_4; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_5; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_6; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_7; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_8; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_9; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_10; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_11; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_12; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_13; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_14; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_15; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_16; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_17; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_18; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_19; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_20; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_21; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_22; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_23; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_24; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_25; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_26; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_27; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_28; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_29; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_30; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_31; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_32; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_33; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_34; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_35; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_36; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_37; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_38; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_39; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_40; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_41; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_42; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_43; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_44; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_45; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_46; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_47; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_48; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_49; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_50; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_51; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_52; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_53; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_54; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_55; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_56; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_57; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_58; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_59; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_60; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_61; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_62; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_63; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_64; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_65; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_66; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_67; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_68; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_69; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_70; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_71; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_72; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_73; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_74; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_75; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_76; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_77; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_78; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_79; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_80; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_81; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_82; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_83; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_84; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_85; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_86; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_87; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_88; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_89; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_90; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_91; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_92; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_93; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_94; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_95; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_0; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_1; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_2; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_3; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_4; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_5; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_6; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_7; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_8; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_9; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_10; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_11; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_12; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_13; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_14; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_15; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_parse_current_state; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 266:26]
  wire [1:0] pipe3to8_io_pipe_phv_in_next_processor_id; // @[matcher.scala 266:26]
  wire  pipe3to8_io_pipe_phv_in_next_config_id; // @[matcher.scala 266:26]
  wire  pipe3to8_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_0; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_1; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_2; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_3; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_4; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_5; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_6; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_7; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_8; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_9; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_10; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_11; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_12; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_13; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_14; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_15; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_16; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_17; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_18; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_19; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_20; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_21; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_22; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_23; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_24; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_25; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_26; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_27; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_28; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_29; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_30; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_31; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_32; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_33; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_34; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_35; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_36; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_37; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_38; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_39; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_40; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_41; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_42; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_43; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_44; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_45; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_46; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_47; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_48; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_49; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_50; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_51; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_52; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_53; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_54; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_55; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_56; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_57; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_58; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_59; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_60; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_61; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_62; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_63; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_64; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_65; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_66; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_67; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_68; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_69; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_70; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_71; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_72; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_73; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_74; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_75; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_76; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_77; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_78; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_79; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_80; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_81; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_82; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_83; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_84; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_85; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_86; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_87; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_88; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_89; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_90; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_91; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_92; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_93; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_94; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_95; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_0; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_1; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_2; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_3; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_4; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_5; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_6; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_7; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_8; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_9; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_10; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_11; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_12; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_13; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_14; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_15; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_parse_current_state; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 266:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 266:26]
  wire [1:0] pipe3to8_io_pipe_phv_out_next_processor_id; // @[matcher.scala 266:26]
  wire  pipe3to8_io_pipe_phv_out_next_config_id; // @[matcher.scala 266:26]
  wire  pipe3to8_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 266:26]
  wire  pipe3to8_io_mod_hash_depth_mod; // @[matcher.scala 266:26]
  wire  pipe3to8_io_mod_config_id; // @[matcher.scala 266:26]
  wire [2:0] pipe3to8_io_mod_hash_depth; // @[matcher.scala 266:26]
  wire [63:0] pipe3to8_io_key_in; // @[matcher.scala 266:26]
  wire [63:0] pipe3to8_io_key_out; // @[matcher.scala 266:26]
  wire [7:0] pipe3to8_io_hash_val; // @[matcher.scala 266:26]
  wire [2:0] pipe3to8_io_hash_val_cs; // @[matcher.scala 266:26]
  wire  pipe9_clock; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_0; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_1; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_2; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_3; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_4; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_5; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_6; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_7; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_8; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_9; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_10; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_11; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_12; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_13; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_14; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_15; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_16; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_17; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_18; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_19; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_20; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_21; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_22; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_23; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_24; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_25; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_26; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_27; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_28; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_29; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_30; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_31; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_32; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_33; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_34; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_35; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_36; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_37; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_38; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_39; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_40; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_41; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_42; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_43; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_44; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_45; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_46; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_47; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_48; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_49; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_50; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_51; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_52; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_53; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_54; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_55; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_56; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_57; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_58; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_59; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_60; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_61; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_62; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_63; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_64; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_65; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_66; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_67; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_68; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_69; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_70; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_71; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_72; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_73; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_74; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_75; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_76; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_77; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_78; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_79; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_80; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_81; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_82; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_83; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_84; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_85; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_86; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_87; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_88; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_89; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_90; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_91; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_92; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_93; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_94; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_95; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_0; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_1; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_2; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_3; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_4; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_5; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_6; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_7; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_8; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_9; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_10; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_11; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_12; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_13; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_14; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_15; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_parse_current_state; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 267:23]
  wire [1:0] pipe9_io_pipe_phv_in_next_processor_id; // @[matcher.scala 267:23]
  wire  pipe9_io_pipe_phv_in_next_config_id; // @[matcher.scala 267:23]
  wire  pipe9_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_0; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_1; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_2; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_3; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_4; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_5; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_6; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_7; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_8; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_9; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_10; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_11; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_12; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_13; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_14; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_15; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_16; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_17; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_18; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_19; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_20; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_21; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_22; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_23; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_24; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_25; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_26; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_27; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_28; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_29; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_30; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_31; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_32; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_33; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_34; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_35; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_36; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_37; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_38; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_39; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_40; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_41; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_42; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_43; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_44; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_45; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_46; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_47; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_48; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_49; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_50; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_51; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_52; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_53; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_54; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_55; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_56; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_57; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_58; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_59; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_60; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_61; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_62; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_63; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_64; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_65; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_66; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_67; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_68; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_69; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_70; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_71; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_72; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_73; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_74; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_75; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_76; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_77; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_78; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_79; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_80; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_81; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_82; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_83; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_84; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_85; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_86; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_87; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_88; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_89; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_90; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_91; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_92; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_93; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_94; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_95; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_0; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_1; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_2; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_3; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_4; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_5; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_6; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_7; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_8; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_9; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_10; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_11; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_12; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_13; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_14; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_15; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_parse_current_state; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 267:23]
  wire [15:0] pipe9_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 267:23]
  wire [1:0] pipe9_io_pipe_phv_out_next_processor_id; // @[matcher.scala 267:23]
  wire  pipe9_io_pipe_phv_out_next_config_id; // @[matcher.scala 267:23]
  wire  pipe9_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 267:23]
  wire [3:0] pipe9_io_table_config_0_table_width; // @[matcher.scala 267:23]
  wire [3:0] pipe9_io_table_config_0_table_depth; // @[matcher.scala 267:23]
  wire [3:0] pipe9_io_table_config_1_table_width; // @[matcher.scala 267:23]
  wire [3:0] pipe9_io_table_config_1_table_depth; // @[matcher.scala 267:23]
  wire [63:0] pipe9_io_key_in; // @[matcher.scala 267:23]
  wire [63:0] pipe9_io_key_out; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_addr_in; // @[matcher.scala 267:23]
  wire [7:0] pipe9_io_addr_out; // @[matcher.scala 267:23]
  wire [2:0] pipe9_io_cs_in; // @[matcher.scala 267:23]
  wire [2:0] pipe9_io_cs_out; // @[matcher.scala 267:23]
  wire  pipe9_io_cs_vec_out_0; // @[matcher.scala 267:23]
  wire  pipe9_io_cs_vec_out_1; // @[matcher.scala 267:23]
  wire  pipe9_io_cs_vec_out_2; // @[matcher.scala 267:23]
  wire  pipe9_io_cs_vec_out_3; // @[matcher.scala 267:23]
  wire  pipe9_io_cs_vec_out_4; // @[matcher.scala 267:23]
  wire  pipe9_io_cs_vec_out_5; // @[matcher.scala 267:23]
  wire  pipe9_io_cs_vec_out_6; // @[matcher.scala 267:23]
  wire  pipe9_io_cs_vec_out_7; // @[matcher.scala 267:23]
  wire  pipe10_clock; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_0; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_1; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_2; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_3; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_4; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_5; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_6; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_7; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_8; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_9; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_10; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_11; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_12; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_13; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_14; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_15; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_16; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_17; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_18; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_19; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_20; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_21; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_22; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_23; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_24; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_25; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_26; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_27; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_28; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_29; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_30; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_31; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_32; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_33; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_34; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_35; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_36; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_37; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_38; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_39; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_40; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_41; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_42; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_43; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_44; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_45; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_46; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_47; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_48; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_49; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_50; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_51; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_52; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_53; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_54; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_55; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_56; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_57; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_58; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_59; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_60; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_61; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_62; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_63; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_64; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_65; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_66; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_67; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_68; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_69; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_70; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_71; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_72; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_73; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_74; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_75; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_76; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_77; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_78; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_79; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_80; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_81; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_82; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_83; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_84; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_85; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_86; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_87; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_88; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_89; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_90; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_91; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_92; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_93; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_94; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_95; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_0; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_1; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_2; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_3; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_4; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_5; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_6; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_7; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_8; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_9; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_10; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_11; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_12; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_13; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_14; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_15; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_parse_current_state; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 268:24]
  wire [1:0] pipe10_io_pipe_phv_in_next_processor_id; // @[matcher.scala 268:24]
  wire  pipe10_io_pipe_phv_in_next_config_id; // @[matcher.scala 268:24]
  wire  pipe10_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_0; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_1; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_2; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_3; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_4; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_5; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_6; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_7; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_8; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_9; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_10; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_11; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_12; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_13; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_14; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_15; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_16; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_17; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_18; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_19; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_20; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_21; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_22; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_23; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_24; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_25; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_26; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_27; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_28; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_29; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_30; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_31; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_32; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_33; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_34; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_35; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_36; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_37; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_38; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_39; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_40; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_41; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_42; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_43; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_44; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_45; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_46; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_47; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_48; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_49; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_50; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_51; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_52; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_53; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_54; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_55; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_56; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_57; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_58; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_59; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_60; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_61; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_62; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_63; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_64; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_65; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_66; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_67; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_68; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_69; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_70; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_71; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_72; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_73; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_74; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_75; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_76; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_77; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_78; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_79; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_80; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_81; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_82; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_83; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_84; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_85; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_86; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_87; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_88; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_89; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_90; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_91; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_92; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_93; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_94; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_95; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_0; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_1; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_2; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_3; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_4; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_5; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_6; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_7; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_8; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_9; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_10; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_11; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_12; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_13; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_14; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_15; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_parse_current_state; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 268:24]
  wire [15:0] pipe10_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 268:24]
  wire [1:0] pipe10_io_pipe_phv_out_next_processor_id; // @[matcher.scala 268:24]
  wire  pipe10_io_pipe_phv_out_next_config_id; // @[matcher.scala 268:24]
  wire  pipe10_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 268:24]
  wire [63:0] pipe10_io_key_in; // @[matcher.scala 268:24]
  wire [63:0] pipe10_io_key_out; // @[matcher.scala 268:24]
  wire [2:0] pipe10_io_cs_in; // @[matcher.scala 268:24]
  wire [2:0] pipe10_io_cs_out; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_addr_in; // @[matcher.scala 268:24]
  wire  pipe10_io_cs_vec_in_0; // @[matcher.scala 268:24]
  wire  pipe10_io_cs_vec_in_1; // @[matcher.scala 268:24]
  wire  pipe10_io_cs_vec_in_2; // @[matcher.scala 268:24]
  wire  pipe10_io_cs_vec_in_3; // @[matcher.scala 268:24]
  wire  pipe10_io_cs_vec_in_4; // @[matcher.scala 268:24]
  wire  pipe10_io_cs_vec_in_5; // @[matcher.scala 268:24]
  wire  pipe10_io_cs_vec_in_6; // @[matcher.scala 268:24]
  wire  pipe10_io_cs_vec_in_7; // @[matcher.scala 268:24]
  wire [63:0] pipe10_io_data_out_0; // @[matcher.scala 268:24]
  wire [63:0] pipe10_io_data_out_1; // @[matcher.scala 268:24]
  wire [63:0] pipe10_io_data_out_2; // @[matcher.scala 268:24]
  wire [63:0] pipe10_io_data_out_3; // @[matcher.scala 268:24]
  wire [63:0] pipe10_io_data_out_4; // @[matcher.scala 268:24]
  wire [63:0] pipe10_io_data_out_5; // @[matcher.scala 268:24]
  wire [63:0] pipe10_io_data_out_6; // @[matcher.scala 268:24]
  wire [63:0] pipe10_io_data_out_7; // @[matcher.scala 268:24]
  wire  pipe10_io_mem_cluster_0_en; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_mem_cluster_0_addr; // @[matcher.scala 268:24]
  wire [63:0] pipe10_io_mem_cluster_0_data; // @[matcher.scala 268:24]
  wire  pipe10_io_mem_cluster_1_en; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_mem_cluster_1_addr; // @[matcher.scala 268:24]
  wire [63:0] pipe10_io_mem_cluster_1_data; // @[matcher.scala 268:24]
  wire  pipe10_io_mem_cluster_2_en; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_mem_cluster_2_addr; // @[matcher.scala 268:24]
  wire [63:0] pipe10_io_mem_cluster_2_data; // @[matcher.scala 268:24]
  wire  pipe10_io_mem_cluster_3_en; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_mem_cluster_3_addr; // @[matcher.scala 268:24]
  wire [63:0] pipe10_io_mem_cluster_3_data; // @[matcher.scala 268:24]
  wire  pipe10_io_mem_cluster_4_en; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_mem_cluster_4_addr; // @[matcher.scala 268:24]
  wire [63:0] pipe10_io_mem_cluster_4_data; // @[matcher.scala 268:24]
  wire  pipe10_io_mem_cluster_5_en; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_mem_cluster_5_addr; // @[matcher.scala 268:24]
  wire [63:0] pipe10_io_mem_cluster_5_data; // @[matcher.scala 268:24]
  wire  pipe10_io_mem_cluster_6_en; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_mem_cluster_6_addr; // @[matcher.scala 268:24]
  wire [63:0] pipe10_io_mem_cluster_6_data; // @[matcher.scala 268:24]
  wire  pipe10_io_mem_cluster_7_en; // @[matcher.scala 268:24]
  wire [7:0] pipe10_io_mem_cluster_7_addr; // @[matcher.scala 268:24]
  wire [63:0] pipe10_io_mem_cluster_7_data; // @[matcher.scala 268:24]
  wire  pipe11_clock; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_0; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_1; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_2; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_3; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_4; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_5; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_6; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_7; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_8; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_9; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_10; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_11; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_12; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_13; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_14; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_15; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_16; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_17; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_18; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_19; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_20; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_21; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_22; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_23; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_24; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_25; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_26; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_27; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_28; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_29; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_30; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_31; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_32; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_33; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_34; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_35; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_36; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_37; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_38; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_39; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_40; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_41; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_42; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_43; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_44; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_45; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_46; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_47; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_48; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_49; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_50; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_51; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_52; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_53; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_54; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_55; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_56; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_57; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_58; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_59; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_60; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_61; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_62; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_63; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_64; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_65; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_66; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_67; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_68; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_69; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_70; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_71; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_72; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_73; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_74; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_75; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_76; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_77; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_78; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_79; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_80; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_81; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_82; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_83; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_84; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_85; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_86; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_87; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_88; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_89; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_90; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_91; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_92; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_93; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_94; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_95; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_0; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_1; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_2; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_3; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_4; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_5; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_6; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_7; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_8; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_9; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_10; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_11; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_12; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_13; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_14; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_15; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_parse_current_state; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 269:24]
  wire [1:0] pipe11_io_pipe_phv_in_next_processor_id; // @[matcher.scala 269:24]
  wire  pipe11_io_pipe_phv_in_next_config_id; // @[matcher.scala 269:24]
  wire  pipe11_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_0; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_1; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_2; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_3; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_4; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_5; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_6; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_7; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_8; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_9; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_10; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_11; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_12; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_13; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_14; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_15; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_16; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_17; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_18; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_19; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_20; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_21; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_22; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_23; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_24; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_25; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_26; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_27; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_28; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_29; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_30; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_31; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_32; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_33; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_34; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_35; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_36; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_37; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_38; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_39; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_40; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_41; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_42; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_43; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_44; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_45; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_46; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_47; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_48; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_49; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_50; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_51; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_52; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_53; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_54; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_55; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_56; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_57; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_58; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_59; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_60; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_61; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_62; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_63; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_64; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_65; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_66; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_67; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_68; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_69; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_70; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_71; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_72; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_73; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_74; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_75; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_76; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_77; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_78; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_79; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_80; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_81; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_82; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_83; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_84; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_85; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_86; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_87; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_88; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_89; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_90; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_91; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_92; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_93; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_94; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_95; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_0; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_1; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_2; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_3; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_4; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_5; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_6; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_7; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_8; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_9; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_10; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_11; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_12; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_13; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_14; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_15; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_parse_current_state; // @[matcher.scala 269:24]
  wire [7:0] pipe11_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 269:24]
  wire [15:0] pipe11_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 269:24]
  wire [1:0] pipe11_io_pipe_phv_out_next_processor_id; // @[matcher.scala 269:24]
  wire  pipe11_io_pipe_phv_out_next_config_id; // @[matcher.scala 269:24]
  wire  pipe11_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 269:24]
  wire [3:0] pipe11_io_table_config_0_table_width; // @[matcher.scala 269:24]
  wire [3:0] pipe11_io_table_config_0_table_depth; // @[matcher.scala 269:24]
  wire [3:0] pipe11_io_table_config_1_table_width; // @[matcher.scala 269:24]
  wire [3:0] pipe11_io_table_config_1_table_depth; // @[matcher.scala 269:24]
  wire [63:0] pipe11_io_key_in; // @[matcher.scala 269:24]
  wire [63:0] pipe11_io_key_out; // @[matcher.scala 269:24]
  wire [2:0] pipe11_io_cs_in; // @[matcher.scala 269:24]
  wire [63:0] pipe11_io_data_in_0; // @[matcher.scala 269:24]
  wire [63:0] pipe11_io_data_in_1; // @[matcher.scala 269:24]
  wire [63:0] pipe11_io_data_in_2; // @[matcher.scala 269:24]
  wire [63:0] pipe11_io_data_in_3; // @[matcher.scala 269:24]
  wire [63:0] pipe11_io_data_in_4; // @[matcher.scala 269:24]
  wire [63:0] pipe11_io_data_in_5; // @[matcher.scala 269:24]
  wire [63:0] pipe11_io_data_in_6; // @[matcher.scala 269:24]
  wire [63:0] pipe11_io_data_in_7; // @[matcher.scala 269:24]
  wire [127:0] pipe11_io_data_out; // @[matcher.scala 269:24]
  wire  pipe12_clock; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_0; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_1; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_2; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_3; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_4; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_5; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_6; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_7; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_8; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_9; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_10; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_11; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_12; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_13; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_14; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_15; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_16; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_17; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_18; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_19; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_20; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_21; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_22; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_23; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_24; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_25; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_26; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_27; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_28; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_29; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_30; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_31; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_32; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_33; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_34; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_35; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_36; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_37; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_38; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_39; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_40; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_41; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_42; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_43; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_44; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_45; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_46; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_47; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_48; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_49; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_50; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_51; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_52; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_53; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_54; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_55; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_56; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_57; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_58; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_59; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_60; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_61; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_62; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_63; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_64; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_65; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_66; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_67; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_68; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_69; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_70; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_71; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_72; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_73; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_74; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_75; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_76; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_77; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_78; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_79; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_80; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_81; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_82; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_83; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_84; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_85; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_86; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_87; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_88; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_89; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_90; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_91; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_92; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_93; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_94; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_95; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_0; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_1; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_2; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_3; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_4; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_5; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_6; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_7; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_8; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_9; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_10; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_11; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_12; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_13; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_14; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_15; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_parse_current_state; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 270:24]
  wire [1:0] pipe12_io_pipe_phv_in_next_processor_id; // @[matcher.scala 270:24]
  wire  pipe12_io_pipe_phv_in_next_config_id; // @[matcher.scala 270:24]
  wire  pipe12_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_0; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_1; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_2; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_3; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_4; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_5; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_6; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_7; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_8; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_9; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_10; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_11; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_12; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_13; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_14; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_15; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_16; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_17; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_18; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_19; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_20; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_21; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_22; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_23; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_24; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_25; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_26; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_27; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_28; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_29; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_30; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_31; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_32; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_33; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_34; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_35; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_36; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_37; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_38; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_39; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_40; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_41; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_42; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_43; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_44; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_45; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_46; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_47; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_48; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_49; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_50; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_51; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_52; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_53; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_54; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_55; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_56; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_57; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_58; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_59; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_60; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_61; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_62; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_63; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_64; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_65; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_66; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_67; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_68; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_69; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_70; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_71; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_72; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_73; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_74; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_75; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_76; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_77; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_78; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_79; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_80; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_81; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_82; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_83; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_84; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_85; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_86; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_87; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_88; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_89; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_90; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_91; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_92; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_93; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_94; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_95; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_0; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_1; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_2; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_3; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_4; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_5; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_6; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_7; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_8; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_9; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_10; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_11; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_12; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_13; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_14; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_15; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_parse_current_state; // @[matcher.scala 270:24]
  wire [7:0] pipe12_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 270:24]
  wire [15:0] pipe12_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 270:24]
  wire [1:0] pipe12_io_pipe_phv_out_next_processor_id; // @[matcher.scala 270:24]
  wire  pipe12_io_pipe_phv_out_next_config_id; // @[matcher.scala 270:24]
  wire  pipe12_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 270:24]
  wire [3:0] pipe12_io_key_config_0_key_length; // @[matcher.scala 270:24]
  wire [3:0] pipe12_io_key_config_1_key_length; // @[matcher.scala 270:24]
  wire [63:0] pipe12_io_key_in; // @[matcher.scala 270:24]
  wire [127:0] pipe12_io_data_in; // @[matcher.scala 270:24]
  wire  pipe12_io_hit; // @[matcher.scala 270:24]
  wire [63:0] pipe12_io_match_value; // @[matcher.scala 270:24]
  reg [7:0] key_config_0_header_id; // @[matcher.scala 17:25]
  reg [7:0] key_config_0_internal_offset; // @[matcher.scala 17:25]
  reg [3:0] key_config_0_key_length; // @[matcher.scala 17:25]
  reg [7:0] key_config_1_header_id; // @[matcher.scala 17:25]
  reg [7:0] key_config_1_internal_offset; // @[matcher.scala 17:25]
  reg [3:0] key_config_1_key_length; // @[matcher.scala 17:25]
  reg [3:0] table_config_0_table_width; // @[matcher.scala 18:27]
  reg [3:0] table_config_0_table_depth; // @[matcher.scala 18:27]
  reg [3:0] table_config_1_table_width; // @[matcher.scala 18:27]
  reg [3:0] table_config_1_table_depth; // @[matcher.scala 18:27]
  MatchGetOffset pipe1 ( // @[matcher.scala 264:23]
    .clock(pipe1_clock),
    .io_pipe_phv_in_data_0(pipe1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe1_io_pipe_phv_out_is_valid_processor),
    .io_key_config_0_header_id(pipe1_io_key_config_0_header_id),
    .io_key_config_0_internal_offset(pipe1_io_key_config_0_internal_offset),
    .io_key_config_1_header_id(pipe1_io_key_config_1_header_id),
    .io_key_config_1_internal_offset(pipe1_io_key_config_1_internal_offset),
    .io_key_offset(pipe1_io_key_offset)
  );
  MatchGetKey pipe2 ( // @[matcher.scala 265:23]
    .clock(pipe2_clock),
    .io_pipe_phv_in_data_0(pipe2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe2_io_pipe_phv_out_is_valid_processor),
    .io_key_config_0_key_length(pipe2_io_key_config_0_key_length),
    .io_key_config_1_key_length(pipe2_io_key_config_1_key_length),
    .io_key_offset(pipe2_io_key_offset),
    .io_match_key(pipe2_io_match_key)
  );
  Hash pipe3to8 ( // @[matcher.scala 266:26]
    .clock(pipe3to8_clock),
    .io_pipe_phv_in_data_0(pipe3to8_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe3to8_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe3to8_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe3to8_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe3to8_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe3to8_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe3to8_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe3to8_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe3to8_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe3to8_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe3to8_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe3to8_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe3to8_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe3to8_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe3to8_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe3to8_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe3to8_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe3to8_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe3to8_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe3to8_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe3to8_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe3to8_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe3to8_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe3to8_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe3to8_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe3to8_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe3to8_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe3to8_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe3to8_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe3to8_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe3to8_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe3to8_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe3to8_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe3to8_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe3to8_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe3to8_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe3to8_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe3to8_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe3to8_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe3to8_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe3to8_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe3to8_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe3to8_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe3to8_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe3to8_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe3to8_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe3to8_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe3to8_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe3to8_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe3to8_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe3to8_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe3to8_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe3to8_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe3to8_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe3to8_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe3to8_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe3to8_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe3to8_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe3to8_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe3to8_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe3to8_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe3to8_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe3to8_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe3to8_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe3to8_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe3to8_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe3to8_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe3to8_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe3to8_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe3to8_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe3to8_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe3to8_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe3to8_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe3to8_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe3to8_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe3to8_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe3to8_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe3to8_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe3to8_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe3to8_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe3to8_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe3to8_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe3to8_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe3to8_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe3to8_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe3to8_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe3to8_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe3to8_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe3to8_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe3to8_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe3to8_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe3to8_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe3to8_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe3to8_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe3to8_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe3to8_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe3to8_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe3to8_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe3to8_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe3to8_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe3to8_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe3to8_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe3to8_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe3to8_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe3to8_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe3to8_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe3to8_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe3to8_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe3to8_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe3to8_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe3to8_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe3to8_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe3to8_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe3to8_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe3to8_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe3to8_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe3to8_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe3to8_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe3to8_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe3to8_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe3to8_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe3to8_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe3to8_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe3to8_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe3to8_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe3to8_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe3to8_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe3to8_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe3to8_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe3to8_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe3to8_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe3to8_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe3to8_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe3to8_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe3to8_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe3to8_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe3to8_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe3to8_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe3to8_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe3to8_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe3to8_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe3to8_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe3to8_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe3to8_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe3to8_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe3to8_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe3to8_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe3to8_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe3to8_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe3to8_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe3to8_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe3to8_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe3to8_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe3to8_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe3to8_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe3to8_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe3to8_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe3to8_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe3to8_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe3to8_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe3to8_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe3to8_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe3to8_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe3to8_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe3to8_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe3to8_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe3to8_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe3to8_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe3to8_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe3to8_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe3to8_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe3to8_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe3to8_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe3to8_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe3to8_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe3to8_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe3to8_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe3to8_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe3to8_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe3to8_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe3to8_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe3to8_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe3to8_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe3to8_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe3to8_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe3to8_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe3to8_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe3to8_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe3to8_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe3to8_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe3to8_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe3to8_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe3to8_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe3to8_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe3to8_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe3to8_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe3to8_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe3to8_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe3to8_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe3to8_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe3to8_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe3to8_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe3to8_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe3to8_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe3to8_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe3to8_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe3to8_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe3to8_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe3to8_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe3to8_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe3to8_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe3to8_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe3to8_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe3to8_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe3to8_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe3to8_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe3to8_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe3to8_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe3to8_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe3to8_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe3to8_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe3to8_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe3to8_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe3to8_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe3to8_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe3to8_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe3to8_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe3to8_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe3to8_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe3to8_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe3to8_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe3to8_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe3to8_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe3to8_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe3to8_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe3to8_io_pipe_phv_out_is_valid_processor),
    .io_mod_hash_depth_mod(pipe3to8_io_mod_hash_depth_mod),
    .io_mod_config_id(pipe3to8_io_mod_config_id),
    .io_mod_hash_depth(pipe3to8_io_mod_hash_depth),
    .io_key_in(pipe3to8_io_key_in),
    .io_key_out(pipe3to8_io_key_out),
    .io_hash_val(pipe3to8_io_hash_val),
    .io_hash_val_cs(pipe3to8_io_hash_val_cs)
  );
  MatchGetCs pipe9 ( // @[matcher.scala 267:23]
    .clock(pipe9_clock),
    .io_pipe_phv_in_data_0(pipe9_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe9_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe9_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe9_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe9_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe9_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe9_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe9_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe9_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe9_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe9_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe9_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe9_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe9_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe9_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe9_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe9_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe9_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe9_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe9_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe9_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe9_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe9_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe9_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe9_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe9_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe9_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe9_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe9_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe9_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe9_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe9_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe9_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe9_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe9_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe9_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe9_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe9_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe9_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe9_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe9_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe9_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe9_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe9_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe9_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe9_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe9_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe9_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe9_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe9_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe9_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe9_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe9_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe9_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe9_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe9_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe9_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe9_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe9_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe9_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe9_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe9_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe9_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe9_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe9_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe9_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe9_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe9_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe9_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe9_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe9_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe9_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe9_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe9_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe9_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe9_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe9_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe9_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe9_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe9_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe9_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe9_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe9_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe9_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe9_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe9_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe9_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe9_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe9_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe9_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe9_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe9_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe9_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe9_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe9_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe9_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe9_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe9_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe9_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe9_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe9_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe9_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe9_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe9_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe9_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe9_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe9_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe9_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe9_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe9_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe9_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe9_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe9_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe9_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe9_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe9_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe9_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe9_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe9_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe9_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe9_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe9_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe9_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe9_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe9_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe9_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe9_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe9_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe9_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe9_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe9_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe9_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe9_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe9_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe9_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe9_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe9_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe9_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe9_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe9_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe9_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe9_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe9_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe9_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe9_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe9_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe9_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe9_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe9_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe9_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe9_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe9_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe9_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe9_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe9_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe9_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe9_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe9_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe9_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe9_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe9_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe9_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe9_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe9_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe9_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe9_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe9_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe9_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe9_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe9_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe9_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe9_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe9_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe9_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe9_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe9_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe9_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe9_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe9_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe9_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe9_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe9_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe9_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe9_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe9_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe9_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe9_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe9_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe9_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe9_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe9_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe9_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe9_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe9_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe9_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe9_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe9_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe9_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe9_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe9_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe9_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe9_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe9_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe9_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe9_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe9_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe9_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe9_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe9_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe9_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe9_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe9_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe9_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe9_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe9_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe9_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe9_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe9_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe9_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe9_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe9_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe9_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe9_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe9_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe9_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe9_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe9_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe9_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe9_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe9_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe9_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe9_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe9_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe9_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe9_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe9_io_pipe_phv_out_is_valid_processor),
    .io_table_config_0_table_width(pipe9_io_table_config_0_table_width),
    .io_table_config_0_table_depth(pipe9_io_table_config_0_table_depth),
    .io_table_config_1_table_width(pipe9_io_table_config_1_table_width),
    .io_table_config_1_table_depth(pipe9_io_table_config_1_table_depth),
    .io_key_in(pipe9_io_key_in),
    .io_key_out(pipe9_io_key_out),
    .io_addr_in(pipe9_io_addr_in),
    .io_addr_out(pipe9_io_addr_out),
    .io_cs_in(pipe9_io_cs_in),
    .io_cs_out(pipe9_io_cs_out),
    .io_cs_vec_out_0(pipe9_io_cs_vec_out_0),
    .io_cs_vec_out_1(pipe9_io_cs_vec_out_1),
    .io_cs_vec_out_2(pipe9_io_cs_vec_out_2),
    .io_cs_vec_out_3(pipe9_io_cs_vec_out_3),
    .io_cs_vec_out_4(pipe9_io_cs_vec_out_4),
    .io_cs_vec_out_5(pipe9_io_cs_vec_out_5),
    .io_cs_vec_out_6(pipe9_io_cs_vec_out_6),
    .io_cs_vec_out_7(pipe9_io_cs_vec_out_7)
  );
  MatchReadData pipe10 ( // @[matcher.scala 268:24]
    .clock(pipe10_clock),
    .io_pipe_phv_in_data_0(pipe10_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe10_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe10_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe10_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe10_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe10_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe10_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe10_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe10_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe10_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe10_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe10_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe10_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe10_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe10_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe10_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe10_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe10_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe10_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe10_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe10_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe10_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe10_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe10_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe10_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe10_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe10_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe10_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe10_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe10_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe10_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe10_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe10_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe10_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe10_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe10_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe10_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe10_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe10_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe10_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe10_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe10_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe10_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe10_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe10_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe10_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe10_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe10_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe10_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe10_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe10_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe10_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe10_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe10_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe10_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe10_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe10_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe10_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe10_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe10_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe10_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe10_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe10_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe10_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe10_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe10_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe10_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe10_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe10_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe10_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe10_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe10_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe10_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe10_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe10_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe10_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe10_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe10_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe10_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe10_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe10_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe10_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe10_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe10_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe10_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe10_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe10_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe10_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe10_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe10_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe10_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe10_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe10_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe10_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe10_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe10_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe10_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe10_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe10_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe10_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe10_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe10_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe10_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe10_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe10_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe10_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe10_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe10_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe10_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe10_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe10_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe10_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe10_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe10_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe10_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe10_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe10_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe10_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe10_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe10_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe10_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe10_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe10_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe10_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe10_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe10_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe10_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe10_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe10_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe10_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe10_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe10_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe10_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe10_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe10_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe10_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe10_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe10_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe10_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe10_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe10_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe10_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe10_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe10_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe10_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe10_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe10_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe10_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe10_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe10_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe10_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe10_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe10_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe10_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe10_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe10_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe10_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe10_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe10_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe10_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe10_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe10_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe10_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe10_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe10_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe10_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe10_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe10_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe10_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe10_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe10_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe10_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe10_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe10_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe10_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe10_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe10_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe10_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe10_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe10_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe10_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe10_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe10_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe10_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe10_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe10_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe10_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe10_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe10_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe10_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe10_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe10_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe10_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe10_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe10_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe10_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe10_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe10_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe10_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe10_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe10_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe10_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe10_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe10_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe10_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe10_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe10_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe10_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe10_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe10_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe10_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe10_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe10_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe10_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe10_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe10_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe10_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe10_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe10_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe10_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe10_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe10_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe10_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe10_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe10_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe10_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe10_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe10_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe10_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe10_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe10_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe10_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe10_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe10_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe10_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe10_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe10_io_key_in),
    .io_key_out(pipe10_io_key_out),
    .io_cs_in(pipe10_io_cs_in),
    .io_cs_out(pipe10_io_cs_out),
    .io_addr_in(pipe10_io_addr_in),
    .io_cs_vec_in_0(pipe10_io_cs_vec_in_0),
    .io_cs_vec_in_1(pipe10_io_cs_vec_in_1),
    .io_cs_vec_in_2(pipe10_io_cs_vec_in_2),
    .io_cs_vec_in_3(pipe10_io_cs_vec_in_3),
    .io_cs_vec_in_4(pipe10_io_cs_vec_in_4),
    .io_cs_vec_in_5(pipe10_io_cs_vec_in_5),
    .io_cs_vec_in_6(pipe10_io_cs_vec_in_6),
    .io_cs_vec_in_7(pipe10_io_cs_vec_in_7),
    .io_data_out_0(pipe10_io_data_out_0),
    .io_data_out_1(pipe10_io_data_out_1),
    .io_data_out_2(pipe10_io_data_out_2),
    .io_data_out_3(pipe10_io_data_out_3),
    .io_data_out_4(pipe10_io_data_out_4),
    .io_data_out_5(pipe10_io_data_out_5),
    .io_data_out_6(pipe10_io_data_out_6),
    .io_data_out_7(pipe10_io_data_out_7),
    .io_mem_cluster_0_en(pipe10_io_mem_cluster_0_en),
    .io_mem_cluster_0_addr(pipe10_io_mem_cluster_0_addr),
    .io_mem_cluster_0_data(pipe10_io_mem_cluster_0_data),
    .io_mem_cluster_1_en(pipe10_io_mem_cluster_1_en),
    .io_mem_cluster_1_addr(pipe10_io_mem_cluster_1_addr),
    .io_mem_cluster_1_data(pipe10_io_mem_cluster_1_data),
    .io_mem_cluster_2_en(pipe10_io_mem_cluster_2_en),
    .io_mem_cluster_2_addr(pipe10_io_mem_cluster_2_addr),
    .io_mem_cluster_2_data(pipe10_io_mem_cluster_2_data),
    .io_mem_cluster_3_en(pipe10_io_mem_cluster_3_en),
    .io_mem_cluster_3_addr(pipe10_io_mem_cluster_3_addr),
    .io_mem_cluster_3_data(pipe10_io_mem_cluster_3_data),
    .io_mem_cluster_4_en(pipe10_io_mem_cluster_4_en),
    .io_mem_cluster_4_addr(pipe10_io_mem_cluster_4_addr),
    .io_mem_cluster_4_data(pipe10_io_mem_cluster_4_data),
    .io_mem_cluster_5_en(pipe10_io_mem_cluster_5_en),
    .io_mem_cluster_5_addr(pipe10_io_mem_cluster_5_addr),
    .io_mem_cluster_5_data(pipe10_io_mem_cluster_5_data),
    .io_mem_cluster_6_en(pipe10_io_mem_cluster_6_en),
    .io_mem_cluster_6_addr(pipe10_io_mem_cluster_6_addr),
    .io_mem_cluster_6_data(pipe10_io_mem_cluster_6_data),
    .io_mem_cluster_7_en(pipe10_io_mem_cluster_7_en),
    .io_mem_cluster_7_addr(pipe10_io_mem_cluster_7_addr),
    .io_mem_cluster_7_data(pipe10_io_mem_cluster_7_data)
  );
  MatchDataReshape pipe11 ( // @[matcher.scala 269:24]
    .clock(pipe11_clock),
    .io_pipe_phv_in_data_0(pipe11_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe11_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe11_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe11_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe11_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe11_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe11_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe11_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe11_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe11_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe11_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe11_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe11_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe11_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe11_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe11_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe11_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe11_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe11_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe11_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe11_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe11_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe11_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe11_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe11_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe11_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe11_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe11_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe11_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe11_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe11_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe11_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe11_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe11_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe11_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe11_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe11_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe11_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe11_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe11_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe11_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe11_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe11_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe11_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe11_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe11_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe11_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe11_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe11_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe11_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe11_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe11_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe11_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe11_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe11_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe11_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe11_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe11_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe11_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe11_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe11_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe11_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe11_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe11_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe11_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe11_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe11_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe11_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe11_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe11_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe11_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe11_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe11_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe11_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe11_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe11_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe11_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe11_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe11_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe11_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe11_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe11_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe11_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe11_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe11_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe11_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe11_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe11_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe11_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe11_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe11_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe11_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe11_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe11_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe11_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe11_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe11_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe11_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe11_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe11_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe11_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe11_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe11_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe11_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe11_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe11_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe11_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe11_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe11_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe11_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe11_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe11_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe11_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe11_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe11_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe11_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe11_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe11_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe11_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe11_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe11_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe11_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe11_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe11_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe11_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe11_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe11_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe11_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe11_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe11_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe11_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe11_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe11_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe11_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe11_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe11_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe11_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe11_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe11_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe11_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe11_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe11_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe11_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe11_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe11_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe11_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe11_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe11_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe11_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe11_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe11_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe11_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe11_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe11_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe11_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe11_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe11_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe11_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe11_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe11_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe11_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe11_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe11_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe11_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe11_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe11_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe11_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe11_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe11_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe11_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe11_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe11_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe11_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe11_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe11_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe11_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe11_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe11_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe11_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe11_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe11_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe11_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe11_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe11_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe11_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe11_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe11_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe11_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe11_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe11_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe11_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe11_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe11_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe11_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe11_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe11_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe11_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe11_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe11_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe11_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe11_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe11_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe11_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe11_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe11_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe11_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe11_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe11_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe11_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe11_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe11_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe11_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe11_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe11_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe11_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe11_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe11_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe11_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe11_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe11_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe11_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe11_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe11_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe11_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe11_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe11_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe11_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe11_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe11_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe11_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe11_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe11_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe11_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe11_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe11_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe11_io_pipe_phv_out_is_valid_processor),
    .io_table_config_0_table_width(pipe11_io_table_config_0_table_width),
    .io_table_config_0_table_depth(pipe11_io_table_config_0_table_depth),
    .io_table_config_1_table_width(pipe11_io_table_config_1_table_width),
    .io_table_config_1_table_depth(pipe11_io_table_config_1_table_depth),
    .io_key_in(pipe11_io_key_in),
    .io_key_out(pipe11_io_key_out),
    .io_cs_in(pipe11_io_cs_in),
    .io_data_in_0(pipe11_io_data_in_0),
    .io_data_in_1(pipe11_io_data_in_1),
    .io_data_in_2(pipe11_io_data_in_2),
    .io_data_in_3(pipe11_io_data_in_3),
    .io_data_in_4(pipe11_io_data_in_4),
    .io_data_in_5(pipe11_io_data_in_5),
    .io_data_in_6(pipe11_io_data_in_6),
    .io_data_in_7(pipe11_io_data_in_7),
    .io_data_out(pipe11_io_data_out)
  );
  MatchResult pipe12 ( // @[matcher.scala 270:24]
    .clock(pipe12_clock),
    .io_pipe_phv_in_data_0(pipe12_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe12_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe12_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe12_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe12_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe12_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe12_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe12_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe12_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe12_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe12_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe12_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe12_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe12_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe12_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe12_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe12_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe12_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe12_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe12_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe12_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe12_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe12_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe12_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe12_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe12_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe12_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe12_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe12_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe12_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe12_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe12_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe12_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe12_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe12_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe12_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe12_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe12_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe12_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe12_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe12_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe12_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe12_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe12_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe12_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe12_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe12_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe12_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe12_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe12_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe12_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe12_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe12_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe12_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe12_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe12_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe12_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe12_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe12_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe12_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe12_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe12_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe12_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe12_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe12_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe12_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe12_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe12_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe12_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe12_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe12_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe12_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe12_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe12_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe12_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe12_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe12_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe12_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe12_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe12_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe12_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe12_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe12_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe12_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe12_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe12_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe12_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe12_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe12_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe12_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe12_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe12_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe12_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe12_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe12_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe12_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe12_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe12_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe12_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe12_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe12_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe12_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe12_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe12_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe12_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe12_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe12_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe12_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe12_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe12_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe12_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe12_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe12_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe12_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe12_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe12_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe12_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe12_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe12_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe12_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe12_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe12_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe12_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe12_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe12_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe12_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe12_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe12_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe12_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe12_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe12_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe12_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe12_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe12_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe12_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe12_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe12_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe12_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe12_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe12_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe12_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe12_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe12_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe12_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe12_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe12_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe12_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe12_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe12_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe12_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe12_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe12_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe12_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe12_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe12_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe12_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe12_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe12_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe12_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe12_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe12_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe12_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe12_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe12_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe12_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe12_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe12_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe12_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe12_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe12_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe12_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe12_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe12_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe12_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe12_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe12_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe12_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe12_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe12_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe12_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe12_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe12_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe12_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe12_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe12_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe12_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe12_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe12_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe12_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe12_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe12_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe12_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe12_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe12_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe12_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe12_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe12_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe12_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe12_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe12_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe12_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe12_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe12_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe12_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe12_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe12_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe12_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe12_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe12_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe12_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe12_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe12_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe12_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe12_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe12_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe12_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe12_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe12_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe12_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe12_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe12_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe12_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe12_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe12_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe12_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe12_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe12_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe12_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe12_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe12_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe12_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe12_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe12_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe12_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe12_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe12_io_pipe_phv_out_is_valid_processor),
    .io_key_config_0_key_length(pipe12_io_key_config_0_key_length),
    .io_key_config_1_key_length(pipe12_io_key_config_1_key_length),
    .io_key_in(pipe12_io_key_in),
    .io_data_in(pipe12_io_data_in),
    .io_hit(pipe12_io_hit),
    .io_match_value(pipe12_io_match_value)
  );
  assign io_pipe_phv_out_data_0 = pipe12_io_pipe_phv_out_data_0; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_1 = pipe12_io_pipe_phv_out_data_1; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_2 = pipe12_io_pipe_phv_out_data_2; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_3 = pipe12_io_pipe_phv_out_data_3; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_4 = pipe12_io_pipe_phv_out_data_4; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_5 = pipe12_io_pipe_phv_out_data_5; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_6 = pipe12_io_pipe_phv_out_data_6; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_7 = pipe12_io_pipe_phv_out_data_7; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_8 = pipe12_io_pipe_phv_out_data_8; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_9 = pipe12_io_pipe_phv_out_data_9; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_10 = pipe12_io_pipe_phv_out_data_10; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_11 = pipe12_io_pipe_phv_out_data_11; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_12 = pipe12_io_pipe_phv_out_data_12; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_13 = pipe12_io_pipe_phv_out_data_13; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_14 = pipe12_io_pipe_phv_out_data_14; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_15 = pipe12_io_pipe_phv_out_data_15; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_16 = pipe12_io_pipe_phv_out_data_16; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_17 = pipe12_io_pipe_phv_out_data_17; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_18 = pipe12_io_pipe_phv_out_data_18; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_19 = pipe12_io_pipe_phv_out_data_19; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_20 = pipe12_io_pipe_phv_out_data_20; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_21 = pipe12_io_pipe_phv_out_data_21; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_22 = pipe12_io_pipe_phv_out_data_22; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_23 = pipe12_io_pipe_phv_out_data_23; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_24 = pipe12_io_pipe_phv_out_data_24; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_25 = pipe12_io_pipe_phv_out_data_25; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_26 = pipe12_io_pipe_phv_out_data_26; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_27 = pipe12_io_pipe_phv_out_data_27; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_28 = pipe12_io_pipe_phv_out_data_28; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_29 = pipe12_io_pipe_phv_out_data_29; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_30 = pipe12_io_pipe_phv_out_data_30; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_31 = pipe12_io_pipe_phv_out_data_31; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_32 = pipe12_io_pipe_phv_out_data_32; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_33 = pipe12_io_pipe_phv_out_data_33; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_34 = pipe12_io_pipe_phv_out_data_34; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_35 = pipe12_io_pipe_phv_out_data_35; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_36 = pipe12_io_pipe_phv_out_data_36; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_37 = pipe12_io_pipe_phv_out_data_37; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_38 = pipe12_io_pipe_phv_out_data_38; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_39 = pipe12_io_pipe_phv_out_data_39; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_40 = pipe12_io_pipe_phv_out_data_40; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_41 = pipe12_io_pipe_phv_out_data_41; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_42 = pipe12_io_pipe_phv_out_data_42; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_43 = pipe12_io_pipe_phv_out_data_43; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_44 = pipe12_io_pipe_phv_out_data_44; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_45 = pipe12_io_pipe_phv_out_data_45; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_46 = pipe12_io_pipe_phv_out_data_46; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_47 = pipe12_io_pipe_phv_out_data_47; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_48 = pipe12_io_pipe_phv_out_data_48; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_49 = pipe12_io_pipe_phv_out_data_49; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_50 = pipe12_io_pipe_phv_out_data_50; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_51 = pipe12_io_pipe_phv_out_data_51; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_52 = pipe12_io_pipe_phv_out_data_52; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_53 = pipe12_io_pipe_phv_out_data_53; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_54 = pipe12_io_pipe_phv_out_data_54; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_55 = pipe12_io_pipe_phv_out_data_55; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_56 = pipe12_io_pipe_phv_out_data_56; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_57 = pipe12_io_pipe_phv_out_data_57; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_58 = pipe12_io_pipe_phv_out_data_58; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_59 = pipe12_io_pipe_phv_out_data_59; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_60 = pipe12_io_pipe_phv_out_data_60; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_61 = pipe12_io_pipe_phv_out_data_61; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_62 = pipe12_io_pipe_phv_out_data_62; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_63 = pipe12_io_pipe_phv_out_data_63; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_64 = pipe12_io_pipe_phv_out_data_64; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_65 = pipe12_io_pipe_phv_out_data_65; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_66 = pipe12_io_pipe_phv_out_data_66; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_67 = pipe12_io_pipe_phv_out_data_67; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_68 = pipe12_io_pipe_phv_out_data_68; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_69 = pipe12_io_pipe_phv_out_data_69; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_70 = pipe12_io_pipe_phv_out_data_70; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_71 = pipe12_io_pipe_phv_out_data_71; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_72 = pipe12_io_pipe_phv_out_data_72; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_73 = pipe12_io_pipe_phv_out_data_73; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_74 = pipe12_io_pipe_phv_out_data_74; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_75 = pipe12_io_pipe_phv_out_data_75; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_76 = pipe12_io_pipe_phv_out_data_76; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_77 = pipe12_io_pipe_phv_out_data_77; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_78 = pipe12_io_pipe_phv_out_data_78; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_79 = pipe12_io_pipe_phv_out_data_79; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_80 = pipe12_io_pipe_phv_out_data_80; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_81 = pipe12_io_pipe_phv_out_data_81; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_82 = pipe12_io_pipe_phv_out_data_82; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_83 = pipe12_io_pipe_phv_out_data_83; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_84 = pipe12_io_pipe_phv_out_data_84; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_85 = pipe12_io_pipe_phv_out_data_85; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_86 = pipe12_io_pipe_phv_out_data_86; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_87 = pipe12_io_pipe_phv_out_data_87; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_88 = pipe12_io_pipe_phv_out_data_88; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_89 = pipe12_io_pipe_phv_out_data_89; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_90 = pipe12_io_pipe_phv_out_data_90; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_91 = pipe12_io_pipe_phv_out_data_91; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_92 = pipe12_io_pipe_phv_out_data_92; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_93 = pipe12_io_pipe_phv_out_data_93; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_94 = pipe12_io_pipe_phv_out_data_94; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_data_95 = pipe12_io_pipe_phv_out_data_95; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_header_0 = pipe12_io_pipe_phv_out_header_0; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_header_1 = pipe12_io_pipe_phv_out_header_1; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_header_2 = pipe12_io_pipe_phv_out_header_2; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_header_3 = pipe12_io_pipe_phv_out_header_3; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_header_4 = pipe12_io_pipe_phv_out_header_4; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_header_5 = pipe12_io_pipe_phv_out_header_5; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_header_6 = pipe12_io_pipe_phv_out_header_6; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_header_7 = pipe12_io_pipe_phv_out_header_7; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_header_8 = pipe12_io_pipe_phv_out_header_8; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_header_9 = pipe12_io_pipe_phv_out_header_9; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_header_10 = pipe12_io_pipe_phv_out_header_10; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_header_11 = pipe12_io_pipe_phv_out_header_11; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_header_12 = pipe12_io_pipe_phv_out_header_12; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_header_13 = pipe12_io_pipe_phv_out_header_13; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_header_14 = pipe12_io_pipe_phv_out_header_14; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_header_15 = pipe12_io_pipe_phv_out_header_15; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_parse_current_state = pipe12_io_pipe_phv_out_parse_current_state; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_parse_current_offset = pipe12_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_parse_transition_field = pipe12_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_next_processor_id = pipe12_io_pipe_phv_out_next_processor_id; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_next_config_id = pipe12_io_pipe_phv_out_next_config_id; // @[matcher.scala 309:27]
  assign io_pipe_phv_out_is_valid_processor = pipe12_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 309:27]
  assign io_hit = pipe12_io_hit; // @[matcher.scala 310:27]
  assign io_match_value = pipe12_io_match_value; // @[matcher.scala 311:27]
  assign io_mem_cluster_0_en = pipe10_io_mem_cluster_0_en; // @[matcher.scala 296:27]
  assign io_mem_cluster_0_addr = pipe10_io_mem_cluster_0_addr; // @[matcher.scala 296:27]
  assign io_mem_cluster_1_en = pipe10_io_mem_cluster_1_en; // @[matcher.scala 296:27]
  assign io_mem_cluster_1_addr = pipe10_io_mem_cluster_1_addr; // @[matcher.scala 296:27]
  assign io_mem_cluster_2_en = pipe10_io_mem_cluster_2_en; // @[matcher.scala 296:27]
  assign io_mem_cluster_2_addr = pipe10_io_mem_cluster_2_addr; // @[matcher.scala 296:27]
  assign io_mem_cluster_3_en = pipe10_io_mem_cluster_3_en; // @[matcher.scala 296:27]
  assign io_mem_cluster_3_addr = pipe10_io_mem_cluster_3_addr; // @[matcher.scala 296:27]
  assign io_mem_cluster_4_en = pipe10_io_mem_cluster_4_en; // @[matcher.scala 296:27]
  assign io_mem_cluster_4_addr = pipe10_io_mem_cluster_4_addr; // @[matcher.scala 296:27]
  assign io_mem_cluster_5_en = pipe10_io_mem_cluster_5_en; // @[matcher.scala 296:27]
  assign io_mem_cluster_5_addr = pipe10_io_mem_cluster_5_addr; // @[matcher.scala 296:27]
  assign io_mem_cluster_6_en = pipe10_io_mem_cluster_6_en; // @[matcher.scala 296:27]
  assign io_mem_cluster_6_addr = pipe10_io_mem_cluster_6_addr; // @[matcher.scala 296:27]
  assign io_mem_cluster_7_en = pipe10_io_mem_cluster_7_en; // @[matcher.scala 296:27]
  assign io_mem_cluster_7_addr = pipe10_io_mem_cluster_7_addr; // @[matcher.scala 296:27]
  assign pipe1_clock = clock;
  assign pipe1_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[matcher.scala 272:26]
  assign pipe1_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[matcher.scala 272:26]
  assign pipe1_io_key_config_0_header_id = key_config_0_header_id; // @[matcher.scala 273:26]
  assign pipe1_io_key_config_0_internal_offset = key_config_0_internal_offset; // @[matcher.scala 273:26]
  assign pipe1_io_key_config_1_header_id = key_config_1_header_id; // @[matcher.scala 273:26]
  assign pipe1_io_key_config_1_internal_offset = key_config_1_internal_offset; // @[matcher.scala 273:26]
  assign pipe2_clock = clock;
  assign pipe2_io_pipe_phv_in_data_0 = pipe1_io_pipe_phv_out_data_0; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_1 = pipe1_io_pipe_phv_out_data_1; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_2 = pipe1_io_pipe_phv_out_data_2; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_3 = pipe1_io_pipe_phv_out_data_3; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_4 = pipe1_io_pipe_phv_out_data_4; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_5 = pipe1_io_pipe_phv_out_data_5; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_6 = pipe1_io_pipe_phv_out_data_6; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_7 = pipe1_io_pipe_phv_out_data_7; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_8 = pipe1_io_pipe_phv_out_data_8; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_9 = pipe1_io_pipe_phv_out_data_9; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_10 = pipe1_io_pipe_phv_out_data_10; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_11 = pipe1_io_pipe_phv_out_data_11; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_12 = pipe1_io_pipe_phv_out_data_12; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_13 = pipe1_io_pipe_phv_out_data_13; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_14 = pipe1_io_pipe_phv_out_data_14; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_15 = pipe1_io_pipe_phv_out_data_15; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_16 = pipe1_io_pipe_phv_out_data_16; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_17 = pipe1_io_pipe_phv_out_data_17; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_18 = pipe1_io_pipe_phv_out_data_18; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_19 = pipe1_io_pipe_phv_out_data_19; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_20 = pipe1_io_pipe_phv_out_data_20; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_21 = pipe1_io_pipe_phv_out_data_21; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_22 = pipe1_io_pipe_phv_out_data_22; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_23 = pipe1_io_pipe_phv_out_data_23; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_24 = pipe1_io_pipe_phv_out_data_24; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_25 = pipe1_io_pipe_phv_out_data_25; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_26 = pipe1_io_pipe_phv_out_data_26; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_27 = pipe1_io_pipe_phv_out_data_27; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_28 = pipe1_io_pipe_phv_out_data_28; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_29 = pipe1_io_pipe_phv_out_data_29; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_30 = pipe1_io_pipe_phv_out_data_30; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_31 = pipe1_io_pipe_phv_out_data_31; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_32 = pipe1_io_pipe_phv_out_data_32; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_33 = pipe1_io_pipe_phv_out_data_33; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_34 = pipe1_io_pipe_phv_out_data_34; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_35 = pipe1_io_pipe_phv_out_data_35; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_36 = pipe1_io_pipe_phv_out_data_36; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_37 = pipe1_io_pipe_phv_out_data_37; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_38 = pipe1_io_pipe_phv_out_data_38; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_39 = pipe1_io_pipe_phv_out_data_39; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_40 = pipe1_io_pipe_phv_out_data_40; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_41 = pipe1_io_pipe_phv_out_data_41; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_42 = pipe1_io_pipe_phv_out_data_42; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_43 = pipe1_io_pipe_phv_out_data_43; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_44 = pipe1_io_pipe_phv_out_data_44; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_45 = pipe1_io_pipe_phv_out_data_45; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_46 = pipe1_io_pipe_phv_out_data_46; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_47 = pipe1_io_pipe_phv_out_data_47; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_48 = pipe1_io_pipe_phv_out_data_48; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_49 = pipe1_io_pipe_phv_out_data_49; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_50 = pipe1_io_pipe_phv_out_data_50; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_51 = pipe1_io_pipe_phv_out_data_51; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_52 = pipe1_io_pipe_phv_out_data_52; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_53 = pipe1_io_pipe_phv_out_data_53; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_54 = pipe1_io_pipe_phv_out_data_54; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_55 = pipe1_io_pipe_phv_out_data_55; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_56 = pipe1_io_pipe_phv_out_data_56; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_57 = pipe1_io_pipe_phv_out_data_57; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_58 = pipe1_io_pipe_phv_out_data_58; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_59 = pipe1_io_pipe_phv_out_data_59; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_60 = pipe1_io_pipe_phv_out_data_60; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_61 = pipe1_io_pipe_phv_out_data_61; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_62 = pipe1_io_pipe_phv_out_data_62; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_63 = pipe1_io_pipe_phv_out_data_63; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_64 = pipe1_io_pipe_phv_out_data_64; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_65 = pipe1_io_pipe_phv_out_data_65; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_66 = pipe1_io_pipe_phv_out_data_66; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_67 = pipe1_io_pipe_phv_out_data_67; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_68 = pipe1_io_pipe_phv_out_data_68; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_69 = pipe1_io_pipe_phv_out_data_69; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_70 = pipe1_io_pipe_phv_out_data_70; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_71 = pipe1_io_pipe_phv_out_data_71; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_72 = pipe1_io_pipe_phv_out_data_72; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_73 = pipe1_io_pipe_phv_out_data_73; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_74 = pipe1_io_pipe_phv_out_data_74; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_75 = pipe1_io_pipe_phv_out_data_75; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_76 = pipe1_io_pipe_phv_out_data_76; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_77 = pipe1_io_pipe_phv_out_data_77; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_78 = pipe1_io_pipe_phv_out_data_78; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_79 = pipe1_io_pipe_phv_out_data_79; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_80 = pipe1_io_pipe_phv_out_data_80; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_81 = pipe1_io_pipe_phv_out_data_81; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_82 = pipe1_io_pipe_phv_out_data_82; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_83 = pipe1_io_pipe_phv_out_data_83; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_84 = pipe1_io_pipe_phv_out_data_84; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_85 = pipe1_io_pipe_phv_out_data_85; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_86 = pipe1_io_pipe_phv_out_data_86; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_87 = pipe1_io_pipe_phv_out_data_87; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_88 = pipe1_io_pipe_phv_out_data_88; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_89 = pipe1_io_pipe_phv_out_data_89; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_90 = pipe1_io_pipe_phv_out_data_90; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_91 = pipe1_io_pipe_phv_out_data_91; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_92 = pipe1_io_pipe_phv_out_data_92; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_93 = pipe1_io_pipe_phv_out_data_93; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_94 = pipe1_io_pipe_phv_out_data_94; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_data_95 = pipe1_io_pipe_phv_out_data_95; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_header_0 = pipe1_io_pipe_phv_out_header_0; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_header_1 = pipe1_io_pipe_phv_out_header_1; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_header_2 = pipe1_io_pipe_phv_out_header_2; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_header_3 = pipe1_io_pipe_phv_out_header_3; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_header_4 = pipe1_io_pipe_phv_out_header_4; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_header_5 = pipe1_io_pipe_phv_out_header_5; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_header_6 = pipe1_io_pipe_phv_out_header_6; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_header_7 = pipe1_io_pipe_phv_out_header_7; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_header_8 = pipe1_io_pipe_phv_out_header_8; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_header_9 = pipe1_io_pipe_phv_out_header_9; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_header_10 = pipe1_io_pipe_phv_out_header_10; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_header_11 = pipe1_io_pipe_phv_out_header_11; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_header_12 = pipe1_io_pipe_phv_out_header_12; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_header_13 = pipe1_io_pipe_phv_out_header_13; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_header_14 = pipe1_io_pipe_phv_out_header_14; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_header_15 = pipe1_io_pipe_phv_out_header_15; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_parse_current_state = pipe1_io_pipe_phv_out_parse_current_state; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_parse_current_offset = pipe1_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_parse_transition_field = pipe1_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_next_processor_id = pipe1_io_pipe_phv_out_next_processor_id; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_next_config_id = pipe1_io_pipe_phv_out_next_config_id; // @[matcher.scala 275:26]
  assign pipe2_io_pipe_phv_in_is_valid_processor = pipe1_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 275:26]
  assign pipe2_io_key_config_0_key_length = key_config_0_key_length; // @[matcher.scala 277:26]
  assign pipe2_io_key_config_1_key_length = key_config_1_key_length; // @[matcher.scala 277:26]
  assign pipe2_io_key_offset = pipe1_io_key_offset; // @[matcher.scala 276:26]
  assign pipe3to8_clock = clock;
  assign pipe3to8_io_pipe_phv_in_data_0 = pipe2_io_pipe_phv_out_data_0; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_1 = pipe2_io_pipe_phv_out_data_1; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_2 = pipe2_io_pipe_phv_out_data_2; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_3 = pipe2_io_pipe_phv_out_data_3; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_4 = pipe2_io_pipe_phv_out_data_4; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_5 = pipe2_io_pipe_phv_out_data_5; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_6 = pipe2_io_pipe_phv_out_data_6; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_7 = pipe2_io_pipe_phv_out_data_7; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_8 = pipe2_io_pipe_phv_out_data_8; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_9 = pipe2_io_pipe_phv_out_data_9; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_10 = pipe2_io_pipe_phv_out_data_10; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_11 = pipe2_io_pipe_phv_out_data_11; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_12 = pipe2_io_pipe_phv_out_data_12; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_13 = pipe2_io_pipe_phv_out_data_13; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_14 = pipe2_io_pipe_phv_out_data_14; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_15 = pipe2_io_pipe_phv_out_data_15; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_16 = pipe2_io_pipe_phv_out_data_16; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_17 = pipe2_io_pipe_phv_out_data_17; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_18 = pipe2_io_pipe_phv_out_data_18; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_19 = pipe2_io_pipe_phv_out_data_19; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_20 = pipe2_io_pipe_phv_out_data_20; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_21 = pipe2_io_pipe_phv_out_data_21; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_22 = pipe2_io_pipe_phv_out_data_22; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_23 = pipe2_io_pipe_phv_out_data_23; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_24 = pipe2_io_pipe_phv_out_data_24; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_25 = pipe2_io_pipe_phv_out_data_25; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_26 = pipe2_io_pipe_phv_out_data_26; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_27 = pipe2_io_pipe_phv_out_data_27; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_28 = pipe2_io_pipe_phv_out_data_28; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_29 = pipe2_io_pipe_phv_out_data_29; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_30 = pipe2_io_pipe_phv_out_data_30; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_31 = pipe2_io_pipe_phv_out_data_31; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_32 = pipe2_io_pipe_phv_out_data_32; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_33 = pipe2_io_pipe_phv_out_data_33; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_34 = pipe2_io_pipe_phv_out_data_34; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_35 = pipe2_io_pipe_phv_out_data_35; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_36 = pipe2_io_pipe_phv_out_data_36; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_37 = pipe2_io_pipe_phv_out_data_37; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_38 = pipe2_io_pipe_phv_out_data_38; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_39 = pipe2_io_pipe_phv_out_data_39; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_40 = pipe2_io_pipe_phv_out_data_40; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_41 = pipe2_io_pipe_phv_out_data_41; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_42 = pipe2_io_pipe_phv_out_data_42; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_43 = pipe2_io_pipe_phv_out_data_43; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_44 = pipe2_io_pipe_phv_out_data_44; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_45 = pipe2_io_pipe_phv_out_data_45; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_46 = pipe2_io_pipe_phv_out_data_46; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_47 = pipe2_io_pipe_phv_out_data_47; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_48 = pipe2_io_pipe_phv_out_data_48; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_49 = pipe2_io_pipe_phv_out_data_49; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_50 = pipe2_io_pipe_phv_out_data_50; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_51 = pipe2_io_pipe_phv_out_data_51; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_52 = pipe2_io_pipe_phv_out_data_52; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_53 = pipe2_io_pipe_phv_out_data_53; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_54 = pipe2_io_pipe_phv_out_data_54; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_55 = pipe2_io_pipe_phv_out_data_55; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_56 = pipe2_io_pipe_phv_out_data_56; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_57 = pipe2_io_pipe_phv_out_data_57; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_58 = pipe2_io_pipe_phv_out_data_58; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_59 = pipe2_io_pipe_phv_out_data_59; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_60 = pipe2_io_pipe_phv_out_data_60; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_61 = pipe2_io_pipe_phv_out_data_61; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_62 = pipe2_io_pipe_phv_out_data_62; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_63 = pipe2_io_pipe_phv_out_data_63; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_64 = pipe2_io_pipe_phv_out_data_64; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_65 = pipe2_io_pipe_phv_out_data_65; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_66 = pipe2_io_pipe_phv_out_data_66; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_67 = pipe2_io_pipe_phv_out_data_67; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_68 = pipe2_io_pipe_phv_out_data_68; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_69 = pipe2_io_pipe_phv_out_data_69; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_70 = pipe2_io_pipe_phv_out_data_70; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_71 = pipe2_io_pipe_phv_out_data_71; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_72 = pipe2_io_pipe_phv_out_data_72; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_73 = pipe2_io_pipe_phv_out_data_73; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_74 = pipe2_io_pipe_phv_out_data_74; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_75 = pipe2_io_pipe_phv_out_data_75; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_76 = pipe2_io_pipe_phv_out_data_76; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_77 = pipe2_io_pipe_phv_out_data_77; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_78 = pipe2_io_pipe_phv_out_data_78; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_79 = pipe2_io_pipe_phv_out_data_79; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_80 = pipe2_io_pipe_phv_out_data_80; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_81 = pipe2_io_pipe_phv_out_data_81; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_82 = pipe2_io_pipe_phv_out_data_82; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_83 = pipe2_io_pipe_phv_out_data_83; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_84 = pipe2_io_pipe_phv_out_data_84; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_85 = pipe2_io_pipe_phv_out_data_85; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_86 = pipe2_io_pipe_phv_out_data_86; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_87 = pipe2_io_pipe_phv_out_data_87; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_88 = pipe2_io_pipe_phv_out_data_88; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_89 = pipe2_io_pipe_phv_out_data_89; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_90 = pipe2_io_pipe_phv_out_data_90; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_91 = pipe2_io_pipe_phv_out_data_91; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_92 = pipe2_io_pipe_phv_out_data_92; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_93 = pipe2_io_pipe_phv_out_data_93; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_94 = pipe2_io_pipe_phv_out_data_94; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_data_95 = pipe2_io_pipe_phv_out_data_95; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_header_0 = pipe2_io_pipe_phv_out_header_0; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_header_1 = pipe2_io_pipe_phv_out_header_1; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_header_2 = pipe2_io_pipe_phv_out_header_2; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_header_3 = pipe2_io_pipe_phv_out_header_3; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_header_4 = pipe2_io_pipe_phv_out_header_4; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_header_5 = pipe2_io_pipe_phv_out_header_5; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_header_6 = pipe2_io_pipe_phv_out_header_6; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_header_7 = pipe2_io_pipe_phv_out_header_7; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_header_8 = pipe2_io_pipe_phv_out_header_8; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_header_9 = pipe2_io_pipe_phv_out_header_9; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_header_10 = pipe2_io_pipe_phv_out_header_10; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_header_11 = pipe2_io_pipe_phv_out_header_11; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_header_12 = pipe2_io_pipe_phv_out_header_12; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_header_13 = pipe2_io_pipe_phv_out_header_13; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_header_14 = pipe2_io_pipe_phv_out_header_14; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_header_15 = pipe2_io_pipe_phv_out_header_15; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_parse_current_state = pipe2_io_pipe_phv_out_parse_current_state; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_parse_current_offset = pipe2_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_parse_transition_field = pipe2_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_next_processor_id = pipe2_io_pipe_phv_out_next_processor_id; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_next_config_id = pipe2_io_pipe_phv_out_next_config_id; // @[matcher.scala 279:29]
  assign pipe3to8_io_pipe_phv_in_is_valid_processor = pipe2_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 279:29]
  assign pipe3to8_io_mod_hash_depth_mod = io_mod_en; // @[matcher.scala 280:36]
  assign pipe3to8_io_mod_config_id = io_mod_config_id; // @[matcher.scala 281:36]
  assign pipe3to8_io_mod_hash_depth = io_mod_table_mod_table_depth[2:0]; // @[matcher.scala 282:36]
  assign pipe3to8_io_key_in = pipe2_io_match_key; // @[matcher.scala 283:26]
  assign pipe9_clock = clock;
  assign pipe9_io_pipe_phv_in_data_0 = pipe3to8_io_pipe_phv_out_data_0; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_1 = pipe3to8_io_pipe_phv_out_data_1; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_2 = pipe3to8_io_pipe_phv_out_data_2; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_3 = pipe3to8_io_pipe_phv_out_data_3; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_4 = pipe3to8_io_pipe_phv_out_data_4; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_5 = pipe3to8_io_pipe_phv_out_data_5; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_6 = pipe3to8_io_pipe_phv_out_data_6; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_7 = pipe3to8_io_pipe_phv_out_data_7; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_8 = pipe3to8_io_pipe_phv_out_data_8; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_9 = pipe3to8_io_pipe_phv_out_data_9; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_10 = pipe3to8_io_pipe_phv_out_data_10; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_11 = pipe3to8_io_pipe_phv_out_data_11; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_12 = pipe3to8_io_pipe_phv_out_data_12; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_13 = pipe3to8_io_pipe_phv_out_data_13; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_14 = pipe3to8_io_pipe_phv_out_data_14; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_15 = pipe3to8_io_pipe_phv_out_data_15; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_16 = pipe3to8_io_pipe_phv_out_data_16; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_17 = pipe3to8_io_pipe_phv_out_data_17; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_18 = pipe3to8_io_pipe_phv_out_data_18; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_19 = pipe3to8_io_pipe_phv_out_data_19; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_20 = pipe3to8_io_pipe_phv_out_data_20; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_21 = pipe3to8_io_pipe_phv_out_data_21; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_22 = pipe3to8_io_pipe_phv_out_data_22; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_23 = pipe3to8_io_pipe_phv_out_data_23; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_24 = pipe3to8_io_pipe_phv_out_data_24; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_25 = pipe3to8_io_pipe_phv_out_data_25; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_26 = pipe3to8_io_pipe_phv_out_data_26; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_27 = pipe3to8_io_pipe_phv_out_data_27; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_28 = pipe3to8_io_pipe_phv_out_data_28; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_29 = pipe3to8_io_pipe_phv_out_data_29; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_30 = pipe3to8_io_pipe_phv_out_data_30; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_31 = pipe3to8_io_pipe_phv_out_data_31; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_32 = pipe3to8_io_pipe_phv_out_data_32; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_33 = pipe3to8_io_pipe_phv_out_data_33; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_34 = pipe3to8_io_pipe_phv_out_data_34; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_35 = pipe3to8_io_pipe_phv_out_data_35; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_36 = pipe3to8_io_pipe_phv_out_data_36; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_37 = pipe3to8_io_pipe_phv_out_data_37; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_38 = pipe3to8_io_pipe_phv_out_data_38; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_39 = pipe3to8_io_pipe_phv_out_data_39; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_40 = pipe3to8_io_pipe_phv_out_data_40; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_41 = pipe3to8_io_pipe_phv_out_data_41; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_42 = pipe3to8_io_pipe_phv_out_data_42; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_43 = pipe3to8_io_pipe_phv_out_data_43; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_44 = pipe3to8_io_pipe_phv_out_data_44; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_45 = pipe3to8_io_pipe_phv_out_data_45; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_46 = pipe3to8_io_pipe_phv_out_data_46; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_47 = pipe3to8_io_pipe_phv_out_data_47; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_48 = pipe3to8_io_pipe_phv_out_data_48; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_49 = pipe3to8_io_pipe_phv_out_data_49; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_50 = pipe3to8_io_pipe_phv_out_data_50; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_51 = pipe3to8_io_pipe_phv_out_data_51; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_52 = pipe3to8_io_pipe_phv_out_data_52; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_53 = pipe3to8_io_pipe_phv_out_data_53; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_54 = pipe3to8_io_pipe_phv_out_data_54; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_55 = pipe3to8_io_pipe_phv_out_data_55; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_56 = pipe3to8_io_pipe_phv_out_data_56; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_57 = pipe3to8_io_pipe_phv_out_data_57; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_58 = pipe3to8_io_pipe_phv_out_data_58; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_59 = pipe3to8_io_pipe_phv_out_data_59; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_60 = pipe3to8_io_pipe_phv_out_data_60; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_61 = pipe3to8_io_pipe_phv_out_data_61; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_62 = pipe3to8_io_pipe_phv_out_data_62; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_63 = pipe3to8_io_pipe_phv_out_data_63; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_64 = pipe3to8_io_pipe_phv_out_data_64; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_65 = pipe3to8_io_pipe_phv_out_data_65; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_66 = pipe3to8_io_pipe_phv_out_data_66; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_67 = pipe3to8_io_pipe_phv_out_data_67; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_68 = pipe3to8_io_pipe_phv_out_data_68; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_69 = pipe3to8_io_pipe_phv_out_data_69; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_70 = pipe3to8_io_pipe_phv_out_data_70; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_71 = pipe3to8_io_pipe_phv_out_data_71; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_72 = pipe3to8_io_pipe_phv_out_data_72; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_73 = pipe3to8_io_pipe_phv_out_data_73; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_74 = pipe3to8_io_pipe_phv_out_data_74; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_75 = pipe3to8_io_pipe_phv_out_data_75; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_76 = pipe3to8_io_pipe_phv_out_data_76; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_77 = pipe3to8_io_pipe_phv_out_data_77; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_78 = pipe3to8_io_pipe_phv_out_data_78; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_79 = pipe3to8_io_pipe_phv_out_data_79; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_80 = pipe3to8_io_pipe_phv_out_data_80; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_81 = pipe3to8_io_pipe_phv_out_data_81; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_82 = pipe3to8_io_pipe_phv_out_data_82; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_83 = pipe3to8_io_pipe_phv_out_data_83; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_84 = pipe3to8_io_pipe_phv_out_data_84; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_85 = pipe3to8_io_pipe_phv_out_data_85; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_86 = pipe3to8_io_pipe_phv_out_data_86; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_87 = pipe3to8_io_pipe_phv_out_data_87; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_88 = pipe3to8_io_pipe_phv_out_data_88; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_89 = pipe3to8_io_pipe_phv_out_data_89; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_90 = pipe3to8_io_pipe_phv_out_data_90; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_91 = pipe3to8_io_pipe_phv_out_data_91; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_92 = pipe3to8_io_pipe_phv_out_data_92; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_93 = pipe3to8_io_pipe_phv_out_data_93; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_94 = pipe3to8_io_pipe_phv_out_data_94; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_data_95 = pipe3to8_io_pipe_phv_out_data_95; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_header_0 = pipe3to8_io_pipe_phv_out_header_0; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_header_1 = pipe3to8_io_pipe_phv_out_header_1; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_header_2 = pipe3to8_io_pipe_phv_out_header_2; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_header_3 = pipe3to8_io_pipe_phv_out_header_3; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_header_4 = pipe3to8_io_pipe_phv_out_header_4; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_header_5 = pipe3to8_io_pipe_phv_out_header_5; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_header_6 = pipe3to8_io_pipe_phv_out_header_6; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_header_7 = pipe3to8_io_pipe_phv_out_header_7; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_header_8 = pipe3to8_io_pipe_phv_out_header_8; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_header_9 = pipe3to8_io_pipe_phv_out_header_9; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_header_10 = pipe3to8_io_pipe_phv_out_header_10; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_header_11 = pipe3to8_io_pipe_phv_out_header_11; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_header_12 = pipe3to8_io_pipe_phv_out_header_12; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_header_13 = pipe3to8_io_pipe_phv_out_header_13; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_header_14 = pipe3to8_io_pipe_phv_out_header_14; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_header_15 = pipe3to8_io_pipe_phv_out_header_15; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_parse_current_state = pipe3to8_io_pipe_phv_out_parse_current_state; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_parse_current_offset = pipe3to8_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_parse_transition_field = pipe3to8_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_next_processor_id = pipe3to8_io_pipe_phv_out_next_processor_id; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_next_config_id = pipe3to8_io_pipe_phv_out_next_config_id; // @[matcher.scala 285:27]
  assign pipe9_io_pipe_phv_in_is_valid_processor = pipe3to8_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 285:27]
  assign pipe9_io_table_config_0_table_width = table_config_0_table_width; // @[matcher.scala 289:27]
  assign pipe9_io_table_config_0_table_depth = table_config_0_table_depth; // @[matcher.scala 289:27]
  assign pipe9_io_table_config_1_table_width = table_config_1_table_width; // @[matcher.scala 289:27]
  assign pipe9_io_table_config_1_table_depth = table_config_1_table_depth; // @[matcher.scala 289:27]
  assign pipe9_io_key_in = pipe3to8_io_key_out; // @[matcher.scala 286:27]
  assign pipe9_io_addr_in = pipe3to8_io_hash_val; // @[matcher.scala 287:27]
  assign pipe9_io_cs_in = pipe3to8_io_hash_val_cs; // @[matcher.scala 288:27]
  assign pipe10_clock = clock;
  assign pipe10_io_pipe_phv_in_data_0 = pipe9_io_pipe_phv_out_data_0; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_1 = pipe9_io_pipe_phv_out_data_1; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_2 = pipe9_io_pipe_phv_out_data_2; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_3 = pipe9_io_pipe_phv_out_data_3; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_4 = pipe9_io_pipe_phv_out_data_4; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_5 = pipe9_io_pipe_phv_out_data_5; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_6 = pipe9_io_pipe_phv_out_data_6; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_7 = pipe9_io_pipe_phv_out_data_7; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_8 = pipe9_io_pipe_phv_out_data_8; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_9 = pipe9_io_pipe_phv_out_data_9; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_10 = pipe9_io_pipe_phv_out_data_10; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_11 = pipe9_io_pipe_phv_out_data_11; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_12 = pipe9_io_pipe_phv_out_data_12; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_13 = pipe9_io_pipe_phv_out_data_13; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_14 = pipe9_io_pipe_phv_out_data_14; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_15 = pipe9_io_pipe_phv_out_data_15; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_16 = pipe9_io_pipe_phv_out_data_16; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_17 = pipe9_io_pipe_phv_out_data_17; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_18 = pipe9_io_pipe_phv_out_data_18; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_19 = pipe9_io_pipe_phv_out_data_19; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_20 = pipe9_io_pipe_phv_out_data_20; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_21 = pipe9_io_pipe_phv_out_data_21; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_22 = pipe9_io_pipe_phv_out_data_22; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_23 = pipe9_io_pipe_phv_out_data_23; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_24 = pipe9_io_pipe_phv_out_data_24; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_25 = pipe9_io_pipe_phv_out_data_25; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_26 = pipe9_io_pipe_phv_out_data_26; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_27 = pipe9_io_pipe_phv_out_data_27; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_28 = pipe9_io_pipe_phv_out_data_28; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_29 = pipe9_io_pipe_phv_out_data_29; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_30 = pipe9_io_pipe_phv_out_data_30; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_31 = pipe9_io_pipe_phv_out_data_31; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_32 = pipe9_io_pipe_phv_out_data_32; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_33 = pipe9_io_pipe_phv_out_data_33; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_34 = pipe9_io_pipe_phv_out_data_34; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_35 = pipe9_io_pipe_phv_out_data_35; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_36 = pipe9_io_pipe_phv_out_data_36; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_37 = pipe9_io_pipe_phv_out_data_37; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_38 = pipe9_io_pipe_phv_out_data_38; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_39 = pipe9_io_pipe_phv_out_data_39; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_40 = pipe9_io_pipe_phv_out_data_40; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_41 = pipe9_io_pipe_phv_out_data_41; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_42 = pipe9_io_pipe_phv_out_data_42; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_43 = pipe9_io_pipe_phv_out_data_43; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_44 = pipe9_io_pipe_phv_out_data_44; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_45 = pipe9_io_pipe_phv_out_data_45; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_46 = pipe9_io_pipe_phv_out_data_46; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_47 = pipe9_io_pipe_phv_out_data_47; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_48 = pipe9_io_pipe_phv_out_data_48; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_49 = pipe9_io_pipe_phv_out_data_49; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_50 = pipe9_io_pipe_phv_out_data_50; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_51 = pipe9_io_pipe_phv_out_data_51; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_52 = pipe9_io_pipe_phv_out_data_52; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_53 = pipe9_io_pipe_phv_out_data_53; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_54 = pipe9_io_pipe_phv_out_data_54; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_55 = pipe9_io_pipe_phv_out_data_55; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_56 = pipe9_io_pipe_phv_out_data_56; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_57 = pipe9_io_pipe_phv_out_data_57; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_58 = pipe9_io_pipe_phv_out_data_58; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_59 = pipe9_io_pipe_phv_out_data_59; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_60 = pipe9_io_pipe_phv_out_data_60; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_61 = pipe9_io_pipe_phv_out_data_61; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_62 = pipe9_io_pipe_phv_out_data_62; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_63 = pipe9_io_pipe_phv_out_data_63; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_64 = pipe9_io_pipe_phv_out_data_64; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_65 = pipe9_io_pipe_phv_out_data_65; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_66 = pipe9_io_pipe_phv_out_data_66; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_67 = pipe9_io_pipe_phv_out_data_67; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_68 = pipe9_io_pipe_phv_out_data_68; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_69 = pipe9_io_pipe_phv_out_data_69; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_70 = pipe9_io_pipe_phv_out_data_70; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_71 = pipe9_io_pipe_phv_out_data_71; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_72 = pipe9_io_pipe_phv_out_data_72; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_73 = pipe9_io_pipe_phv_out_data_73; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_74 = pipe9_io_pipe_phv_out_data_74; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_75 = pipe9_io_pipe_phv_out_data_75; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_76 = pipe9_io_pipe_phv_out_data_76; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_77 = pipe9_io_pipe_phv_out_data_77; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_78 = pipe9_io_pipe_phv_out_data_78; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_79 = pipe9_io_pipe_phv_out_data_79; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_80 = pipe9_io_pipe_phv_out_data_80; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_81 = pipe9_io_pipe_phv_out_data_81; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_82 = pipe9_io_pipe_phv_out_data_82; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_83 = pipe9_io_pipe_phv_out_data_83; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_84 = pipe9_io_pipe_phv_out_data_84; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_85 = pipe9_io_pipe_phv_out_data_85; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_86 = pipe9_io_pipe_phv_out_data_86; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_87 = pipe9_io_pipe_phv_out_data_87; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_88 = pipe9_io_pipe_phv_out_data_88; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_89 = pipe9_io_pipe_phv_out_data_89; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_90 = pipe9_io_pipe_phv_out_data_90; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_91 = pipe9_io_pipe_phv_out_data_91; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_92 = pipe9_io_pipe_phv_out_data_92; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_93 = pipe9_io_pipe_phv_out_data_93; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_94 = pipe9_io_pipe_phv_out_data_94; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_data_95 = pipe9_io_pipe_phv_out_data_95; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_header_0 = pipe9_io_pipe_phv_out_header_0; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_header_1 = pipe9_io_pipe_phv_out_header_1; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_header_2 = pipe9_io_pipe_phv_out_header_2; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_header_3 = pipe9_io_pipe_phv_out_header_3; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_header_4 = pipe9_io_pipe_phv_out_header_4; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_header_5 = pipe9_io_pipe_phv_out_header_5; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_header_6 = pipe9_io_pipe_phv_out_header_6; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_header_7 = pipe9_io_pipe_phv_out_header_7; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_header_8 = pipe9_io_pipe_phv_out_header_8; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_header_9 = pipe9_io_pipe_phv_out_header_9; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_header_10 = pipe9_io_pipe_phv_out_header_10; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_header_11 = pipe9_io_pipe_phv_out_header_11; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_header_12 = pipe9_io_pipe_phv_out_header_12; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_header_13 = pipe9_io_pipe_phv_out_header_13; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_header_14 = pipe9_io_pipe_phv_out_header_14; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_header_15 = pipe9_io_pipe_phv_out_header_15; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_parse_current_state = pipe9_io_pipe_phv_out_parse_current_state; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_parse_current_offset = pipe9_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_parse_transition_field = pipe9_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_next_processor_id = pipe9_io_pipe_phv_out_next_processor_id; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_next_config_id = pipe9_io_pipe_phv_out_next_config_id; // @[matcher.scala 291:27]
  assign pipe10_io_pipe_phv_in_is_valid_processor = pipe9_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 291:27]
  assign pipe10_io_key_in = pipe9_io_key_out; // @[matcher.scala 292:27]
  assign pipe10_io_cs_in = pipe9_io_cs_out; // @[matcher.scala 293:27]
  assign pipe10_io_addr_in = pipe9_io_addr_out; // @[matcher.scala 294:27]
  assign pipe10_io_cs_vec_in_0 = pipe9_io_cs_vec_out_0; // @[matcher.scala 295:27]
  assign pipe10_io_cs_vec_in_1 = pipe9_io_cs_vec_out_1; // @[matcher.scala 295:27]
  assign pipe10_io_cs_vec_in_2 = pipe9_io_cs_vec_out_2; // @[matcher.scala 295:27]
  assign pipe10_io_cs_vec_in_3 = pipe9_io_cs_vec_out_3; // @[matcher.scala 295:27]
  assign pipe10_io_cs_vec_in_4 = pipe9_io_cs_vec_out_4; // @[matcher.scala 295:27]
  assign pipe10_io_cs_vec_in_5 = pipe9_io_cs_vec_out_5; // @[matcher.scala 295:27]
  assign pipe10_io_cs_vec_in_6 = pipe9_io_cs_vec_out_6; // @[matcher.scala 295:27]
  assign pipe10_io_cs_vec_in_7 = pipe9_io_cs_vec_out_7; // @[matcher.scala 295:27]
  assign pipe10_io_mem_cluster_0_data = io_mem_cluster_0_data; // @[matcher.scala 296:27]
  assign pipe10_io_mem_cluster_1_data = io_mem_cluster_1_data; // @[matcher.scala 296:27]
  assign pipe10_io_mem_cluster_2_data = io_mem_cluster_2_data; // @[matcher.scala 296:27]
  assign pipe10_io_mem_cluster_3_data = io_mem_cluster_3_data; // @[matcher.scala 296:27]
  assign pipe10_io_mem_cluster_4_data = io_mem_cluster_4_data; // @[matcher.scala 296:27]
  assign pipe10_io_mem_cluster_5_data = io_mem_cluster_5_data; // @[matcher.scala 296:27]
  assign pipe10_io_mem_cluster_6_data = io_mem_cluster_6_data; // @[matcher.scala 296:27]
  assign pipe10_io_mem_cluster_7_data = io_mem_cluster_7_data; // @[matcher.scala 296:27]
  assign pipe11_clock = clock;
  assign pipe11_io_pipe_phv_in_data_0 = pipe10_io_pipe_phv_out_data_0; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_1 = pipe10_io_pipe_phv_out_data_1; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_2 = pipe10_io_pipe_phv_out_data_2; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_3 = pipe10_io_pipe_phv_out_data_3; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_4 = pipe10_io_pipe_phv_out_data_4; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_5 = pipe10_io_pipe_phv_out_data_5; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_6 = pipe10_io_pipe_phv_out_data_6; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_7 = pipe10_io_pipe_phv_out_data_7; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_8 = pipe10_io_pipe_phv_out_data_8; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_9 = pipe10_io_pipe_phv_out_data_9; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_10 = pipe10_io_pipe_phv_out_data_10; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_11 = pipe10_io_pipe_phv_out_data_11; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_12 = pipe10_io_pipe_phv_out_data_12; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_13 = pipe10_io_pipe_phv_out_data_13; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_14 = pipe10_io_pipe_phv_out_data_14; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_15 = pipe10_io_pipe_phv_out_data_15; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_16 = pipe10_io_pipe_phv_out_data_16; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_17 = pipe10_io_pipe_phv_out_data_17; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_18 = pipe10_io_pipe_phv_out_data_18; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_19 = pipe10_io_pipe_phv_out_data_19; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_20 = pipe10_io_pipe_phv_out_data_20; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_21 = pipe10_io_pipe_phv_out_data_21; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_22 = pipe10_io_pipe_phv_out_data_22; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_23 = pipe10_io_pipe_phv_out_data_23; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_24 = pipe10_io_pipe_phv_out_data_24; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_25 = pipe10_io_pipe_phv_out_data_25; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_26 = pipe10_io_pipe_phv_out_data_26; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_27 = pipe10_io_pipe_phv_out_data_27; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_28 = pipe10_io_pipe_phv_out_data_28; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_29 = pipe10_io_pipe_phv_out_data_29; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_30 = pipe10_io_pipe_phv_out_data_30; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_31 = pipe10_io_pipe_phv_out_data_31; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_32 = pipe10_io_pipe_phv_out_data_32; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_33 = pipe10_io_pipe_phv_out_data_33; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_34 = pipe10_io_pipe_phv_out_data_34; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_35 = pipe10_io_pipe_phv_out_data_35; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_36 = pipe10_io_pipe_phv_out_data_36; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_37 = pipe10_io_pipe_phv_out_data_37; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_38 = pipe10_io_pipe_phv_out_data_38; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_39 = pipe10_io_pipe_phv_out_data_39; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_40 = pipe10_io_pipe_phv_out_data_40; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_41 = pipe10_io_pipe_phv_out_data_41; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_42 = pipe10_io_pipe_phv_out_data_42; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_43 = pipe10_io_pipe_phv_out_data_43; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_44 = pipe10_io_pipe_phv_out_data_44; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_45 = pipe10_io_pipe_phv_out_data_45; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_46 = pipe10_io_pipe_phv_out_data_46; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_47 = pipe10_io_pipe_phv_out_data_47; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_48 = pipe10_io_pipe_phv_out_data_48; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_49 = pipe10_io_pipe_phv_out_data_49; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_50 = pipe10_io_pipe_phv_out_data_50; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_51 = pipe10_io_pipe_phv_out_data_51; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_52 = pipe10_io_pipe_phv_out_data_52; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_53 = pipe10_io_pipe_phv_out_data_53; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_54 = pipe10_io_pipe_phv_out_data_54; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_55 = pipe10_io_pipe_phv_out_data_55; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_56 = pipe10_io_pipe_phv_out_data_56; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_57 = pipe10_io_pipe_phv_out_data_57; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_58 = pipe10_io_pipe_phv_out_data_58; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_59 = pipe10_io_pipe_phv_out_data_59; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_60 = pipe10_io_pipe_phv_out_data_60; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_61 = pipe10_io_pipe_phv_out_data_61; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_62 = pipe10_io_pipe_phv_out_data_62; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_63 = pipe10_io_pipe_phv_out_data_63; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_64 = pipe10_io_pipe_phv_out_data_64; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_65 = pipe10_io_pipe_phv_out_data_65; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_66 = pipe10_io_pipe_phv_out_data_66; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_67 = pipe10_io_pipe_phv_out_data_67; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_68 = pipe10_io_pipe_phv_out_data_68; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_69 = pipe10_io_pipe_phv_out_data_69; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_70 = pipe10_io_pipe_phv_out_data_70; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_71 = pipe10_io_pipe_phv_out_data_71; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_72 = pipe10_io_pipe_phv_out_data_72; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_73 = pipe10_io_pipe_phv_out_data_73; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_74 = pipe10_io_pipe_phv_out_data_74; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_75 = pipe10_io_pipe_phv_out_data_75; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_76 = pipe10_io_pipe_phv_out_data_76; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_77 = pipe10_io_pipe_phv_out_data_77; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_78 = pipe10_io_pipe_phv_out_data_78; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_79 = pipe10_io_pipe_phv_out_data_79; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_80 = pipe10_io_pipe_phv_out_data_80; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_81 = pipe10_io_pipe_phv_out_data_81; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_82 = pipe10_io_pipe_phv_out_data_82; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_83 = pipe10_io_pipe_phv_out_data_83; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_84 = pipe10_io_pipe_phv_out_data_84; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_85 = pipe10_io_pipe_phv_out_data_85; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_86 = pipe10_io_pipe_phv_out_data_86; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_87 = pipe10_io_pipe_phv_out_data_87; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_88 = pipe10_io_pipe_phv_out_data_88; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_89 = pipe10_io_pipe_phv_out_data_89; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_90 = pipe10_io_pipe_phv_out_data_90; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_91 = pipe10_io_pipe_phv_out_data_91; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_92 = pipe10_io_pipe_phv_out_data_92; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_93 = pipe10_io_pipe_phv_out_data_93; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_94 = pipe10_io_pipe_phv_out_data_94; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_data_95 = pipe10_io_pipe_phv_out_data_95; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_header_0 = pipe10_io_pipe_phv_out_header_0; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_header_1 = pipe10_io_pipe_phv_out_header_1; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_header_2 = pipe10_io_pipe_phv_out_header_2; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_header_3 = pipe10_io_pipe_phv_out_header_3; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_header_4 = pipe10_io_pipe_phv_out_header_4; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_header_5 = pipe10_io_pipe_phv_out_header_5; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_header_6 = pipe10_io_pipe_phv_out_header_6; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_header_7 = pipe10_io_pipe_phv_out_header_7; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_header_8 = pipe10_io_pipe_phv_out_header_8; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_header_9 = pipe10_io_pipe_phv_out_header_9; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_header_10 = pipe10_io_pipe_phv_out_header_10; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_header_11 = pipe10_io_pipe_phv_out_header_11; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_header_12 = pipe10_io_pipe_phv_out_header_12; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_header_13 = pipe10_io_pipe_phv_out_header_13; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_header_14 = pipe10_io_pipe_phv_out_header_14; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_header_15 = pipe10_io_pipe_phv_out_header_15; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_parse_current_state = pipe10_io_pipe_phv_out_parse_current_state; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_parse_current_offset = pipe10_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_parse_transition_field = pipe10_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_next_processor_id = pipe10_io_pipe_phv_out_next_processor_id; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_next_config_id = pipe10_io_pipe_phv_out_next_config_id; // @[matcher.scala 298:27]
  assign pipe11_io_pipe_phv_in_is_valid_processor = pipe10_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 298:27]
  assign pipe11_io_table_config_0_table_width = table_config_0_table_width; // @[matcher.scala 302:28]
  assign pipe11_io_table_config_0_table_depth = table_config_0_table_depth; // @[matcher.scala 302:28]
  assign pipe11_io_table_config_1_table_width = table_config_1_table_width; // @[matcher.scala 302:28]
  assign pipe11_io_table_config_1_table_depth = table_config_1_table_depth; // @[matcher.scala 302:28]
  assign pipe11_io_key_in = pipe10_io_key_out; // @[matcher.scala 299:27]
  assign pipe11_io_cs_in = pipe10_io_cs_out; // @[matcher.scala 300:27]
  assign pipe11_io_data_in_0 = pipe10_io_data_out_0; // @[matcher.scala 301:27]
  assign pipe11_io_data_in_1 = pipe10_io_data_out_1; // @[matcher.scala 301:27]
  assign pipe11_io_data_in_2 = pipe10_io_data_out_2; // @[matcher.scala 301:27]
  assign pipe11_io_data_in_3 = pipe10_io_data_out_3; // @[matcher.scala 301:27]
  assign pipe11_io_data_in_4 = pipe10_io_data_out_4; // @[matcher.scala 301:27]
  assign pipe11_io_data_in_5 = pipe10_io_data_out_5; // @[matcher.scala 301:27]
  assign pipe11_io_data_in_6 = pipe10_io_data_out_6; // @[matcher.scala 301:27]
  assign pipe11_io_data_in_7 = pipe10_io_data_out_7; // @[matcher.scala 301:27]
  assign pipe12_clock = clock;
  assign pipe12_io_pipe_phv_in_data_0 = pipe11_io_pipe_phv_out_data_0; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_1 = pipe11_io_pipe_phv_out_data_1; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_2 = pipe11_io_pipe_phv_out_data_2; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_3 = pipe11_io_pipe_phv_out_data_3; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_4 = pipe11_io_pipe_phv_out_data_4; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_5 = pipe11_io_pipe_phv_out_data_5; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_6 = pipe11_io_pipe_phv_out_data_6; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_7 = pipe11_io_pipe_phv_out_data_7; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_8 = pipe11_io_pipe_phv_out_data_8; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_9 = pipe11_io_pipe_phv_out_data_9; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_10 = pipe11_io_pipe_phv_out_data_10; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_11 = pipe11_io_pipe_phv_out_data_11; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_12 = pipe11_io_pipe_phv_out_data_12; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_13 = pipe11_io_pipe_phv_out_data_13; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_14 = pipe11_io_pipe_phv_out_data_14; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_15 = pipe11_io_pipe_phv_out_data_15; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_16 = pipe11_io_pipe_phv_out_data_16; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_17 = pipe11_io_pipe_phv_out_data_17; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_18 = pipe11_io_pipe_phv_out_data_18; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_19 = pipe11_io_pipe_phv_out_data_19; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_20 = pipe11_io_pipe_phv_out_data_20; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_21 = pipe11_io_pipe_phv_out_data_21; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_22 = pipe11_io_pipe_phv_out_data_22; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_23 = pipe11_io_pipe_phv_out_data_23; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_24 = pipe11_io_pipe_phv_out_data_24; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_25 = pipe11_io_pipe_phv_out_data_25; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_26 = pipe11_io_pipe_phv_out_data_26; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_27 = pipe11_io_pipe_phv_out_data_27; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_28 = pipe11_io_pipe_phv_out_data_28; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_29 = pipe11_io_pipe_phv_out_data_29; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_30 = pipe11_io_pipe_phv_out_data_30; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_31 = pipe11_io_pipe_phv_out_data_31; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_32 = pipe11_io_pipe_phv_out_data_32; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_33 = pipe11_io_pipe_phv_out_data_33; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_34 = pipe11_io_pipe_phv_out_data_34; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_35 = pipe11_io_pipe_phv_out_data_35; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_36 = pipe11_io_pipe_phv_out_data_36; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_37 = pipe11_io_pipe_phv_out_data_37; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_38 = pipe11_io_pipe_phv_out_data_38; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_39 = pipe11_io_pipe_phv_out_data_39; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_40 = pipe11_io_pipe_phv_out_data_40; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_41 = pipe11_io_pipe_phv_out_data_41; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_42 = pipe11_io_pipe_phv_out_data_42; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_43 = pipe11_io_pipe_phv_out_data_43; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_44 = pipe11_io_pipe_phv_out_data_44; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_45 = pipe11_io_pipe_phv_out_data_45; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_46 = pipe11_io_pipe_phv_out_data_46; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_47 = pipe11_io_pipe_phv_out_data_47; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_48 = pipe11_io_pipe_phv_out_data_48; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_49 = pipe11_io_pipe_phv_out_data_49; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_50 = pipe11_io_pipe_phv_out_data_50; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_51 = pipe11_io_pipe_phv_out_data_51; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_52 = pipe11_io_pipe_phv_out_data_52; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_53 = pipe11_io_pipe_phv_out_data_53; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_54 = pipe11_io_pipe_phv_out_data_54; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_55 = pipe11_io_pipe_phv_out_data_55; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_56 = pipe11_io_pipe_phv_out_data_56; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_57 = pipe11_io_pipe_phv_out_data_57; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_58 = pipe11_io_pipe_phv_out_data_58; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_59 = pipe11_io_pipe_phv_out_data_59; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_60 = pipe11_io_pipe_phv_out_data_60; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_61 = pipe11_io_pipe_phv_out_data_61; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_62 = pipe11_io_pipe_phv_out_data_62; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_63 = pipe11_io_pipe_phv_out_data_63; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_64 = pipe11_io_pipe_phv_out_data_64; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_65 = pipe11_io_pipe_phv_out_data_65; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_66 = pipe11_io_pipe_phv_out_data_66; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_67 = pipe11_io_pipe_phv_out_data_67; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_68 = pipe11_io_pipe_phv_out_data_68; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_69 = pipe11_io_pipe_phv_out_data_69; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_70 = pipe11_io_pipe_phv_out_data_70; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_71 = pipe11_io_pipe_phv_out_data_71; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_72 = pipe11_io_pipe_phv_out_data_72; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_73 = pipe11_io_pipe_phv_out_data_73; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_74 = pipe11_io_pipe_phv_out_data_74; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_75 = pipe11_io_pipe_phv_out_data_75; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_76 = pipe11_io_pipe_phv_out_data_76; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_77 = pipe11_io_pipe_phv_out_data_77; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_78 = pipe11_io_pipe_phv_out_data_78; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_79 = pipe11_io_pipe_phv_out_data_79; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_80 = pipe11_io_pipe_phv_out_data_80; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_81 = pipe11_io_pipe_phv_out_data_81; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_82 = pipe11_io_pipe_phv_out_data_82; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_83 = pipe11_io_pipe_phv_out_data_83; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_84 = pipe11_io_pipe_phv_out_data_84; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_85 = pipe11_io_pipe_phv_out_data_85; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_86 = pipe11_io_pipe_phv_out_data_86; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_87 = pipe11_io_pipe_phv_out_data_87; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_88 = pipe11_io_pipe_phv_out_data_88; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_89 = pipe11_io_pipe_phv_out_data_89; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_90 = pipe11_io_pipe_phv_out_data_90; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_91 = pipe11_io_pipe_phv_out_data_91; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_92 = pipe11_io_pipe_phv_out_data_92; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_93 = pipe11_io_pipe_phv_out_data_93; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_94 = pipe11_io_pipe_phv_out_data_94; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_data_95 = pipe11_io_pipe_phv_out_data_95; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_header_0 = pipe11_io_pipe_phv_out_header_0; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_header_1 = pipe11_io_pipe_phv_out_header_1; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_header_2 = pipe11_io_pipe_phv_out_header_2; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_header_3 = pipe11_io_pipe_phv_out_header_3; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_header_4 = pipe11_io_pipe_phv_out_header_4; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_header_5 = pipe11_io_pipe_phv_out_header_5; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_header_6 = pipe11_io_pipe_phv_out_header_6; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_header_7 = pipe11_io_pipe_phv_out_header_7; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_header_8 = pipe11_io_pipe_phv_out_header_8; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_header_9 = pipe11_io_pipe_phv_out_header_9; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_header_10 = pipe11_io_pipe_phv_out_header_10; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_header_11 = pipe11_io_pipe_phv_out_header_11; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_header_12 = pipe11_io_pipe_phv_out_header_12; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_header_13 = pipe11_io_pipe_phv_out_header_13; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_header_14 = pipe11_io_pipe_phv_out_header_14; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_header_15 = pipe11_io_pipe_phv_out_header_15; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_parse_current_state = pipe11_io_pipe_phv_out_parse_current_state; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_parse_current_offset = pipe11_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_parse_transition_field = pipe11_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_next_processor_id = pipe11_io_pipe_phv_out_next_processor_id; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_next_config_id = pipe11_io_pipe_phv_out_next_config_id; // @[matcher.scala 304:27]
  assign pipe12_io_pipe_phv_in_is_valid_processor = pipe11_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 304:27]
  assign pipe12_io_key_config_0_key_length = key_config_0_key_length; // @[matcher.scala 307:27]
  assign pipe12_io_key_config_1_key_length = key_config_1_key_length; // @[matcher.scala 307:27]
  assign pipe12_io_key_in = pipe11_io_key_out; // @[matcher.scala 305:27]
  assign pipe12_io_data_in = pipe11_io_data_out; // @[matcher.scala 306:27]
  always @(posedge clock) begin
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_0_header_id <= io_mod_key_mod_header_id; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_0_internal_offset <= io_mod_key_mod_internal_offset; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_0_key_length <= io_mod_key_mod_key_length; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_1_header_id <= io_mod_key_mod_header_id; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_1_internal_offset <= io_mod_key_mod_internal_offset; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_1_key_length <= io_mod_key_mod_key_length; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_table_width <= io_mod_table_mod_table_width; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_table_depth <= io_mod_table_mod_table_depth; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_table_width <= io_mod_table_mod_table_width; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_table_depth <= io_mod_table_mod_table_depth; // @[matcher.scala 22:40]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  key_config_0_header_id = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  key_config_0_internal_offset = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  key_config_0_key_length = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  key_config_1_header_id = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  key_config_1_internal_offset = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  key_config_1_key_length = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  table_config_0_table_width = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  table_config_0_table_depth = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  table_config_1_table_width = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  table_config_1_table_depth = _RAND_9[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
