module IPSA(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  input         io_mod_proc_mod_0_par_mod_en,
  input         io_mod_proc_mod_0_par_mod_last_mau_id_mod,
  input  [1:0]  io_mod_proc_mod_0_par_mod_last_mau_id,
  input  [1:0]  io_mod_proc_mod_0_par_mod_cs,
  input         io_mod_proc_mod_0_par_mod_module_mod_state_id_mod,
  input  [7:0]  io_mod_proc_mod_0_par_mod_module_mod_state_id,
  input         io_mod_proc_mod_0_par_mod_module_mod_sram_w_cs,
  input         io_mod_proc_mod_0_par_mod_module_mod_sram_w_en,
  input  [7:0]  io_mod_proc_mod_0_par_mod_module_mod_sram_w_addr,
  input  [63:0] io_mod_proc_mod_0_par_mod_module_mod_sram_w_data,
  input         io_mod_proc_mod_0_mat_mod_en,
  input         io_mod_proc_mod_0_mat_mod_config_id,
  input  [7:0]  io_mod_proc_mod_0_mat_mod_key_mod_header_id,
  input  [7:0]  io_mod_proc_mod_0_mat_mod_key_mod_internal_offset,
  input  [7:0]  io_mod_proc_mod_0_mat_mod_key_mod_key_length,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_0,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_1,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_2,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_3,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_4,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_5,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_6,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_7,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_8,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_9,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_10,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_11,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_12,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_13,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_14,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_15,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_16,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_17,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_18,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_19,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_20,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_21,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_22,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_23,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_24,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_25,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_26,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_27,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_28,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_29,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_30,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_31,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_32,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_33,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_34,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_35,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_36,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_37,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_38,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_39,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_40,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_41,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_42,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_43,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_44,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_45,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_46,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_47,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_48,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_49,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_50,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_51,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_52,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_53,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_54,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_55,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_56,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_57,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_58,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_59,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_60,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_61,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_62,
  input  [5:0]  io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_63,
  input  [6:0]  io_mod_proc_mod_0_mat_mod_table_mod_table_width,
  input  [6:0]  io_mod_proc_mod_0_mat_mod_table_mod_table_depth,
  input         io_mod_proc_mod_0_act_mod_en_0,
  input         io_mod_proc_mod_0_act_mod_en_1,
  input  [7:0]  io_mod_proc_mod_0_act_mod_addr,
  input  [63:0] io_mod_proc_mod_0_act_mod_data_0,
  input  [63:0] io_mod_proc_mod_0_act_mod_data_1,
  input         io_mod_proc_mod_1_par_mod_en,
  input         io_mod_proc_mod_1_par_mod_last_mau_id_mod,
  input  [1:0]  io_mod_proc_mod_1_par_mod_last_mau_id,
  input  [1:0]  io_mod_proc_mod_1_par_mod_cs,
  input         io_mod_proc_mod_1_par_mod_module_mod_state_id_mod,
  input  [7:0]  io_mod_proc_mod_1_par_mod_module_mod_state_id,
  input         io_mod_proc_mod_1_par_mod_module_mod_sram_w_cs,
  input         io_mod_proc_mod_1_par_mod_module_mod_sram_w_en,
  input  [7:0]  io_mod_proc_mod_1_par_mod_module_mod_sram_w_addr,
  input  [63:0] io_mod_proc_mod_1_par_mod_module_mod_sram_w_data,
  input         io_mod_proc_mod_1_mat_mod_en,
  input         io_mod_proc_mod_1_mat_mod_config_id,
  input  [7:0]  io_mod_proc_mod_1_mat_mod_key_mod_header_id,
  input  [7:0]  io_mod_proc_mod_1_mat_mod_key_mod_internal_offset,
  input  [7:0]  io_mod_proc_mod_1_mat_mod_key_mod_key_length,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_0,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_1,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_2,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_3,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_4,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_5,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_6,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_7,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_8,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_9,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_10,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_11,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_12,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_13,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_14,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_15,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_16,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_17,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_18,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_19,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_20,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_21,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_22,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_23,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_24,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_25,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_26,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_27,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_28,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_29,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_30,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_31,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_32,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_33,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_34,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_35,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_36,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_37,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_38,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_39,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_40,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_41,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_42,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_43,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_44,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_45,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_46,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_47,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_48,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_49,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_50,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_51,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_52,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_53,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_54,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_55,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_56,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_57,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_58,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_59,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_60,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_61,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_62,
  input  [5:0]  io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_63,
  input  [6:0]  io_mod_proc_mod_1_mat_mod_table_mod_table_width,
  input  [6:0]  io_mod_proc_mod_1_mat_mod_table_mod_table_depth,
  input         io_mod_proc_mod_1_act_mod_en_0,
  input         io_mod_proc_mod_1_act_mod_en_1,
  input  [7:0]  io_mod_proc_mod_1_act_mod_addr,
  input  [63:0] io_mod_proc_mod_1_act_mod_data_0,
  input  [63:0] io_mod_proc_mod_1_act_mod_data_1,
  input         io_mod_proc_mod_2_par_mod_en,
  input         io_mod_proc_mod_2_par_mod_last_mau_id_mod,
  input  [1:0]  io_mod_proc_mod_2_par_mod_last_mau_id,
  input  [1:0]  io_mod_proc_mod_2_par_mod_cs,
  input         io_mod_proc_mod_2_par_mod_module_mod_state_id_mod,
  input  [7:0]  io_mod_proc_mod_2_par_mod_module_mod_state_id,
  input         io_mod_proc_mod_2_par_mod_module_mod_sram_w_cs,
  input         io_mod_proc_mod_2_par_mod_module_mod_sram_w_en,
  input  [7:0]  io_mod_proc_mod_2_par_mod_module_mod_sram_w_addr,
  input  [63:0] io_mod_proc_mod_2_par_mod_module_mod_sram_w_data,
  input         io_mod_proc_mod_2_mat_mod_en,
  input         io_mod_proc_mod_2_mat_mod_config_id,
  input  [7:0]  io_mod_proc_mod_2_mat_mod_key_mod_header_id,
  input  [7:0]  io_mod_proc_mod_2_mat_mod_key_mod_internal_offset,
  input  [7:0]  io_mod_proc_mod_2_mat_mod_key_mod_key_length,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_0,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_1,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_2,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_3,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_4,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_5,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_6,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_7,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_8,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_9,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_10,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_11,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_12,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_13,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_14,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_15,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_16,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_17,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_18,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_19,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_20,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_21,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_22,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_23,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_24,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_25,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_26,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_27,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_28,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_29,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_30,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_31,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_32,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_33,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_34,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_35,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_36,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_37,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_38,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_39,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_40,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_41,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_42,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_43,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_44,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_45,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_46,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_47,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_48,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_49,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_50,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_51,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_52,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_53,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_54,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_55,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_56,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_57,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_58,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_59,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_60,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_61,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_62,
  input  [5:0]  io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_63,
  input  [6:0]  io_mod_proc_mod_2_mat_mod_table_mod_table_width,
  input  [6:0]  io_mod_proc_mod_2_mat_mod_table_mod_table_depth,
  input         io_mod_proc_mod_2_act_mod_en_0,
  input         io_mod_proc_mod_2_act_mod_en_1,
  input  [7:0]  io_mod_proc_mod_2_act_mod_addr,
  input  [63:0] io_mod_proc_mod_2_act_mod_data_0,
  input  [63:0] io_mod_proc_mod_2_act_mod_data_1,
  input         io_mod_proc_mod_3_par_mod_en,
  input         io_mod_proc_mod_3_par_mod_last_mau_id_mod,
  input  [1:0]  io_mod_proc_mod_3_par_mod_last_mau_id,
  input  [1:0]  io_mod_proc_mod_3_par_mod_cs,
  input         io_mod_proc_mod_3_par_mod_module_mod_state_id_mod,
  input  [7:0]  io_mod_proc_mod_3_par_mod_module_mod_state_id,
  input         io_mod_proc_mod_3_par_mod_module_mod_sram_w_cs,
  input         io_mod_proc_mod_3_par_mod_module_mod_sram_w_en,
  input  [7:0]  io_mod_proc_mod_3_par_mod_module_mod_sram_w_addr,
  input  [63:0] io_mod_proc_mod_3_par_mod_module_mod_sram_w_data,
  input         io_mod_proc_mod_3_mat_mod_en,
  input         io_mod_proc_mod_3_mat_mod_config_id,
  input  [7:0]  io_mod_proc_mod_3_mat_mod_key_mod_header_id,
  input  [7:0]  io_mod_proc_mod_3_mat_mod_key_mod_internal_offset,
  input  [7:0]  io_mod_proc_mod_3_mat_mod_key_mod_key_length,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_0,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_1,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_2,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_3,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_4,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_5,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_6,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_7,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_8,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_9,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_10,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_11,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_12,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_13,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_14,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_15,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_16,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_17,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_18,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_19,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_20,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_21,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_22,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_23,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_24,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_25,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_26,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_27,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_28,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_29,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_30,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_31,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_32,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_33,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_34,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_35,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_36,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_37,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_38,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_39,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_40,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_41,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_42,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_43,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_44,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_45,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_46,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_47,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_48,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_49,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_50,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_51,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_52,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_53,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_54,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_55,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_56,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_57,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_58,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_59,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_60,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_61,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_62,
  input  [5:0]  io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_63,
  input  [6:0]  io_mod_proc_mod_3_mat_mod_table_mod_table_width,
  input  [6:0]  io_mod_proc_mod_3_mat_mod_table_mod_table_depth,
  input         io_mod_proc_mod_3_act_mod_en_0,
  input         io_mod_proc_mod_3_act_mod_en_1,
  input  [7:0]  io_mod_proc_mod_3_act_mod_addr,
  input  [63:0] io_mod_proc_mod_3_act_mod_data_0,
  input  [63:0] io_mod_proc_mod_3_act_mod_data_1,
  input         io_mod_xbar_mod_en,
  input  [1:0]  io_mod_xbar_mod_first_proc_id,
  input  [1:0]  io_mod_xbar_mod_last_proc_id,
  input  [1:0]  io_mod_xbar_mod_next_proc_id_0,
  input  [1:0]  io_mod_xbar_mod_next_proc_id_1,
  input  [1:0]  io_mod_xbar_mod_next_proc_id_2,
  input  [1:0]  io_mod_xbar_mod_next_proc_id_3,
  input  [5:0]  io_w_0_wcs,
  input         io_w_0_w_en,
  input  [7:0]  io_w_0_w_addr,
  input  [63:0] io_w_0_w_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1561;
  reg [31:0] _RAND_1562;
  reg [31:0] _RAND_1563;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [31:0] _RAND_1566;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [31:0] _RAND_1569;
  reg [31:0] _RAND_1570;
  reg [31:0] _RAND_1571;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1573;
  reg [31:0] _RAND_1574;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [31:0] _RAND_1578;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1581;
  reg [31:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1585;
  reg [31:0] _RAND_1586;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1588;
  reg [31:0] _RAND_1589;
  reg [31:0] _RAND_1590;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1593;
  reg [31:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1597;
  reg [31:0] _RAND_1598;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [31:0] _RAND_1602;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1605;
  reg [31:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1609;
  reg [31:0] _RAND_1610;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [31:0] _RAND_1614;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [31:0] _RAND_1617;
  reg [31:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1621;
  reg [31:0] _RAND_1622;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [31:0] _RAND_1626;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1629;
  reg [31:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1632;
  reg [31:0] _RAND_1633;
  reg [31:0] _RAND_1634;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [31:0] _RAND_1638;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [31:0] _RAND_1641;
  reg [31:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1645;
  reg [31:0] _RAND_1646;
  reg [31:0] _RAND_1647;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [31:0] _RAND_1650;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1653;
  reg [31:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1657;
  reg [31:0] _RAND_1658;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [31:0] _RAND_1662;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1665;
  reg [31:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1668;
  reg [31:0] _RAND_1669;
  reg [31:0] _RAND_1670;
  reg [31:0] _RAND_1671;
  reg [31:0] _RAND_1672;
  reg [31:0] _RAND_1673;
  reg [31:0] _RAND_1674;
  reg [31:0] _RAND_1675;
  reg [31:0] _RAND_1676;
  reg [31:0] _RAND_1677;
  reg [31:0] _RAND_1678;
  reg [31:0] _RAND_1679;
  reg [31:0] _RAND_1680;
  reg [31:0] _RAND_1681;
  reg [31:0] _RAND_1682;
  reg [31:0] _RAND_1683;
  reg [31:0] _RAND_1684;
  reg [31:0] _RAND_1685;
  reg [31:0] _RAND_1686;
  reg [31:0] _RAND_1687;
  reg [31:0] _RAND_1688;
  reg [31:0] _RAND_1689;
  reg [31:0] _RAND_1690;
  reg [31:0] _RAND_1691;
  reg [31:0] _RAND_1692;
  reg [31:0] _RAND_1693;
  reg [31:0] _RAND_1694;
  reg [31:0] _RAND_1695;
  reg [31:0] _RAND_1696;
  reg [31:0] _RAND_1697;
  reg [31:0] _RAND_1698;
  reg [31:0] _RAND_1699;
  reg [31:0] _RAND_1700;
  reg [31:0] _RAND_1701;
  reg [31:0] _RAND_1702;
  reg [31:0] _RAND_1703;
  reg [31:0] _RAND_1704;
  reg [31:0] _RAND_1705;
  reg [31:0] _RAND_1706;
  reg [31:0] _RAND_1707;
  reg [31:0] _RAND_1708;
  reg [31:0] _RAND_1709;
  reg [31:0] _RAND_1710;
  reg [31:0] _RAND_1711;
  reg [31:0] _RAND_1712;
  reg [31:0] _RAND_1713;
  reg [31:0] _RAND_1714;
  reg [31:0] _RAND_1715;
  reg [31:0] _RAND_1716;
  reg [31:0] _RAND_1717;
  reg [31:0] _RAND_1718;
  reg [31:0] _RAND_1719;
  reg [31:0] _RAND_1720;
  reg [31:0] _RAND_1721;
  reg [31:0] _RAND_1722;
  reg [31:0] _RAND_1723;
  reg [31:0] _RAND_1724;
  reg [31:0] _RAND_1725;
  reg [31:0] _RAND_1726;
  reg [31:0] _RAND_1727;
  reg [31:0] _RAND_1728;
  reg [31:0] _RAND_1729;
  reg [31:0] _RAND_1730;
  reg [31:0] _RAND_1731;
  reg [31:0] _RAND_1732;
  reg [31:0] _RAND_1733;
  reg [31:0] _RAND_1734;
  reg [31:0] _RAND_1735;
  reg [31:0] _RAND_1736;
  reg [31:0] _RAND_1737;
  reg [31:0] _RAND_1738;
  reg [31:0] _RAND_1739;
  reg [31:0] _RAND_1740;
  reg [31:0] _RAND_1741;
  reg [31:0] _RAND_1742;
  reg [31:0] _RAND_1743;
  reg [31:0] _RAND_1744;
  reg [31:0] _RAND_1745;
  reg [31:0] _RAND_1746;
  reg [31:0] _RAND_1747;
  reg [31:0] _RAND_1748;
  reg [31:0] _RAND_1749;
  reg [31:0] _RAND_1750;
  reg [31:0] _RAND_1751;
  reg [31:0] _RAND_1752;
  reg [31:0] _RAND_1753;
  reg [31:0] _RAND_1754;
  reg [31:0] _RAND_1755;
  reg [31:0] _RAND_1756;
  reg [31:0] _RAND_1757;
  reg [31:0] _RAND_1758;
  reg [31:0] _RAND_1759;
  reg [31:0] _RAND_1760;
  reg [31:0] _RAND_1761;
  reg [31:0] _RAND_1762;
  reg [31:0] _RAND_1763;
  reg [31:0] _RAND_1764;
  reg [31:0] _RAND_1765;
  reg [31:0] _RAND_1766;
  reg [31:0] _RAND_1767;
  reg [31:0] _RAND_1768;
  reg [31:0] _RAND_1769;
  reg [31:0] _RAND_1770;
  reg [31:0] _RAND_1771;
  reg [31:0] _RAND_1772;
  reg [31:0] _RAND_1773;
  reg [31:0] _RAND_1774;
  reg [31:0] _RAND_1775;
  reg [31:0] _RAND_1776;
  reg [31:0] _RAND_1777;
  reg [31:0] _RAND_1778;
  reg [31:0] _RAND_1779;
  reg [31:0] _RAND_1780;
  reg [31:0] _RAND_1781;
  reg [31:0] _RAND_1782;
  reg [31:0] _RAND_1783;
  reg [31:0] _RAND_1784;
  reg [31:0] _RAND_1785;
  reg [31:0] _RAND_1786;
  reg [31:0] _RAND_1787;
  reg [31:0] _RAND_1788;
  reg [31:0] _RAND_1789;
  reg [31:0] _RAND_1790;
  reg [31:0] _RAND_1791;
  reg [31:0] _RAND_1792;
  reg [31:0] _RAND_1793;
  reg [31:0] _RAND_1794;
  reg [31:0] _RAND_1795;
  reg [31:0] _RAND_1796;
  reg [31:0] _RAND_1797;
  reg [31:0] _RAND_1798;
  reg [31:0] _RAND_1799;
  reg [31:0] _RAND_1800;
  reg [31:0] _RAND_1801;
  reg [31:0] _RAND_1802;
  reg [31:0] _RAND_1803;
  reg [31:0] _RAND_1804;
  reg [31:0] _RAND_1805;
  reg [31:0] _RAND_1806;
  reg [31:0] _RAND_1807;
  reg [31:0] _RAND_1808;
  reg [31:0] _RAND_1809;
  reg [31:0] _RAND_1810;
  reg [31:0] _RAND_1811;
  reg [31:0] _RAND_1812;
  reg [31:0] _RAND_1813;
  reg [31:0] _RAND_1814;
  reg [31:0] _RAND_1815;
  reg [31:0] _RAND_1816;
  reg [31:0] _RAND_1817;
  reg [31:0] _RAND_1818;
  reg [31:0] _RAND_1819;
  reg [31:0] _RAND_1820;
  reg [31:0] _RAND_1821;
  reg [31:0] _RAND_1822;
  reg [31:0] _RAND_1823;
  reg [31:0] _RAND_1824;
  reg [31:0] _RAND_1825;
  reg [31:0] _RAND_1826;
  reg [31:0] _RAND_1827;
  reg [31:0] _RAND_1828;
  reg [31:0] _RAND_1829;
  reg [31:0] _RAND_1830;
  reg [31:0] _RAND_1831;
  reg [31:0] _RAND_1832;
  reg [31:0] _RAND_1833;
  reg [31:0] _RAND_1834;
  reg [31:0] _RAND_1835;
  reg [31:0] _RAND_1836;
  reg [31:0] _RAND_1837;
  reg [31:0] _RAND_1838;
  reg [31:0] _RAND_1839;
  reg [31:0] _RAND_1840;
  reg [31:0] _RAND_1841;
  reg [31:0] _RAND_1842;
  reg [31:0] _RAND_1843;
  reg [31:0] _RAND_1844;
  reg [31:0] _RAND_1845;
  reg [31:0] _RAND_1846;
  reg [31:0] _RAND_1847;
  reg [31:0] _RAND_1848;
  reg [31:0] _RAND_1849;
  reg [31:0] _RAND_1850;
  reg [31:0] _RAND_1851;
  reg [31:0] _RAND_1852;
  reg [31:0] _RAND_1853;
  reg [31:0] _RAND_1854;
  reg [31:0] _RAND_1855;
  reg [31:0] _RAND_1856;
  reg [31:0] _RAND_1857;
  reg [31:0] _RAND_1858;
  reg [31:0] _RAND_1859;
  reg [31:0] _RAND_1860;
  reg [31:0] _RAND_1861;
  reg [31:0] _RAND_1862;
  reg [31:0] _RAND_1863;
  reg [31:0] _RAND_1864;
  reg [31:0] _RAND_1865;
  reg [31:0] _RAND_1866;
  reg [31:0] _RAND_1867;
  reg [31:0] _RAND_1868;
  reg [31:0] _RAND_1869;
  reg [31:0] _RAND_1870;
  reg [31:0] _RAND_1871;
  reg [31:0] _RAND_1872;
  reg [31:0] _RAND_1873;
  reg [31:0] _RAND_1874;
  reg [31:0] _RAND_1875;
  reg [31:0] _RAND_1876;
  reg [31:0] _RAND_1877;
  reg [31:0] _RAND_1878;
  reg [31:0] _RAND_1879;
  reg [31:0] _RAND_1880;
  reg [31:0] _RAND_1881;
  reg [31:0] _RAND_1882;
  reg [31:0] _RAND_1883;
  reg [31:0] _RAND_1884;
  reg [31:0] _RAND_1885;
  reg [31:0] _RAND_1886;
  reg [31:0] _RAND_1887;
  reg [31:0] _RAND_1888;
  reg [31:0] _RAND_1889;
  reg [31:0] _RAND_1890;
  reg [31:0] _RAND_1891;
  reg [31:0] _RAND_1892;
  reg [31:0] _RAND_1893;
  reg [31:0] _RAND_1894;
  reg [31:0] _RAND_1895;
  reg [31:0] _RAND_1896;
  reg [31:0] _RAND_1897;
  reg [31:0] _RAND_1898;
  reg [31:0] _RAND_1899;
  reg [31:0] _RAND_1900;
  reg [31:0] _RAND_1901;
  reg [31:0] _RAND_1902;
  reg [31:0] _RAND_1903;
  reg [31:0] _RAND_1904;
  reg [31:0] _RAND_1905;
  reg [31:0] _RAND_1906;
  reg [31:0] _RAND_1907;
  reg [31:0] _RAND_1908;
  reg [31:0] _RAND_1909;
  reg [31:0] _RAND_1910;
  reg [31:0] _RAND_1911;
  reg [31:0] _RAND_1912;
  reg [31:0] _RAND_1913;
  reg [31:0] _RAND_1914;
  reg [31:0] _RAND_1915;
  reg [31:0] _RAND_1916;
  reg [31:0] _RAND_1917;
  reg [31:0] _RAND_1918;
  reg [31:0] _RAND_1919;
  reg [31:0] _RAND_1920;
  reg [31:0] _RAND_1921;
  reg [31:0] _RAND_1922;
  reg [31:0] _RAND_1923;
  reg [31:0] _RAND_1924;
  reg [31:0] _RAND_1925;
  reg [31:0] _RAND_1926;
  reg [31:0] _RAND_1927;
  reg [31:0] _RAND_1928;
  reg [31:0] _RAND_1929;
  reg [31:0] _RAND_1930;
  reg [31:0] _RAND_1931;
  reg [31:0] _RAND_1932;
  reg [31:0] _RAND_1933;
  reg [31:0] _RAND_1934;
  reg [31:0] _RAND_1935;
  reg [31:0] _RAND_1936;
  reg [31:0] _RAND_1937;
  reg [31:0] _RAND_1938;
  reg [31:0] _RAND_1939;
  reg [31:0] _RAND_1940;
  reg [31:0] _RAND_1941;
  reg [31:0] _RAND_1942;
  reg [31:0] _RAND_1943;
  reg [31:0] _RAND_1944;
  reg [31:0] _RAND_1945;
  reg [31:0] _RAND_1946;
  reg [31:0] _RAND_1947;
  reg [31:0] _RAND_1948;
  reg [31:0] _RAND_1949;
  reg [31:0] _RAND_1950;
  reg [31:0] _RAND_1951;
  reg [31:0] _RAND_1952;
  reg [31:0] _RAND_1953;
  reg [31:0] _RAND_1954;
  reg [31:0] _RAND_1955;
  reg [31:0] _RAND_1956;
  reg [31:0] _RAND_1957;
  reg [31:0] _RAND_1958;
  reg [31:0] _RAND_1959;
  reg [31:0] _RAND_1960;
  reg [31:0] _RAND_1961;
  reg [31:0] _RAND_1962;
  reg [31:0] _RAND_1963;
  reg [31:0] _RAND_1964;
  reg [31:0] _RAND_1965;
  reg [31:0] _RAND_1966;
  reg [31:0] _RAND_1967;
  reg [31:0] _RAND_1968;
  reg [31:0] _RAND_1969;
  reg [31:0] _RAND_1970;
  reg [31:0] _RAND_1971;
  reg [31:0] _RAND_1972;
  reg [31:0] _RAND_1973;
  reg [31:0] _RAND_1974;
  reg [31:0] _RAND_1975;
  reg [31:0] _RAND_1976;
  reg [31:0] _RAND_1977;
  reg [31:0] _RAND_1978;
  reg [31:0] _RAND_1979;
  reg [31:0] _RAND_1980;
  reg [31:0] _RAND_1981;
  reg [31:0] _RAND_1982;
  reg [31:0] _RAND_1983;
  reg [31:0] _RAND_1984;
  reg [31:0] _RAND_1985;
  reg [31:0] _RAND_1986;
  reg [31:0] _RAND_1987;
  reg [31:0] _RAND_1988;
  reg [31:0] _RAND_1989;
  reg [31:0] _RAND_1990;
  reg [31:0] _RAND_1991;
  reg [31:0] _RAND_1992;
  reg [31:0] _RAND_1993;
  reg [31:0] _RAND_1994;
  reg [31:0] _RAND_1995;
  reg [31:0] _RAND_1996;
  reg [31:0] _RAND_1997;
  reg [31:0] _RAND_1998;
  reg [31:0] _RAND_1999;
  reg [31:0] _RAND_2000;
  reg [31:0] _RAND_2001;
  reg [31:0] _RAND_2002;
  reg [31:0] _RAND_2003;
  reg [31:0] _RAND_2004;
  reg [31:0] _RAND_2005;
  reg [31:0] _RAND_2006;
  reg [31:0] _RAND_2007;
  reg [31:0] _RAND_2008;
  reg [31:0] _RAND_2009;
  reg [31:0] _RAND_2010;
  reg [31:0] _RAND_2011;
  reg [31:0] _RAND_2012;
  reg [31:0] _RAND_2013;
  reg [31:0] _RAND_2014;
  reg [31:0] _RAND_2015;
  reg [31:0] _RAND_2016;
  reg [31:0] _RAND_2017;
  reg [31:0] _RAND_2018;
  reg [31:0] _RAND_2019;
  reg [31:0] _RAND_2020;
  reg [31:0] _RAND_2021;
  reg [31:0] _RAND_2022;
  reg [31:0] _RAND_2023;
  reg [31:0] _RAND_2024;
  reg [31:0] _RAND_2025;
  reg [31:0] _RAND_2026;
  reg [31:0] _RAND_2027;
  reg [31:0] _RAND_2028;
  reg [31:0] _RAND_2029;
  reg [31:0] _RAND_2030;
  reg [31:0] _RAND_2031;
  reg [31:0] _RAND_2032;
  reg [31:0] _RAND_2033;
  reg [31:0] _RAND_2034;
  reg [31:0] _RAND_2035;
  reg [31:0] _RAND_2036;
  reg [31:0] _RAND_2037;
  reg [31:0] _RAND_2038;
  reg [31:0] _RAND_2039;
  reg [31:0] _RAND_2040;
  reg [31:0] _RAND_2041;
  reg [31:0] _RAND_2042;
  reg [31:0] _RAND_2043;
  reg [31:0] _RAND_2044;
  reg [31:0] _RAND_2045;
  reg [31:0] _RAND_2046;
  reg [31:0] _RAND_2047;
  reg [31:0] _RAND_2048;
  reg [31:0] _RAND_2049;
  reg [31:0] _RAND_2050;
  reg [31:0] _RAND_2051;
  reg [31:0] _RAND_2052;
  reg [31:0] _RAND_2053;
  reg [31:0] _RAND_2054;
  reg [31:0] _RAND_2055;
  reg [31:0] _RAND_2056;
  reg [31:0] _RAND_2057;
  reg [31:0] _RAND_2058;
  reg [31:0] _RAND_2059;
  reg [31:0] _RAND_2060;
  reg [31:0] _RAND_2061;
  reg [31:0] _RAND_2062;
  reg [31:0] _RAND_2063;
  reg [31:0] _RAND_2064;
  reg [31:0] _RAND_2065;
  reg [31:0] _RAND_2066;
  reg [31:0] _RAND_2067;
  reg [31:0] _RAND_2068;
  reg [31:0] _RAND_2069;
  reg [31:0] _RAND_2070;
  reg [31:0] _RAND_2071;
  reg [31:0] _RAND_2072;
  reg [31:0] _RAND_2073;
  reg [31:0] _RAND_2074;
  reg [31:0] _RAND_2075;
  reg [31:0] _RAND_2076;
  reg [31:0] _RAND_2077;
  reg [31:0] _RAND_2078;
  reg [31:0] _RAND_2079;
  reg [31:0] _RAND_2080;
  reg [31:0] _RAND_2081;
  reg [31:0] _RAND_2082;
  reg [31:0] _RAND_2083;
  reg [31:0] _RAND_2084;
  reg [31:0] _RAND_2085;
  reg [31:0] _RAND_2086;
  reg [31:0] _RAND_2087;
  reg [31:0] _RAND_2088;
  reg [31:0] _RAND_2089;
  reg [31:0] _RAND_2090;
  reg [31:0] _RAND_2091;
  reg [31:0] _RAND_2092;
  reg [31:0] _RAND_2093;
  reg [31:0] _RAND_2094;
  reg [31:0] _RAND_2095;
  reg [31:0] _RAND_2096;
  reg [31:0] _RAND_2097;
  reg [31:0] _RAND_2098;
  reg [31:0] _RAND_2099;
  reg [31:0] _RAND_2100;
  reg [31:0] _RAND_2101;
  reg [31:0] _RAND_2102;
  reg [31:0] _RAND_2103;
  reg [31:0] _RAND_2104;
  reg [31:0] _RAND_2105;
  reg [31:0] _RAND_2106;
  reg [31:0] _RAND_2107;
  reg [31:0] _RAND_2108;
  reg [31:0] _RAND_2109;
  reg [31:0] _RAND_2110;
  reg [31:0] _RAND_2111;
  reg [31:0] _RAND_2112;
  reg [31:0] _RAND_2113;
  reg [31:0] _RAND_2114;
  reg [31:0] _RAND_2115;
  reg [31:0] _RAND_2116;
  reg [31:0] _RAND_2117;
  reg [31:0] _RAND_2118;
  reg [31:0] _RAND_2119;
  reg [31:0] _RAND_2120;
  reg [31:0] _RAND_2121;
  reg [31:0] _RAND_2122;
  reg [31:0] _RAND_2123;
  reg [31:0] _RAND_2124;
  reg [31:0] _RAND_2125;
  reg [31:0] _RAND_2126;
  reg [31:0] _RAND_2127;
  reg [31:0] _RAND_2128;
  reg [31:0] _RAND_2129;
  reg [31:0] _RAND_2130;
  reg [31:0] _RAND_2131;
  reg [31:0] _RAND_2132;
  reg [31:0] _RAND_2133;
  reg [31:0] _RAND_2134;
  reg [31:0] _RAND_2135;
  reg [31:0] _RAND_2136;
  reg [31:0] _RAND_2137;
  reg [31:0] _RAND_2138;
  reg [31:0] _RAND_2139;
  reg [31:0] _RAND_2140;
  reg [31:0] _RAND_2141;
  reg [31:0] _RAND_2142;
  reg [31:0] _RAND_2143;
  reg [31:0] _RAND_2144;
  reg [31:0] _RAND_2145;
  reg [31:0] _RAND_2146;
  reg [31:0] _RAND_2147;
  reg [31:0] _RAND_2148;
  reg [31:0] _RAND_2149;
  reg [31:0] _RAND_2150;
  reg [31:0] _RAND_2151;
  reg [31:0] _RAND_2152;
  reg [31:0] _RAND_2153;
  reg [31:0] _RAND_2154;
  reg [31:0] _RAND_2155;
  reg [31:0] _RAND_2156;
  reg [31:0] _RAND_2157;
  reg [31:0] _RAND_2158;
  reg [31:0] _RAND_2159;
  reg [31:0] _RAND_2160;
  reg [31:0] _RAND_2161;
  reg [31:0] _RAND_2162;
  reg [31:0] _RAND_2163;
  reg [31:0] _RAND_2164;
  reg [31:0] _RAND_2165;
  reg [31:0] _RAND_2166;
  reg [31:0] _RAND_2167;
  reg [31:0] _RAND_2168;
  reg [31:0] _RAND_2169;
  reg [31:0] _RAND_2170;
  reg [31:0] _RAND_2171;
  reg [31:0] _RAND_2172;
  reg [31:0] _RAND_2173;
  reg [31:0] _RAND_2174;
  reg [31:0] _RAND_2175;
  reg [31:0] _RAND_2176;
  reg [31:0] _RAND_2177;
  reg [31:0] _RAND_2178;
  reg [31:0] _RAND_2179;
  reg [31:0] _RAND_2180;
  reg [31:0] _RAND_2181;
  reg [31:0] _RAND_2182;
  reg [31:0] _RAND_2183;
  reg [31:0] _RAND_2184;
  reg [31:0] _RAND_2185;
  reg [31:0] _RAND_2186;
  reg [31:0] _RAND_2187;
  reg [31:0] _RAND_2188;
  reg [31:0] _RAND_2189;
  reg [31:0] _RAND_2190;
  reg [31:0] _RAND_2191;
  reg [31:0] _RAND_2192;
  reg [31:0] _RAND_2193;
  reg [31:0] _RAND_2194;
  reg [31:0] _RAND_2195;
  reg [31:0] _RAND_2196;
  reg [31:0] _RAND_2197;
  reg [31:0] _RAND_2198;
  reg [31:0] _RAND_2199;
  reg [31:0] _RAND_2200;
  reg [31:0] _RAND_2201;
  reg [31:0] _RAND_2202;
  reg [31:0] _RAND_2203;
  reg [31:0] _RAND_2204;
  reg [31:0] _RAND_2205;
  reg [31:0] _RAND_2206;
  reg [31:0] _RAND_2207;
  reg [31:0] _RAND_2208;
  reg [31:0] _RAND_2209;
  reg [31:0] _RAND_2210;
  reg [31:0] _RAND_2211;
  reg [31:0] _RAND_2212;
  reg [31:0] _RAND_2213;
  reg [31:0] _RAND_2214;
  reg [31:0] _RAND_2215;
  reg [31:0] _RAND_2216;
  reg [31:0] _RAND_2217;
  reg [31:0] _RAND_2218;
  reg [31:0] _RAND_2219;
  reg [31:0] _RAND_2220;
  reg [31:0] _RAND_2221;
  reg [31:0] _RAND_2222;
  reg [31:0] _RAND_2223;
  reg [31:0] _RAND_2224;
  reg [31:0] _RAND_2225;
  reg [31:0] _RAND_2226;
  reg [31:0] _RAND_2227;
  reg [31:0] _RAND_2228;
  reg [31:0] _RAND_2229;
  reg [31:0] _RAND_2230;
  reg [31:0] _RAND_2231;
  reg [31:0] _RAND_2232;
  reg [31:0] _RAND_2233;
  reg [31:0] _RAND_2234;
  reg [31:0] _RAND_2235;
  reg [31:0] _RAND_2236;
  reg [31:0] _RAND_2237;
  reg [31:0] _RAND_2238;
  reg [31:0] _RAND_2239;
  reg [31:0] _RAND_2240;
  reg [31:0] _RAND_2241;
  reg [31:0] _RAND_2242;
  reg [31:0] _RAND_2243;
  reg [31:0] _RAND_2244;
  reg [31:0] _RAND_2245;
  reg [31:0] _RAND_2246;
  reg [31:0] _RAND_2247;
  reg [31:0] _RAND_2248;
  reg [31:0] _RAND_2249;
  reg [31:0] _RAND_2250;
  reg [31:0] _RAND_2251;
  reg [31:0] _RAND_2252;
  reg [31:0] _RAND_2253;
  reg [31:0] _RAND_2254;
  reg [31:0] _RAND_2255;
  reg [31:0] _RAND_2256;
  reg [31:0] _RAND_2257;
  reg [31:0] _RAND_2258;
  reg [31:0] _RAND_2259;
  reg [31:0] _RAND_2260;
  reg [31:0] _RAND_2261;
  reg [31:0] _RAND_2262;
  reg [31:0] _RAND_2263;
  reg [31:0] _RAND_2264;
  reg [31:0] _RAND_2265;
  reg [31:0] _RAND_2266;
  reg [31:0] _RAND_2267;
  reg [31:0] _RAND_2268;
  reg [31:0] _RAND_2269;
  reg [31:0] _RAND_2270;
  reg [31:0] _RAND_2271;
  reg [31:0] _RAND_2272;
  reg [31:0] _RAND_2273;
  reg [31:0] _RAND_2274;
  reg [31:0] _RAND_2275;
  reg [31:0] _RAND_2276;
  reg [31:0] _RAND_2277;
  reg [31:0] _RAND_2278;
  reg [31:0] _RAND_2279;
  reg [31:0] _RAND_2280;
  reg [31:0] _RAND_2281;
  reg [31:0] _RAND_2282;
  reg [31:0] _RAND_2283;
  reg [31:0] _RAND_2284;
  reg [31:0] _RAND_2285;
  reg [31:0] _RAND_2286;
  reg [31:0] _RAND_2287;
  reg [31:0] _RAND_2288;
  reg [31:0] _RAND_2289;
  reg [31:0] _RAND_2290;
  reg [31:0] _RAND_2291;
  reg [31:0] _RAND_2292;
  reg [31:0] _RAND_2293;
  reg [31:0] _RAND_2294;
  reg [31:0] _RAND_2295;
  reg [31:0] _RAND_2296;
  reg [31:0] _RAND_2297;
  reg [31:0] _RAND_2298;
  reg [31:0] _RAND_2299;
  reg [31:0] _RAND_2300;
  reg [31:0] _RAND_2301;
  reg [31:0] _RAND_2302;
  reg [31:0] _RAND_2303;
  reg [31:0] _RAND_2304;
  reg [31:0] _RAND_2305;
  reg [31:0] _RAND_2306;
  reg [31:0] _RAND_2307;
  reg [31:0] _RAND_2308;
  reg [31:0] _RAND_2309;
  reg [31:0] _RAND_2310;
  reg [31:0] _RAND_2311;
  reg [31:0] _RAND_2312;
  reg [31:0] _RAND_2313;
  reg [31:0] _RAND_2314;
  reg [31:0] _RAND_2315;
  reg [31:0] _RAND_2316;
  reg [31:0] _RAND_2317;
  reg [31:0] _RAND_2318;
  reg [31:0] _RAND_2319;
  reg [31:0] _RAND_2320;
  reg [31:0] _RAND_2321;
  reg [31:0] _RAND_2322;
  reg [31:0] _RAND_2323;
  reg [31:0] _RAND_2324;
  reg [31:0] _RAND_2325;
  reg [31:0] _RAND_2326;
  reg [31:0] _RAND_2327;
  reg [31:0] _RAND_2328;
  reg [31:0] _RAND_2329;
  reg [31:0] _RAND_2330;
  reg [31:0] _RAND_2331;
  reg [31:0] _RAND_2332;
  reg [31:0] _RAND_2333;
  reg [31:0] _RAND_2334;
  reg [31:0] _RAND_2335;
  reg [31:0] _RAND_2336;
  reg [31:0] _RAND_2337;
  reg [31:0] _RAND_2338;
  reg [31:0] _RAND_2339;
  reg [31:0] _RAND_2340;
  reg [31:0] _RAND_2341;
  reg [31:0] _RAND_2342;
  reg [31:0] _RAND_2343;
  reg [31:0] _RAND_2344;
  reg [31:0] _RAND_2345;
  reg [31:0] _RAND_2346;
  reg [31:0] _RAND_2347;
  reg [31:0] _RAND_2348;
  reg [31:0] _RAND_2349;
  reg [31:0] _RAND_2350;
  reg [31:0] _RAND_2351;
  reg [31:0] _RAND_2352;
  reg [31:0] _RAND_2353;
  reg [31:0] _RAND_2354;
  reg [31:0] _RAND_2355;
  reg [31:0] _RAND_2356;
  reg [31:0] _RAND_2357;
  reg [31:0] _RAND_2358;
  reg [31:0] _RAND_2359;
  reg [31:0] _RAND_2360;
  reg [31:0] _RAND_2361;
  reg [31:0] _RAND_2362;
  reg [31:0] _RAND_2363;
  reg [31:0] _RAND_2364;
  reg [31:0] _RAND_2365;
  reg [31:0] _RAND_2366;
  reg [31:0] _RAND_2367;
  reg [31:0] _RAND_2368;
  reg [31:0] _RAND_2369;
  reg [31:0] _RAND_2370;
  reg [31:0] _RAND_2371;
  reg [31:0] _RAND_2372;
  reg [31:0] _RAND_2373;
  reg [31:0] _RAND_2374;
  reg [31:0] _RAND_2375;
  reg [31:0] _RAND_2376;
  reg [31:0] _RAND_2377;
  reg [31:0] _RAND_2378;
  reg [31:0] _RAND_2379;
  reg [31:0] _RAND_2380;
  reg [31:0] _RAND_2381;
  reg [31:0] _RAND_2382;
  reg [31:0] _RAND_2383;
  reg [31:0] _RAND_2384;
  reg [31:0] _RAND_2385;
  reg [31:0] _RAND_2386;
  reg [31:0] _RAND_2387;
  reg [31:0] _RAND_2388;
  reg [31:0] _RAND_2389;
  reg [31:0] _RAND_2390;
  reg [31:0] _RAND_2391;
  reg [31:0] _RAND_2392;
  reg [31:0] _RAND_2393;
  reg [31:0] _RAND_2394;
  reg [31:0] _RAND_2395;
  reg [31:0] _RAND_2396;
  reg [31:0] _RAND_2397;
  reg [31:0] _RAND_2398;
  reg [31:0] _RAND_2399;
  reg [31:0] _RAND_2400;
  reg [31:0] _RAND_2401;
  reg [31:0] _RAND_2402;
  reg [31:0] _RAND_2403;
  reg [31:0] _RAND_2404;
  reg [31:0] _RAND_2405;
  reg [31:0] _RAND_2406;
  reg [31:0] _RAND_2407;
  reg [31:0] _RAND_2408;
  reg [31:0] _RAND_2409;
  reg [31:0] _RAND_2410;
  reg [31:0] _RAND_2411;
  reg [31:0] _RAND_2412;
  reg [31:0] _RAND_2413;
  reg [31:0] _RAND_2414;
  reg [31:0] _RAND_2415;
  reg [31:0] _RAND_2416;
  reg [31:0] _RAND_2417;
  reg [31:0] _RAND_2418;
  reg [31:0] _RAND_2419;
  reg [31:0] _RAND_2420;
  reg [31:0] _RAND_2421;
  reg [31:0] _RAND_2422;
  reg [31:0] _RAND_2423;
  reg [31:0] _RAND_2424;
  reg [31:0] _RAND_2425;
  reg [31:0] _RAND_2426;
  reg [31:0] _RAND_2427;
  reg [31:0] _RAND_2428;
  reg [31:0] _RAND_2429;
  reg [31:0] _RAND_2430;
  reg [31:0] _RAND_2431;
  reg [31:0] _RAND_2432;
  reg [31:0] _RAND_2433;
  reg [31:0] _RAND_2434;
  reg [31:0] _RAND_2435;
  reg [31:0] _RAND_2436;
  reg [31:0] _RAND_2437;
  reg [31:0] _RAND_2438;
  reg [31:0] _RAND_2439;
  reg [31:0] _RAND_2440;
  reg [31:0] _RAND_2441;
  reg [31:0] _RAND_2442;
  reg [31:0] _RAND_2443;
  reg [31:0] _RAND_2444;
  reg [31:0] _RAND_2445;
  reg [31:0] _RAND_2446;
  reg [31:0] _RAND_2447;
  reg [31:0] _RAND_2448;
  reg [31:0] _RAND_2449;
  reg [31:0] _RAND_2450;
  reg [31:0] _RAND_2451;
  reg [31:0] _RAND_2452;
  reg [31:0] _RAND_2453;
  reg [31:0] _RAND_2454;
  reg [31:0] _RAND_2455;
  reg [31:0] _RAND_2456;
  reg [31:0] _RAND_2457;
  reg [31:0] _RAND_2458;
  reg [31:0] _RAND_2459;
  reg [31:0] _RAND_2460;
  reg [31:0] _RAND_2461;
  reg [31:0] _RAND_2462;
  reg [31:0] _RAND_2463;
  reg [31:0] _RAND_2464;
  reg [31:0] _RAND_2465;
  reg [31:0] _RAND_2466;
  reg [31:0] _RAND_2467;
  reg [31:0] _RAND_2468;
  reg [31:0] _RAND_2469;
  reg [31:0] _RAND_2470;
  reg [31:0] _RAND_2471;
  reg [31:0] _RAND_2472;
  reg [31:0] _RAND_2473;
  reg [31:0] _RAND_2474;
  reg [31:0] _RAND_2475;
  reg [31:0] _RAND_2476;
  reg [31:0] _RAND_2477;
  reg [31:0] _RAND_2478;
  reg [31:0] _RAND_2479;
  reg [31:0] _RAND_2480;
  reg [31:0] _RAND_2481;
  reg [31:0] _RAND_2482;
  reg [31:0] _RAND_2483;
  reg [31:0] _RAND_2484;
  reg [31:0] _RAND_2485;
  reg [31:0] _RAND_2486;
  reg [31:0] _RAND_2487;
  reg [31:0] _RAND_2488;
  reg [31:0] _RAND_2489;
  reg [31:0] _RAND_2490;
  reg [31:0] _RAND_2491;
  reg [31:0] _RAND_2492;
  reg [31:0] _RAND_2493;
  reg [31:0] _RAND_2494;
  reg [31:0] _RAND_2495;
  reg [31:0] _RAND_2496;
  reg [31:0] _RAND_2497;
  reg [31:0] _RAND_2498;
  reg [31:0] _RAND_2499;
  reg [31:0] _RAND_2500;
  reg [31:0] _RAND_2501;
  reg [31:0] _RAND_2502;
  reg [31:0] _RAND_2503;
  reg [31:0] _RAND_2504;
  reg [31:0] _RAND_2505;
  reg [31:0] _RAND_2506;
  reg [31:0] _RAND_2507;
  reg [31:0] _RAND_2508;
  reg [31:0] _RAND_2509;
  reg [31:0] _RAND_2510;
  reg [31:0] _RAND_2511;
  reg [31:0] _RAND_2512;
  reg [31:0] _RAND_2513;
  reg [31:0] _RAND_2514;
  reg [31:0] _RAND_2515;
  reg [31:0] _RAND_2516;
  reg [31:0] _RAND_2517;
  reg [31:0] _RAND_2518;
  reg [31:0] _RAND_2519;
  reg [31:0] _RAND_2520;
  reg [31:0] _RAND_2521;
  reg [31:0] _RAND_2522;
  reg [31:0] _RAND_2523;
  reg [31:0] _RAND_2524;
  reg [31:0] _RAND_2525;
  reg [31:0] _RAND_2526;
  reg [31:0] _RAND_2527;
  reg [31:0] _RAND_2528;
  reg [31:0] _RAND_2529;
  reg [31:0] _RAND_2530;
  reg [31:0] _RAND_2531;
  reg [31:0] _RAND_2532;
  reg [31:0] _RAND_2533;
  reg [31:0] _RAND_2534;
  reg [31:0] _RAND_2535;
  reg [31:0] _RAND_2536;
  reg [31:0] _RAND_2537;
  reg [31:0] _RAND_2538;
  reg [31:0] _RAND_2539;
  reg [31:0] _RAND_2540;
  reg [31:0] _RAND_2541;
  reg [31:0] _RAND_2542;
  reg [31:0] _RAND_2543;
  reg [31:0] _RAND_2544;
  reg [31:0] _RAND_2545;
  reg [31:0] _RAND_2546;
  reg [31:0] _RAND_2547;
  reg [31:0] _RAND_2548;
  reg [31:0] _RAND_2549;
  reg [31:0] _RAND_2550;
  reg [31:0] _RAND_2551;
  reg [31:0] _RAND_2552;
  reg [31:0] _RAND_2553;
  reg [31:0] _RAND_2554;
  reg [31:0] _RAND_2555;
  reg [31:0] _RAND_2556;
  reg [31:0] _RAND_2557;
  reg [31:0] _RAND_2558;
  reg [31:0] _RAND_2559;
  reg [31:0] _RAND_2560;
  reg [31:0] _RAND_2561;
  reg [31:0] _RAND_2562;
  reg [31:0] _RAND_2563;
  reg [31:0] _RAND_2564;
  reg [31:0] _RAND_2565;
  reg [31:0] _RAND_2566;
  reg [31:0] _RAND_2567;
  reg [31:0] _RAND_2568;
  reg [31:0] _RAND_2569;
  reg [31:0] _RAND_2570;
  reg [31:0] _RAND_2571;
  reg [31:0] _RAND_2572;
  reg [31:0] _RAND_2573;
  reg [31:0] _RAND_2574;
  reg [31:0] _RAND_2575;
  reg [31:0] _RAND_2576;
  reg [31:0] _RAND_2577;
  reg [31:0] _RAND_2578;
  reg [31:0] _RAND_2579;
  reg [31:0] _RAND_2580;
  reg [31:0] _RAND_2581;
  reg [31:0] _RAND_2582;
  reg [31:0] _RAND_2583;
  reg [31:0] _RAND_2584;
  reg [31:0] _RAND_2585;
  reg [31:0] _RAND_2586;
  reg [31:0] _RAND_2587;
  reg [31:0] _RAND_2588;
  reg [31:0] _RAND_2589;
  reg [31:0] _RAND_2590;
  reg [31:0] _RAND_2591;
  reg [31:0] _RAND_2592;
  reg [31:0] _RAND_2593;
  reg [31:0] _RAND_2594;
  reg [31:0] _RAND_2595;
  reg [31:0] _RAND_2596;
  reg [31:0] _RAND_2597;
  reg [31:0] _RAND_2598;
  reg [31:0] _RAND_2599;
  reg [31:0] _RAND_2600;
  reg [31:0] _RAND_2601;
  reg [31:0] _RAND_2602;
  reg [31:0] _RAND_2603;
  reg [31:0] _RAND_2604;
  reg [31:0] _RAND_2605;
  reg [31:0] _RAND_2606;
  reg [31:0] _RAND_2607;
  reg [31:0] _RAND_2608;
  reg [31:0] _RAND_2609;
  reg [31:0] _RAND_2610;
  reg [31:0] _RAND_2611;
  reg [31:0] _RAND_2612;
  reg [31:0] _RAND_2613;
  reg [31:0] _RAND_2614;
  reg [31:0] _RAND_2615;
  reg [31:0] _RAND_2616;
  reg [31:0] _RAND_2617;
  reg [31:0] _RAND_2618;
  reg [31:0] _RAND_2619;
  reg [31:0] _RAND_2620;
  reg [31:0] _RAND_2621;
  reg [31:0] _RAND_2622;
  reg [31:0] _RAND_2623;
  reg [31:0] _RAND_2624;
  reg [31:0] _RAND_2625;
  reg [31:0] _RAND_2626;
  reg [31:0] _RAND_2627;
  reg [31:0] _RAND_2628;
  reg [31:0] _RAND_2629;
  reg [31:0] _RAND_2630;
  reg [31:0] _RAND_2631;
  reg [31:0] _RAND_2632;
  reg [31:0] _RAND_2633;
  reg [31:0] _RAND_2634;
  reg [31:0] _RAND_2635;
  reg [31:0] _RAND_2636;
  reg [31:0] _RAND_2637;
  reg [31:0] _RAND_2638;
  reg [31:0] _RAND_2639;
  reg [31:0] _RAND_2640;
  reg [31:0] _RAND_2641;
  reg [31:0] _RAND_2642;
  reg [31:0] _RAND_2643;
  reg [31:0] _RAND_2644;
  reg [31:0] _RAND_2645;
  reg [31:0] _RAND_2646;
  reg [31:0] _RAND_2647;
  reg [31:0] _RAND_2648;
  reg [31:0] _RAND_2649;
  reg [31:0] _RAND_2650;
  reg [31:0] _RAND_2651;
  reg [31:0] _RAND_2652;
  reg [31:0] _RAND_2653;
  reg [31:0] _RAND_2654;
  reg [31:0] _RAND_2655;
  reg [31:0] _RAND_2656;
  reg [31:0] _RAND_2657;
  reg [31:0] _RAND_2658;
  reg [31:0] _RAND_2659;
  reg [31:0] _RAND_2660;
  reg [31:0] _RAND_2661;
  reg [31:0] _RAND_2662;
  reg [31:0] _RAND_2663;
  reg [31:0] _RAND_2664;
  reg [31:0] _RAND_2665;
  reg [31:0] _RAND_2666;
  reg [31:0] _RAND_2667;
  reg [31:0] _RAND_2668;
  reg [31:0] _RAND_2669;
  reg [31:0] _RAND_2670;
  reg [31:0] _RAND_2671;
  reg [31:0] _RAND_2672;
  reg [31:0] _RAND_2673;
  reg [31:0] _RAND_2674;
  reg [31:0] _RAND_2675;
  reg [31:0] _RAND_2676;
  reg [31:0] _RAND_2677;
  reg [31:0] _RAND_2678;
  reg [31:0] _RAND_2679;
  reg [31:0] _RAND_2680;
  reg [31:0] _RAND_2681;
  reg [31:0] _RAND_2682;
  reg [31:0] _RAND_2683;
  reg [31:0] _RAND_2684;
  reg [31:0] _RAND_2685;
  reg [31:0] _RAND_2686;
  reg [31:0] _RAND_2687;
  reg [31:0] _RAND_2688;
  reg [31:0] _RAND_2689;
  reg [31:0] _RAND_2690;
  reg [31:0] _RAND_2691;
  reg [31:0] _RAND_2692;
  reg [31:0] _RAND_2693;
  reg [31:0] _RAND_2694;
  reg [31:0] _RAND_2695;
  reg [31:0] _RAND_2696;
  reg [31:0] _RAND_2697;
  reg [31:0] _RAND_2698;
  reg [31:0] _RAND_2699;
  reg [31:0] _RAND_2700;
  reg [31:0] _RAND_2701;
  reg [31:0] _RAND_2702;
  reg [31:0] _RAND_2703;
  reg [31:0] _RAND_2704;
  reg [31:0] _RAND_2705;
  reg [31:0] _RAND_2706;
  reg [31:0] _RAND_2707;
  reg [31:0] _RAND_2708;
  reg [31:0] _RAND_2709;
  reg [31:0] _RAND_2710;
  reg [31:0] _RAND_2711;
  reg [31:0] _RAND_2712;
  reg [31:0] _RAND_2713;
  reg [31:0] _RAND_2714;
  reg [31:0] _RAND_2715;
  reg [31:0] _RAND_2716;
  reg [31:0] _RAND_2717;
  reg [31:0] _RAND_2718;
  reg [31:0] _RAND_2719;
  reg [31:0] _RAND_2720;
  reg [31:0] _RAND_2721;
  reg [31:0] _RAND_2722;
  reg [31:0] _RAND_2723;
  reg [31:0] _RAND_2724;
  reg [31:0] _RAND_2725;
  reg [31:0] _RAND_2726;
  reg [31:0] _RAND_2727;
  reg [31:0] _RAND_2728;
  reg [31:0] _RAND_2729;
  reg [31:0] _RAND_2730;
  reg [31:0] _RAND_2731;
  reg [31:0] _RAND_2732;
  reg [31:0] _RAND_2733;
  reg [31:0] _RAND_2734;
  reg [31:0] _RAND_2735;
  reg [31:0] _RAND_2736;
  reg [31:0] _RAND_2737;
  reg [31:0] _RAND_2738;
  reg [31:0] _RAND_2739;
  reg [31:0] _RAND_2740;
  reg [31:0] _RAND_2741;
  reg [31:0] _RAND_2742;
  reg [31:0] _RAND_2743;
  reg [31:0] _RAND_2744;
  reg [31:0] _RAND_2745;
  reg [31:0] _RAND_2746;
  reg [31:0] _RAND_2747;
  reg [31:0] _RAND_2748;
  reg [31:0] _RAND_2749;
  reg [31:0] _RAND_2750;
  reg [31:0] _RAND_2751;
  reg [31:0] _RAND_2752;
  reg [31:0] _RAND_2753;
  reg [31:0] _RAND_2754;
  reg [31:0] _RAND_2755;
  reg [31:0] _RAND_2756;
  reg [31:0] _RAND_2757;
  reg [31:0] _RAND_2758;
  reg [31:0] _RAND_2759;
  reg [31:0] _RAND_2760;
  reg [31:0] _RAND_2761;
  reg [31:0] _RAND_2762;
  reg [31:0] _RAND_2763;
  reg [31:0] _RAND_2764;
  reg [31:0] _RAND_2765;
  reg [31:0] _RAND_2766;
  reg [31:0] _RAND_2767;
  reg [31:0] _RAND_2768;
  reg [31:0] _RAND_2769;
  reg [31:0] _RAND_2770;
  reg [31:0] _RAND_2771;
  reg [31:0] _RAND_2772;
  reg [31:0] _RAND_2773;
  reg [31:0] _RAND_2774;
  reg [31:0] _RAND_2775;
  reg [31:0] _RAND_2776;
  reg [31:0] _RAND_2777;
  reg [31:0] _RAND_2778;
  reg [31:0] _RAND_2779;
  reg [31:0] _RAND_2780;
  reg [31:0] _RAND_2781;
  reg [31:0] _RAND_2782;
  reg [31:0] _RAND_2783;
  reg [31:0] _RAND_2784;
  reg [31:0] _RAND_2785;
  reg [31:0] _RAND_2786;
  reg [31:0] _RAND_2787;
  reg [31:0] _RAND_2788;
  reg [31:0] _RAND_2789;
  reg [31:0] _RAND_2790;
  reg [31:0] _RAND_2791;
  reg [31:0] _RAND_2792;
  reg [31:0] _RAND_2793;
  reg [31:0] _RAND_2794;
  reg [31:0] _RAND_2795;
  reg [31:0] _RAND_2796;
  reg [31:0] _RAND_2797;
  reg [31:0] _RAND_2798;
  reg [31:0] _RAND_2799;
  reg [31:0] _RAND_2800;
  reg [31:0] _RAND_2801;
  reg [31:0] _RAND_2802;
  reg [31:0] _RAND_2803;
  reg [31:0] _RAND_2804;
  reg [31:0] _RAND_2805;
  reg [31:0] _RAND_2806;
  reg [31:0] _RAND_2807;
  reg [31:0] _RAND_2808;
  reg [31:0] _RAND_2809;
  reg [31:0] _RAND_2810;
  reg [31:0] _RAND_2811;
  reg [31:0] _RAND_2812;
  reg [31:0] _RAND_2813;
  reg [31:0] _RAND_2814;
  reg [31:0] _RAND_2815;
  reg [31:0] _RAND_2816;
  reg [31:0] _RAND_2817;
  reg [31:0] _RAND_2818;
  reg [31:0] _RAND_2819;
  reg [31:0] _RAND_2820;
  reg [31:0] _RAND_2821;
  reg [31:0] _RAND_2822;
  reg [31:0] _RAND_2823;
  reg [31:0] _RAND_2824;
  reg [31:0] _RAND_2825;
  reg [31:0] _RAND_2826;
  reg [31:0] _RAND_2827;
  reg [31:0] _RAND_2828;
  reg [31:0] _RAND_2829;
  reg [31:0] _RAND_2830;
  reg [31:0] _RAND_2831;
  reg [31:0] _RAND_2832;
  reg [31:0] _RAND_2833;
  reg [31:0] _RAND_2834;
  reg [31:0] _RAND_2835;
  reg [31:0] _RAND_2836;
  reg [31:0] _RAND_2837;
  reg [31:0] _RAND_2838;
  reg [31:0] _RAND_2839;
  reg [31:0] _RAND_2840;
  reg [31:0] _RAND_2841;
  reg [31:0] _RAND_2842;
  reg [31:0] _RAND_2843;
  reg [31:0] _RAND_2844;
  reg [31:0] _RAND_2845;
  reg [31:0] _RAND_2846;
  reg [31:0] _RAND_2847;
  reg [31:0] _RAND_2848;
  reg [31:0] _RAND_2849;
  reg [31:0] _RAND_2850;
  reg [31:0] _RAND_2851;
  reg [31:0] _RAND_2852;
  reg [31:0] _RAND_2853;
  reg [31:0] _RAND_2854;
  reg [31:0] _RAND_2855;
  reg [31:0] _RAND_2856;
  reg [31:0] _RAND_2857;
  reg [31:0] _RAND_2858;
  reg [31:0] _RAND_2859;
  reg [31:0] _RAND_2860;
  reg [31:0] _RAND_2861;
  reg [31:0] _RAND_2862;
  reg [31:0] _RAND_2863;
  reg [31:0] _RAND_2864;
  reg [31:0] _RAND_2865;
  reg [31:0] _RAND_2866;
  reg [31:0] _RAND_2867;
  reg [31:0] _RAND_2868;
  reg [31:0] _RAND_2869;
  reg [31:0] _RAND_2870;
  reg [31:0] _RAND_2871;
  reg [31:0] _RAND_2872;
  reg [31:0] _RAND_2873;
  reg [31:0] _RAND_2874;
  reg [31:0] _RAND_2875;
  reg [31:0] _RAND_2876;
  reg [31:0] _RAND_2877;
  reg [31:0] _RAND_2878;
  reg [31:0] _RAND_2879;
  reg [31:0] _RAND_2880;
  reg [31:0] _RAND_2881;
  reg [31:0] _RAND_2882;
  reg [31:0] _RAND_2883;
  reg [31:0] _RAND_2884;
  reg [31:0] _RAND_2885;
  reg [31:0] _RAND_2886;
  reg [31:0] _RAND_2887;
  reg [31:0] _RAND_2888;
  reg [31:0] _RAND_2889;
  reg [31:0] _RAND_2890;
  reg [31:0] _RAND_2891;
  reg [31:0] _RAND_2892;
  reg [31:0] _RAND_2893;
  reg [31:0] _RAND_2894;
  reg [31:0] _RAND_2895;
  reg [31:0] _RAND_2896;
  reg [31:0] _RAND_2897;
  reg [31:0] _RAND_2898;
  reg [31:0] _RAND_2899;
  reg [31:0] _RAND_2900;
  reg [31:0] _RAND_2901;
  reg [31:0] _RAND_2902;
  reg [31:0] _RAND_2903;
  reg [31:0] _RAND_2904;
  reg [31:0] _RAND_2905;
  reg [31:0] _RAND_2906;
  reg [31:0] _RAND_2907;
  reg [31:0] _RAND_2908;
  reg [31:0] _RAND_2909;
  reg [31:0] _RAND_2910;
  reg [31:0] _RAND_2911;
  reg [31:0] _RAND_2912;
  reg [31:0] _RAND_2913;
  reg [31:0] _RAND_2914;
  reg [31:0] _RAND_2915;
  reg [31:0] _RAND_2916;
  reg [31:0] _RAND_2917;
  reg [31:0] _RAND_2918;
  reg [31:0] _RAND_2919;
  reg [31:0] _RAND_2920;
  reg [31:0] _RAND_2921;
  reg [31:0] _RAND_2922;
  reg [31:0] _RAND_2923;
  reg [31:0] _RAND_2924;
  reg [31:0] _RAND_2925;
  reg [31:0] _RAND_2926;
  reg [31:0] _RAND_2927;
  reg [31:0] _RAND_2928;
  reg [31:0] _RAND_2929;
  reg [31:0] _RAND_2930;
  reg [31:0] _RAND_2931;
  reg [31:0] _RAND_2932;
  reg [31:0] _RAND_2933;
  reg [31:0] _RAND_2934;
  reg [31:0] _RAND_2935;
  reg [31:0] _RAND_2936;
  reg [31:0] _RAND_2937;
  reg [31:0] _RAND_2938;
  reg [31:0] _RAND_2939;
  reg [31:0] _RAND_2940;
  reg [31:0] _RAND_2941;
  reg [31:0] _RAND_2942;
  reg [31:0] _RAND_2943;
  reg [31:0] _RAND_2944;
  reg [31:0] _RAND_2945;
  reg [31:0] _RAND_2946;
  reg [31:0] _RAND_2947;
  reg [31:0] _RAND_2948;
  reg [31:0] _RAND_2949;
  reg [31:0] _RAND_2950;
  reg [31:0] _RAND_2951;
  reg [31:0] _RAND_2952;
  reg [31:0] _RAND_2953;
  reg [31:0] _RAND_2954;
  reg [31:0] _RAND_2955;
  reg [31:0] _RAND_2956;
  reg [31:0] _RAND_2957;
  reg [31:0] _RAND_2958;
  reg [31:0] _RAND_2959;
  reg [31:0] _RAND_2960;
  reg [31:0] _RAND_2961;
  reg [31:0] _RAND_2962;
  reg [31:0] _RAND_2963;
  reg [31:0] _RAND_2964;
  reg [31:0] _RAND_2965;
  reg [31:0] _RAND_2966;
  reg [31:0] _RAND_2967;
  reg [31:0] _RAND_2968;
  reg [31:0] _RAND_2969;
  reg [31:0] _RAND_2970;
  reg [31:0] _RAND_2971;
  reg [31:0] _RAND_2972;
  reg [31:0] _RAND_2973;
  reg [31:0] _RAND_2974;
  reg [31:0] _RAND_2975;
  reg [31:0] _RAND_2976;
  reg [31:0] _RAND_2977;
  reg [31:0] _RAND_2978;
  reg [31:0] _RAND_2979;
  reg [31:0] _RAND_2980;
  reg [31:0] _RAND_2981;
  reg [31:0] _RAND_2982;
  reg [31:0] _RAND_2983;
  reg [31:0] _RAND_2984;
  reg [31:0] _RAND_2985;
  reg [31:0] _RAND_2986;
  reg [31:0] _RAND_2987;
  reg [31:0] _RAND_2988;
  reg [31:0] _RAND_2989;
  reg [31:0] _RAND_2990;
  reg [31:0] _RAND_2991;
  reg [31:0] _RAND_2992;
  reg [31:0] _RAND_2993;
  reg [31:0] _RAND_2994;
  reg [31:0] _RAND_2995;
  reg [31:0] _RAND_2996;
  reg [31:0] _RAND_2997;
  reg [31:0] _RAND_2998;
  reg [31:0] _RAND_2999;
  reg [31:0] _RAND_3000;
  reg [31:0] _RAND_3001;
  reg [31:0] _RAND_3002;
  reg [31:0] _RAND_3003;
  reg [31:0] _RAND_3004;
  reg [31:0] _RAND_3005;
  reg [31:0] _RAND_3006;
  reg [31:0] _RAND_3007;
  reg [31:0] _RAND_3008;
  reg [31:0] _RAND_3009;
  reg [31:0] _RAND_3010;
  reg [31:0] _RAND_3011;
  reg [31:0] _RAND_3012;
  reg [31:0] _RAND_3013;
  reg [31:0] _RAND_3014;
  reg [31:0] _RAND_3015;
  reg [31:0] _RAND_3016;
  reg [31:0] _RAND_3017;
  reg [31:0] _RAND_3018;
  reg [31:0] _RAND_3019;
  reg [31:0] _RAND_3020;
  reg [31:0] _RAND_3021;
  reg [31:0] _RAND_3022;
  reg [31:0] _RAND_3023;
  reg [31:0] _RAND_3024;
  reg [31:0] _RAND_3025;
  reg [31:0] _RAND_3026;
  reg [31:0] _RAND_3027;
  reg [31:0] _RAND_3028;
  reg [31:0] _RAND_3029;
  reg [31:0] _RAND_3030;
  reg [31:0] _RAND_3031;
  reg [31:0] _RAND_3032;
  reg [31:0] _RAND_3033;
  reg [31:0] _RAND_3034;
  reg [31:0] _RAND_3035;
  reg [31:0] _RAND_3036;
  reg [31:0] _RAND_3037;
  reg [31:0] _RAND_3038;
  reg [31:0] _RAND_3039;
  reg [31:0] _RAND_3040;
  reg [31:0] _RAND_3041;
  reg [31:0] _RAND_3042;
  reg [31:0] _RAND_3043;
  reg [31:0] _RAND_3044;
  reg [31:0] _RAND_3045;
  reg [31:0] _RAND_3046;
  reg [31:0] _RAND_3047;
  reg [31:0] _RAND_3048;
  reg [31:0] _RAND_3049;
  reg [31:0] _RAND_3050;
  reg [31:0] _RAND_3051;
  reg [31:0] _RAND_3052;
  reg [31:0] _RAND_3053;
  reg [31:0] _RAND_3054;
  reg [31:0] _RAND_3055;
  reg [31:0] _RAND_3056;
  reg [31:0] _RAND_3057;
  reg [31:0] _RAND_3058;
  reg [31:0] _RAND_3059;
  reg [31:0] _RAND_3060;
  reg [31:0] _RAND_3061;
  reg [31:0] _RAND_3062;
  reg [31:0] _RAND_3063;
  reg [31:0] _RAND_3064;
  reg [31:0] _RAND_3065;
  reg [31:0] _RAND_3066;
  reg [31:0] _RAND_3067;
  reg [31:0] _RAND_3068;
  reg [31:0] _RAND_3069;
  reg [31:0] _RAND_3070;
  reg [31:0] _RAND_3071;
  reg [31:0] _RAND_3072;
  reg [31:0] _RAND_3073;
  reg [31:0] _RAND_3074;
  reg [31:0] _RAND_3075;
  reg [31:0] _RAND_3076;
  reg [31:0] _RAND_3077;
  reg [31:0] _RAND_3078;
  reg [31:0] _RAND_3079;
  reg [31:0] _RAND_3080;
  reg [31:0] _RAND_3081;
  reg [31:0] _RAND_3082;
  reg [31:0] _RAND_3083;
  reg [31:0] _RAND_3084;
  reg [31:0] _RAND_3085;
  reg [31:0] _RAND_3086;
  reg [31:0] _RAND_3087;
  reg [31:0] _RAND_3088;
  reg [31:0] _RAND_3089;
  reg [31:0] _RAND_3090;
  reg [31:0] _RAND_3091;
  reg [31:0] _RAND_3092;
  reg [31:0] _RAND_3093;
  reg [31:0] _RAND_3094;
  reg [31:0] _RAND_3095;
  reg [31:0] _RAND_3096;
  reg [31:0] _RAND_3097;
  reg [31:0] _RAND_3098;
  reg [31:0] _RAND_3099;
  reg [31:0] _RAND_3100;
  reg [31:0] _RAND_3101;
  reg [31:0] _RAND_3102;
  reg [31:0] _RAND_3103;
  reg [31:0] _RAND_3104;
  reg [31:0] _RAND_3105;
  reg [31:0] _RAND_3106;
  reg [31:0] _RAND_3107;
  reg [31:0] _RAND_3108;
  reg [31:0] _RAND_3109;
  reg [31:0] _RAND_3110;
  reg [31:0] _RAND_3111;
  reg [31:0] _RAND_3112;
  reg [31:0] _RAND_3113;
  reg [31:0] _RAND_3114;
  reg [31:0] _RAND_3115;
  reg [31:0] _RAND_3116;
  reg [31:0] _RAND_3117;
  reg [31:0] _RAND_3118;
  reg [31:0] _RAND_3119;
  reg [31:0] _RAND_3120;
  reg [31:0] _RAND_3121;
  reg [31:0] _RAND_3122;
  reg [31:0] _RAND_3123;
  reg [31:0] _RAND_3124;
  reg [31:0] _RAND_3125;
  reg [31:0] _RAND_3126;
  reg [31:0] _RAND_3127;
  reg [31:0] _RAND_3128;
  reg [31:0] _RAND_3129;
  reg [31:0] _RAND_3130;
  reg [31:0] _RAND_3131;
  reg [31:0] _RAND_3132;
  reg [31:0] _RAND_3133;
  reg [31:0] _RAND_3134;
  reg [31:0] _RAND_3135;
  reg [31:0] _RAND_3136;
  reg [31:0] _RAND_3137;
  reg [31:0] _RAND_3138;
  reg [31:0] _RAND_3139;
  reg [31:0] _RAND_3140;
  reg [31:0] _RAND_3141;
  reg [31:0] _RAND_3142;
  reg [31:0] _RAND_3143;
  reg [31:0] _RAND_3144;
  reg [31:0] _RAND_3145;
  reg [31:0] _RAND_3146;
  reg [31:0] _RAND_3147;
  reg [31:0] _RAND_3148;
  reg [31:0] _RAND_3149;
  reg [31:0] _RAND_3150;
  reg [31:0] _RAND_3151;
  reg [31:0] _RAND_3152;
  reg [31:0] _RAND_3153;
  reg [31:0] _RAND_3154;
  reg [31:0] _RAND_3155;
  reg [31:0] _RAND_3156;
  reg [31:0] _RAND_3157;
  reg [31:0] _RAND_3158;
  reg [31:0] _RAND_3159;
  reg [31:0] _RAND_3160;
  reg [31:0] _RAND_3161;
  reg [31:0] _RAND_3162;
  reg [31:0] _RAND_3163;
  reg [31:0] _RAND_3164;
  reg [31:0] _RAND_3165;
  reg [31:0] _RAND_3166;
  reg [31:0] _RAND_3167;
  reg [31:0] _RAND_3168;
  reg [31:0] _RAND_3169;
  reg [31:0] _RAND_3170;
  reg [31:0] _RAND_3171;
  reg [31:0] _RAND_3172;
  reg [31:0] _RAND_3173;
  reg [31:0] _RAND_3174;
  reg [31:0] _RAND_3175;
  reg [31:0] _RAND_3176;
  reg [31:0] _RAND_3177;
  reg [31:0] _RAND_3178;
  reg [31:0] _RAND_3179;
  reg [31:0] _RAND_3180;
  reg [31:0] _RAND_3181;
  reg [31:0] _RAND_3182;
  reg [31:0] _RAND_3183;
  reg [31:0] _RAND_3184;
  reg [31:0] _RAND_3185;
  reg [31:0] _RAND_3186;
  reg [31:0] _RAND_3187;
  reg [31:0] _RAND_3188;
  reg [31:0] _RAND_3189;
  reg [31:0] _RAND_3190;
  reg [31:0] _RAND_3191;
  reg [31:0] _RAND_3192;
  reg [31:0] _RAND_3193;
  reg [31:0] _RAND_3194;
  reg [31:0] _RAND_3195;
  reg [31:0] _RAND_3196;
  reg [31:0] _RAND_3197;
  reg [31:0] _RAND_3198;
  reg [31:0] _RAND_3199;
  reg [31:0] _RAND_3200;
  reg [31:0] _RAND_3201;
  reg [31:0] _RAND_3202;
  reg [31:0] _RAND_3203;
  reg [31:0] _RAND_3204;
  reg [31:0] _RAND_3205;
  reg [31:0] _RAND_3206;
  reg [31:0] _RAND_3207;
  reg [31:0] _RAND_3208;
  reg [31:0] _RAND_3209;
  reg [31:0] _RAND_3210;
  reg [31:0] _RAND_3211;
  reg [31:0] _RAND_3212;
  reg [31:0] _RAND_3213;
  reg [31:0] _RAND_3214;
  reg [31:0] _RAND_3215;
  reg [31:0] _RAND_3216;
  reg [31:0] _RAND_3217;
  reg [31:0] _RAND_3218;
  reg [31:0] _RAND_3219;
  reg [31:0] _RAND_3220;
  reg [31:0] _RAND_3221;
  reg [31:0] _RAND_3222;
  reg [31:0] _RAND_3223;
  reg [31:0] _RAND_3224;
  reg [31:0] _RAND_3225;
  reg [31:0] _RAND_3226;
  reg [31:0] _RAND_3227;
  reg [31:0] _RAND_3228;
  reg [31:0] _RAND_3229;
  reg [31:0] _RAND_3230;
  reg [31:0] _RAND_3231;
  reg [31:0] _RAND_3232;
  reg [31:0] _RAND_3233;
  reg [31:0] _RAND_3234;
  reg [31:0] _RAND_3235;
  reg [31:0] _RAND_3236;
  reg [31:0] _RAND_3237;
  reg [31:0] _RAND_3238;
  reg [31:0] _RAND_3239;
  reg [31:0] _RAND_3240;
  reg [31:0] _RAND_3241;
  reg [31:0] _RAND_3242;
  reg [31:0] _RAND_3243;
  reg [31:0] _RAND_3244;
  reg [31:0] _RAND_3245;
  reg [31:0] _RAND_3246;
  reg [31:0] _RAND_3247;
  reg [31:0] _RAND_3248;
  reg [31:0] _RAND_3249;
  reg [31:0] _RAND_3250;
  reg [31:0] _RAND_3251;
  reg [31:0] _RAND_3252;
  reg [31:0] _RAND_3253;
  reg [31:0] _RAND_3254;
  reg [31:0] _RAND_3255;
  reg [31:0] _RAND_3256;
  reg [31:0] _RAND_3257;
  reg [31:0] _RAND_3258;
  reg [31:0] _RAND_3259;
  reg [31:0] _RAND_3260;
  reg [31:0] _RAND_3261;
  reg [31:0] _RAND_3262;
  reg [31:0] _RAND_3263;
  reg [31:0] _RAND_3264;
  reg [31:0] _RAND_3265;
  reg [31:0] _RAND_3266;
  reg [31:0] _RAND_3267;
  reg [31:0] _RAND_3268;
  reg [31:0] _RAND_3269;
  reg [31:0] _RAND_3270;
  reg [31:0] _RAND_3271;
  reg [31:0] _RAND_3272;
  reg [31:0] _RAND_3273;
  reg [31:0] _RAND_3274;
  reg [31:0] _RAND_3275;
  reg [31:0] _RAND_3276;
  reg [31:0] _RAND_3277;
  reg [31:0] _RAND_3278;
  reg [31:0] _RAND_3279;
  reg [31:0] _RAND_3280;
  reg [31:0] _RAND_3281;
  reg [31:0] _RAND_3282;
  reg [31:0] _RAND_3283;
  reg [31:0] _RAND_3284;
  reg [31:0] _RAND_3285;
  reg [31:0] _RAND_3286;
  reg [31:0] _RAND_3287;
  reg [31:0] _RAND_3288;
  reg [31:0] _RAND_3289;
  reg [31:0] _RAND_3290;
  reg [31:0] _RAND_3291;
  reg [31:0] _RAND_3292;
  reg [31:0] _RAND_3293;
  reg [31:0] _RAND_3294;
  reg [31:0] _RAND_3295;
  reg [31:0] _RAND_3296;
  reg [31:0] _RAND_3297;
  reg [31:0] _RAND_3298;
  reg [31:0] _RAND_3299;
  reg [31:0] _RAND_3300;
  reg [31:0] _RAND_3301;
  reg [31:0] _RAND_3302;
  reg [31:0] _RAND_3303;
  reg [31:0] _RAND_3304;
  reg [31:0] _RAND_3305;
  reg [31:0] _RAND_3306;
  reg [31:0] _RAND_3307;
  reg [31:0] _RAND_3308;
  reg [31:0] _RAND_3309;
  reg [31:0] _RAND_3310;
  reg [31:0] _RAND_3311;
  reg [31:0] _RAND_3312;
  reg [31:0] _RAND_3313;
  reg [31:0] _RAND_3314;
  reg [31:0] _RAND_3315;
  reg [31:0] _RAND_3316;
  reg [31:0] _RAND_3317;
  reg [31:0] _RAND_3318;
  reg [31:0] _RAND_3319;
  reg [31:0] _RAND_3320;
  reg [31:0] _RAND_3321;
  reg [31:0] _RAND_3322;
  reg [31:0] _RAND_3323;
  reg [31:0] _RAND_3324;
  reg [31:0] _RAND_3325;
  reg [31:0] _RAND_3326;
  reg [31:0] _RAND_3327;
  reg [31:0] _RAND_3328;
  reg [31:0] _RAND_3329;
  reg [31:0] _RAND_3330;
  reg [31:0] _RAND_3331;
  reg [31:0] _RAND_3332;
  reg [31:0] _RAND_3333;
  reg [31:0] _RAND_3334;
  reg [31:0] _RAND_3335;
  reg [31:0] _RAND_3336;
  reg [31:0] _RAND_3337;
  reg [31:0] _RAND_3338;
  reg [31:0] _RAND_3339;
  reg [31:0] _RAND_3340;
  reg [31:0] _RAND_3341;
  reg [31:0] _RAND_3342;
  reg [31:0] _RAND_3343;
  reg [31:0] _RAND_3344;
  reg [31:0] _RAND_3345;
  reg [31:0] _RAND_3346;
  reg [31:0] _RAND_3347;
  reg [31:0] _RAND_3348;
  reg [31:0] _RAND_3349;
`endif // RANDOMIZE_REG_INIT
  wire  proc_0_clock; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_0; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_1; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_2; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_3; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_4; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_5; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_6; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_7; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_8; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_9; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_10; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_11; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_12; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_13; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_14; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_15; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_16; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_17; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_18; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_19; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_20; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_21; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_22; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_23; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_24; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_25; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_26; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_27; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_28; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_29; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_30; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_31; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_32; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_33; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_34; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_35; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_36; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_37; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_38; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_39; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_40; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_41; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_42; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_43; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_44; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_45; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_46; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_47; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_48; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_49; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_50; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_51; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_52; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_53; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_54; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_55; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_56; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_57; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_58; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_59; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_60; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_61; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_62; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_63; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_64; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_65; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_66; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_67; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_68; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_69; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_70; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_71; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_72; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_73; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_74; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_75; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_76; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_77; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_78; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_79; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_80; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_81; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_82; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_83; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_84; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_85; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_86; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_87; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_88; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_89; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_90; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_91; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_92; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_93; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_94; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_95; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_96; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_97; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_98; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_99; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_100; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_101; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_102; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_103; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_104; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_105; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_106; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_107; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_108; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_109; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_110; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_111; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_112; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_113; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_114; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_115; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_116; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_117; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_118; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_119; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_120; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_121; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_122; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_123; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_124; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_125; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_126; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_127; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_128; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_129; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_130; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_131; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_132; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_133; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_134; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_135; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_136; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_137; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_138; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_139; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_140; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_141; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_142; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_143; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_144; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_145; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_146; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_147; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_148; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_149; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_150; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_151; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_152; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_153; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_154; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_155; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_156; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_157; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_158; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_159; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_160; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_161; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_162; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_163; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_164; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_165; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_166; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_167; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_168; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_169; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_170; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_171; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_172; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_173; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_174; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_175; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_176; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_177; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_178; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_179; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_180; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_181; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_182; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_183; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_184; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_185; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_186; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_187; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_188; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_189; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_190; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_191; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_192; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_193; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_194; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_195; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_196; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_197; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_198; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_199; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_200; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_201; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_202; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_203; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_204; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_205; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_206; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_207; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_208; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_209; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_210; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_211; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_212; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_213; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_214; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_215; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_216; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_217; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_218; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_219; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_220; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_221; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_222; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_223; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_224; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_225; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_226; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_227; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_228; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_229; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_230; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_231; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_232; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_233; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_234; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_235; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_236; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_237; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_238; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_239; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_240; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_241; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_242; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_243; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_244; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_245; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_246; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_247; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_248; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_249; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_250; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_251; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_252; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_253; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_254; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_255; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_0; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_1; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_2; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_3; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_4; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_5; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_6; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_7; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_8; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_9; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_10; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_11; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_12; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_13; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_14; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_in_header_15; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 62:25]
  wire [1:0] proc_0_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 62:25]
  wire  proc_0_io_pipe_phv_in_next_config_id; // @[ipsa.scala 62:25]
  wire  proc_0_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_0; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_1; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_2; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_3; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_4; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_5; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_6; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_7; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_8; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_9; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_10; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_11; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_12; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_13; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_14; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_15; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_16; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_17; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_18; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_19; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_20; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_21; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_22; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_23; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_24; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_25; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_26; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_27; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_28; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_29; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_30; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_31; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_32; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_33; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_34; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_35; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_36; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_37; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_38; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_39; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_40; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_41; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_42; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_43; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_44; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_45; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_46; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_47; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_48; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_49; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_50; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_51; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_52; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_53; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_54; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_55; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_56; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_57; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_58; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_59; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_60; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_61; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_62; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_63; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_64; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_65; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_66; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_67; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_68; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_69; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_70; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_71; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_72; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_73; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_74; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_75; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_76; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_77; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_78; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_79; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_80; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_81; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_82; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_83; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_84; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_85; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_86; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_87; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_88; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_89; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_90; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_91; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_92; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_93; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_94; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_95; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_96; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_97; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_98; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_99; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_100; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_101; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_102; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_103; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_104; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_105; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_106; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_107; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_108; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_109; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_110; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_111; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_112; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_113; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_114; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_115; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_116; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_117; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_118; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_119; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_120; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_121; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_122; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_123; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_124; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_125; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_126; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_127; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_128; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_129; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_130; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_131; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_132; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_133; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_134; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_135; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_136; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_137; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_138; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_139; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_140; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_141; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_142; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_143; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_144; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_145; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_146; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_147; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_148; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_149; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_150; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_151; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_152; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_153; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_154; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_155; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_156; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_157; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_158; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_159; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_160; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_161; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_162; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_163; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_164; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_165; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_166; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_167; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_168; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_169; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_170; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_171; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_172; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_173; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_174; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_175; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_176; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_177; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_178; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_179; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_180; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_181; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_182; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_183; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_184; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_185; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_186; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_187; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_188; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_189; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_190; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_191; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_192; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_193; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_194; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_195; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_196; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_197; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_198; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_199; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_200; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_201; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_202; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_203; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_204; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_205; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_206; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_207; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_208; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_209; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_210; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_211; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_212; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_213; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_214; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_215; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_216; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_217; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_218; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_219; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_220; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_221; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_222; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_223; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_224; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_225; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_226; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_227; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_228; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_229; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_230; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_231; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_232; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_233; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_234; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_235; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_236; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_237; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_238; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_239; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_240; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_241; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_242; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_243; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_244; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_245; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_246; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_247; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_248; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_249; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_250; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_251; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_252; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_253; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_254; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_255; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_0; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_1; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_2; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_3; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_4; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_5; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_6; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_7; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_8; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_9; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_10; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_11; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_12; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_13; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_14; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_out_header_15; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 62:25]
  wire [15:0] proc_0_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 62:25]
  wire [1:0] proc_0_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 62:25]
  wire  proc_0_io_pipe_phv_out_next_config_id; // @[ipsa.scala 62:25]
  wire  proc_0_io_mod_par_mod_en; // @[ipsa.scala 62:25]
  wire  proc_0_io_mod_par_mod_last_mau_id_mod; // @[ipsa.scala 62:25]
  wire [1:0] proc_0_io_mod_par_mod_last_mau_id; // @[ipsa.scala 62:25]
  wire [1:0] proc_0_io_mod_par_mod_cs; // @[ipsa.scala 62:25]
  wire  proc_0_io_mod_par_mod_module_mod_state_id_mod; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mod_par_mod_module_mod_state_id; // @[ipsa.scala 62:25]
  wire  proc_0_io_mod_par_mod_module_mod_sram_w_cs; // @[ipsa.scala 62:25]
  wire  proc_0_io_mod_par_mod_module_mod_sram_w_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mod_par_mod_module_mod_sram_w_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mod_par_mod_module_mod_sram_w_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mod_mat_mod_en; // @[ipsa.scala 62:25]
  wire  proc_0_io_mod_mat_mod_config_id; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mod_mat_mod_key_mod_header_id; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mod_mat_mod_key_mod_internal_offset; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mod_mat_mod_key_mod_key_length; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_0; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_1; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_2; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_3; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_4; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_5; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_6; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_7; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_8; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_9; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_10; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_11; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_12; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_13; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_14; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_15; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_16; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_17; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_18; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_19; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_20; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_21; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_22; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_23; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_24; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_25; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_26; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_27; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_28; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_29; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_30; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_31; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_32; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_33; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_34; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_35; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_36; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_37; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_38; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_39; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_40; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_41; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_42; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_43; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_44; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_45; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_46; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_47; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_48; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_49; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_50; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_51; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_52; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_53; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_54; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_55; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_56; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_57; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_58; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_59; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_60; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_61; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_62; // @[ipsa.scala 62:25]
  wire [5:0] proc_0_io_mod_mat_mod_table_mod_sram_id_table_63; // @[ipsa.scala 62:25]
  wire [6:0] proc_0_io_mod_mat_mod_table_mod_table_width; // @[ipsa.scala 62:25]
  wire [6:0] proc_0_io_mod_mat_mod_table_mod_table_depth; // @[ipsa.scala 62:25]
  wire  proc_0_io_mod_act_mod_en_0; // @[ipsa.scala 62:25]
  wire  proc_0_io_mod_act_mod_en_1; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mod_act_mod_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mod_act_mod_data_0; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mod_act_mod_data_1; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_0_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_0_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_0_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_1_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_1_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_1_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_2_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_2_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_2_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_3_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_3_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_3_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_4_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_4_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_4_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_5_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_5_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_5_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_6_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_6_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_6_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_7_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_7_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_7_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_8_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_8_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_8_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_9_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_9_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_9_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_10_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_10_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_10_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_11_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_11_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_11_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_12_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_12_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_12_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_13_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_13_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_13_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_14_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_14_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_14_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_15_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_15_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_15_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_16_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_16_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_16_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_17_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_17_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_17_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_18_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_18_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_18_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_19_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_19_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_19_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_20_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_20_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_20_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_21_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_21_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_21_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_22_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_22_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_22_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_23_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_23_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_23_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_24_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_24_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_24_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_25_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_25_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_25_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_26_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_26_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_26_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_27_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_27_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_27_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_28_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_28_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_28_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_29_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_29_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_29_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_30_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_30_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_30_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_31_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_31_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_31_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_32_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_32_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_32_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_33_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_33_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_33_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_34_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_34_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_34_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_35_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_35_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_35_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_36_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_36_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_36_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_37_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_37_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_37_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_38_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_38_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_38_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_39_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_39_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_39_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_40_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_40_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_40_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_41_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_41_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_41_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_42_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_42_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_42_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_43_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_43_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_43_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_44_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_44_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_44_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_45_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_45_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_45_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_46_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_46_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_46_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_47_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_47_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_47_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_48_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_48_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_48_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_49_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_49_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_49_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_50_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_50_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_50_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_51_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_51_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_51_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_52_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_52_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_52_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_53_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_53_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_53_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_54_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_54_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_54_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_55_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_55_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_55_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_56_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_56_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_56_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_57_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_57_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_57_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_58_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_58_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_58_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_59_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_59_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_59_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_60_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_60_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_60_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_61_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_61_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_61_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_62_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_62_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_62_data; // @[ipsa.scala 62:25]
  wire  proc_0_io_mem_cluster_63_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_0_io_mem_cluster_63_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_0_io_mem_cluster_63_data; // @[ipsa.scala 62:25]
  wire  proc_1_clock; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_0; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_1; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_2; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_3; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_4; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_5; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_6; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_7; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_8; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_9; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_10; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_11; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_12; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_13; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_14; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_15; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_16; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_17; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_18; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_19; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_20; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_21; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_22; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_23; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_24; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_25; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_26; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_27; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_28; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_29; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_30; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_31; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_32; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_33; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_34; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_35; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_36; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_37; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_38; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_39; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_40; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_41; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_42; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_43; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_44; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_45; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_46; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_47; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_48; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_49; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_50; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_51; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_52; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_53; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_54; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_55; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_56; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_57; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_58; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_59; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_60; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_61; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_62; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_63; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_64; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_65; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_66; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_67; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_68; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_69; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_70; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_71; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_72; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_73; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_74; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_75; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_76; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_77; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_78; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_79; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_80; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_81; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_82; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_83; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_84; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_85; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_86; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_87; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_88; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_89; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_90; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_91; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_92; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_93; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_94; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_95; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_96; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_97; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_98; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_99; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_100; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_101; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_102; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_103; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_104; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_105; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_106; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_107; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_108; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_109; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_110; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_111; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_112; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_113; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_114; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_115; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_116; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_117; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_118; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_119; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_120; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_121; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_122; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_123; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_124; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_125; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_126; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_127; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_128; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_129; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_130; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_131; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_132; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_133; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_134; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_135; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_136; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_137; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_138; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_139; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_140; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_141; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_142; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_143; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_144; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_145; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_146; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_147; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_148; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_149; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_150; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_151; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_152; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_153; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_154; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_155; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_156; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_157; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_158; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_159; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_160; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_161; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_162; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_163; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_164; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_165; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_166; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_167; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_168; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_169; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_170; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_171; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_172; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_173; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_174; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_175; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_176; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_177; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_178; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_179; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_180; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_181; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_182; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_183; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_184; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_185; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_186; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_187; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_188; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_189; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_190; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_191; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_192; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_193; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_194; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_195; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_196; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_197; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_198; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_199; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_200; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_201; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_202; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_203; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_204; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_205; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_206; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_207; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_208; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_209; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_210; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_211; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_212; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_213; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_214; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_215; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_216; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_217; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_218; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_219; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_220; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_221; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_222; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_223; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_224; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_225; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_226; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_227; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_228; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_229; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_230; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_231; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_232; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_233; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_234; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_235; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_236; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_237; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_238; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_239; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_240; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_241; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_242; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_243; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_244; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_245; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_246; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_247; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_248; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_249; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_250; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_251; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_252; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_253; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_254; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_255; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_0; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_1; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_2; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_3; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_4; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_5; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_6; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_7; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_8; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_9; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_10; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_11; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_12; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_13; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_14; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_in_header_15; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 62:25]
  wire [1:0] proc_1_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 62:25]
  wire  proc_1_io_pipe_phv_in_next_config_id; // @[ipsa.scala 62:25]
  wire  proc_1_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_0; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_1; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_2; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_3; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_4; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_5; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_6; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_7; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_8; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_9; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_10; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_11; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_12; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_13; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_14; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_15; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_16; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_17; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_18; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_19; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_20; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_21; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_22; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_23; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_24; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_25; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_26; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_27; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_28; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_29; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_30; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_31; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_32; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_33; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_34; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_35; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_36; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_37; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_38; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_39; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_40; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_41; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_42; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_43; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_44; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_45; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_46; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_47; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_48; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_49; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_50; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_51; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_52; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_53; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_54; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_55; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_56; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_57; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_58; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_59; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_60; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_61; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_62; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_63; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_64; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_65; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_66; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_67; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_68; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_69; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_70; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_71; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_72; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_73; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_74; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_75; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_76; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_77; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_78; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_79; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_80; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_81; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_82; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_83; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_84; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_85; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_86; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_87; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_88; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_89; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_90; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_91; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_92; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_93; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_94; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_95; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_96; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_97; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_98; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_99; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_100; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_101; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_102; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_103; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_104; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_105; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_106; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_107; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_108; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_109; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_110; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_111; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_112; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_113; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_114; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_115; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_116; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_117; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_118; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_119; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_120; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_121; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_122; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_123; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_124; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_125; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_126; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_127; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_128; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_129; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_130; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_131; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_132; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_133; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_134; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_135; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_136; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_137; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_138; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_139; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_140; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_141; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_142; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_143; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_144; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_145; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_146; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_147; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_148; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_149; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_150; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_151; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_152; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_153; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_154; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_155; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_156; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_157; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_158; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_159; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_160; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_161; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_162; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_163; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_164; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_165; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_166; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_167; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_168; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_169; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_170; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_171; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_172; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_173; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_174; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_175; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_176; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_177; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_178; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_179; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_180; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_181; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_182; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_183; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_184; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_185; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_186; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_187; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_188; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_189; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_190; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_191; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_192; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_193; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_194; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_195; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_196; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_197; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_198; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_199; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_200; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_201; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_202; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_203; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_204; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_205; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_206; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_207; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_208; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_209; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_210; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_211; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_212; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_213; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_214; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_215; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_216; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_217; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_218; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_219; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_220; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_221; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_222; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_223; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_224; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_225; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_226; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_227; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_228; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_229; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_230; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_231; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_232; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_233; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_234; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_235; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_236; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_237; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_238; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_239; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_240; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_241; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_242; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_243; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_244; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_245; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_246; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_247; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_248; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_249; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_250; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_251; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_252; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_253; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_254; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_255; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_0; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_1; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_2; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_3; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_4; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_5; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_6; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_7; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_8; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_9; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_10; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_11; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_12; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_13; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_14; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_out_header_15; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 62:25]
  wire [15:0] proc_1_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 62:25]
  wire [1:0] proc_1_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 62:25]
  wire  proc_1_io_pipe_phv_out_next_config_id; // @[ipsa.scala 62:25]
  wire  proc_1_io_mod_par_mod_en; // @[ipsa.scala 62:25]
  wire  proc_1_io_mod_par_mod_last_mau_id_mod; // @[ipsa.scala 62:25]
  wire [1:0] proc_1_io_mod_par_mod_last_mau_id; // @[ipsa.scala 62:25]
  wire [1:0] proc_1_io_mod_par_mod_cs; // @[ipsa.scala 62:25]
  wire  proc_1_io_mod_par_mod_module_mod_state_id_mod; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mod_par_mod_module_mod_state_id; // @[ipsa.scala 62:25]
  wire  proc_1_io_mod_par_mod_module_mod_sram_w_cs; // @[ipsa.scala 62:25]
  wire  proc_1_io_mod_par_mod_module_mod_sram_w_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mod_par_mod_module_mod_sram_w_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mod_par_mod_module_mod_sram_w_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mod_mat_mod_en; // @[ipsa.scala 62:25]
  wire  proc_1_io_mod_mat_mod_config_id; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mod_mat_mod_key_mod_header_id; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mod_mat_mod_key_mod_internal_offset; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mod_mat_mod_key_mod_key_length; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_0; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_1; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_2; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_3; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_4; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_5; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_6; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_7; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_8; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_9; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_10; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_11; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_12; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_13; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_14; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_15; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_16; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_17; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_18; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_19; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_20; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_21; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_22; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_23; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_24; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_25; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_26; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_27; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_28; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_29; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_30; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_31; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_32; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_33; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_34; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_35; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_36; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_37; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_38; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_39; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_40; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_41; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_42; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_43; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_44; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_45; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_46; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_47; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_48; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_49; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_50; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_51; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_52; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_53; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_54; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_55; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_56; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_57; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_58; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_59; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_60; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_61; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_62; // @[ipsa.scala 62:25]
  wire [5:0] proc_1_io_mod_mat_mod_table_mod_sram_id_table_63; // @[ipsa.scala 62:25]
  wire [6:0] proc_1_io_mod_mat_mod_table_mod_table_width; // @[ipsa.scala 62:25]
  wire [6:0] proc_1_io_mod_mat_mod_table_mod_table_depth; // @[ipsa.scala 62:25]
  wire  proc_1_io_mod_act_mod_en_0; // @[ipsa.scala 62:25]
  wire  proc_1_io_mod_act_mod_en_1; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mod_act_mod_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mod_act_mod_data_0; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mod_act_mod_data_1; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_0_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_0_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_0_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_1_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_1_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_1_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_2_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_2_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_2_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_3_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_3_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_3_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_4_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_4_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_4_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_5_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_5_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_5_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_6_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_6_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_6_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_7_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_7_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_7_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_8_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_8_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_8_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_9_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_9_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_9_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_10_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_10_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_10_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_11_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_11_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_11_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_12_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_12_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_12_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_13_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_13_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_13_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_14_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_14_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_14_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_15_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_15_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_15_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_16_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_16_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_16_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_17_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_17_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_17_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_18_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_18_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_18_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_19_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_19_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_19_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_20_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_20_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_20_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_21_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_21_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_21_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_22_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_22_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_22_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_23_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_23_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_23_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_24_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_24_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_24_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_25_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_25_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_25_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_26_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_26_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_26_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_27_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_27_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_27_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_28_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_28_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_28_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_29_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_29_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_29_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_30_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_30_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_30_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_31_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_31_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_31_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_32_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_32_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_32_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_33_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_33_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_33_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_34_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_34_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_34_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_35_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_35_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_35_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_36_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_36_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_36_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_37_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_37_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_37_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_38_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_38_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_38_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_39_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_39_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_39_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_40_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_40_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_40_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_41_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_41_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_41_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_42_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_42_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_42_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_43_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_43_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_43_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_44_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_44_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_44_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_45_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_45_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_45_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_46_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_46_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_46_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_47_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_47_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_47_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_48_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_48_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_48_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_49_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_49_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_49_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_50_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_50_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_50_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_51_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_51_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_51_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_52_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_52_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_52_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_53_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_53_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_53_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_54_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_54_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_54_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_55_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_55_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_55_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_56_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_56_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_56_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_57_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_57_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_57_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_58_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_58_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_58_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_59_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_59_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_59_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_60_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_60_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_60_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_61_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_61_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_61_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_62_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_62_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_62_data; // @[ipsa.scala 62:25]
  wire  proc_1_io_mem_cluster_63_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_1_io_mem_cluster_63_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_1_io_mem_cluster_63_data; // @[ipsa.scala 62:25]
  wire  proc_2_clock; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_0; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_1; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_2; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_3; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_4; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_5; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_6; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_7; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_8; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_9; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_10; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_11; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_12; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_13; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_14; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_15; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_16; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_17; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_18; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_19; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_20; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_21; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_22; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_23; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_24; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_25; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_26; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_27; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_28; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_29; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_30; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_31; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_32; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_33; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_34; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_35; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_36; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_37; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_38; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_39; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_40; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_41; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_42; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_43; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_44; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_45; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_46; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_47; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_48; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_49; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_50; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_51; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_52; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_53; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_54; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_55; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_56; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_57; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_58; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_59; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_60; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_61; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_62; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_63; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_64; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_65; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_66; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_67; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_68; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_69; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_70; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_71; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_72; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_73; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_74; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_75; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_76; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_77; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_78; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_79; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_80; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_81; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_82; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_83; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_84; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_85; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_86; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_87; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_88; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_89; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_90; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_91; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_92; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_93; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_94; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_95; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_96; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_97; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_98; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_99; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_100; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_101; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_102; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_103; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_104; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_105; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_106; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_107; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_108; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_109; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_110; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_111; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_112; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_113; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_114; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_115; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_116; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_117; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_118; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_119; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_120; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_121; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_122; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_123; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_124; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_125; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_126; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_127; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_128; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_129; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_130; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_131; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_132; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_133; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_134; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_135; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_136; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_137; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_138; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_139; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_140; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_141; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_142; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_143; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_144; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_145; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_146; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_147; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_148; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_149; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_150; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_151; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_152; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_153; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_154; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_155; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_156; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_157; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_158; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_159; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_160; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_161; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_162; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_163; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_164; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_165; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_166; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_167; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_168; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_169; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_170; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_171; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_172; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_173; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_174; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_175; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_176; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_177; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_178; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_179; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_180; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_181; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_182; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_183; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_184; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_185; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_186; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_187; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_188; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_189; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_190; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_191; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_192; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_193; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_194; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_195; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_196; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_197; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_198; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_199; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_200; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_201; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_202; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_203; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_204; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_205; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_206; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_207; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_208; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_209; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_210; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_211; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_212; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_213; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_214; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_215; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_216; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_217; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_218; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_219; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_220; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_221; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_222; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_223; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_224; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_225; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_226; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_227; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_228; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_229; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_230; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_231; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_232; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_233; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_234; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_235; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_236; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_237; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_238; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_239; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_240; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_241; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_242; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_243; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_244; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_245; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_246; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_247; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_248; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_249; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_250; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_251; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_252; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_253; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_254; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_255; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_0; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_1; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_2; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_3; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_4; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_5; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_6; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_7; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_8; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_9; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_10; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_11; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_12; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_13; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_14; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_in_header_15; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 62:25]
  wire [1:0] proc_2_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 62:25]
  wire  proc_2_io_pipe_phv_in_next_config_id; // @[ipsa.scala 62:25]
  wire  proc_2_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_0; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_1; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_2; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_3; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_4; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_5; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_6; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_7; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_8; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_9; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_10; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_11; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_12; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_13; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_14; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_15; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_16; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_17; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_18; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_19; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_20; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_21; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_22; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_23; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_24; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_25; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_26; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_27; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_28; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_29; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_30; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_31; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_32; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_33; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_34; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_35; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_36; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_37; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_38; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_39; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_40; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_41; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_42; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_43; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_44; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_45; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_46; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_47; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_48; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_49; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_50; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_51; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_52; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_53; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_54; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_55; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_56; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_57; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_58; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_59; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_60; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_61; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_62; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_63; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_64; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_65; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_66; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_67; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_68; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_69; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_70; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_71; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_72; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_73; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_74; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_75; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_76; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_77; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_78; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_79; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_80; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_81; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_82; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_83; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_84; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_85; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_86; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_87; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_88; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_89; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_90; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_91; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_92; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_93; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_94; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_95; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_96; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_97; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_98; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_99; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_100; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_101; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_102; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_103; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_104; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_105; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_106; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_107; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_108; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_109; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_110; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_111; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_112; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_113; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_114; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_115; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_116; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_117; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_118; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_119; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_120; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_121; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_122; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_123; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_124; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_125; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_126; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_127; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_128; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_129; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_130; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_131; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_132; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_133; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_134; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_135; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_136; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_137; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_138; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_139; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_140; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_141; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_142; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_143; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_144; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_145; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_146; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_147; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_148; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_149; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_150; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_151; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_152; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_153; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_154; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_155; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_156; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_157; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_158; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_159; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_160; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_161; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_162; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_163; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_164; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_165; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_166; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_167; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_168; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_169; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_170; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_171; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_172; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_173; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_174; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_175; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_176; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_177; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_178; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_179; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_180; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_181; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_182; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_183; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_184; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_185; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_186; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_187; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_188; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_189; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_190; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_191; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_192; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_193; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_194; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_195; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_196; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_197; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_198; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_199; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_200; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_201; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_202; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_203; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_204; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_205; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_206; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_207; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_208; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_209; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_210; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_211; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_212; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_213; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_214; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_215; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_216; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_217; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_218; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_219; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_220; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_221; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_222; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_223; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_224; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_225; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_226; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_227; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_228; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_229; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_230; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_231; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_232; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_233; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_234; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_235; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_236; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_237; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_238; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_239; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_240; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_241; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_242; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_243; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_244; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_245; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_246; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_247; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_248; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_249; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_250; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_251; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_252; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_253; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_254; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_255; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_0; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_1; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_2; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_3; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_4; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_5; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_6; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_7; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_8; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_9; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_10; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_11; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_12; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_13; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_14; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_out_header_15; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 62:25]
  wire [15:0] proc_2_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 62:25]
  wire [1:0] proc_2_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 62:25]
  wire  proc_2_io_pipe_phv_out_next_config_id; // @[ipsa.scala 62:25]
  wire  proc_2_io_mod_par_mod_en; // @[ipsa.scala 62:25]
  wire  proc_2_io_mod_par_mod_last_mau_id_mod; // @[ipsa.scala 62:25]
  wire [1:0] proc_2_io_mod_par_mod_last_mau_id; // @[ipsa.scala 62:25]
  wire [1:0] proc_2_io_mod_par_mod_cs; // @[ipsa.scala 62:25]
  wire  proc_2_io_mod_par_mod_module_mod_state_id_mod; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mod_par_mod_module_mod_state_id; // @[ipsa.scala 62:25]
  wire  proc_2_io_mod_par_mod_module_mod_sram_w_cs; // @[ipsa.scala 62:25]
  wire  proc_2_io_mod_par_mod_module_mod_sram_w_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mod_par_mod_module_mod_sram_w_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mod_par_mod_module_mod_sram_w_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mod_mat_mod_en; // @[ipsa.scala 62:25]
  wire  proc_2_io_mod_mat_mod_config_id; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mod_mat_mod_key_mod_header_id; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mod_mat_mod_key_mod_internal_offset; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mod_mat_mod_key_mod_key_length; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_0; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_1; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_2; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_3; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_4; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_5; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_6; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_7; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_8; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_9; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_10; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_11; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_12; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_13; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_14; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_15; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_16; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_17; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_18; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_19; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_20; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_21; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_22; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_23; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_24; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_25; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_26; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_27; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_28; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_29; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_30; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_31; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_32; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_33; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_34; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_35; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_36; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_37; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_38; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_39; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_40; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_41; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_42; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_43; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_44; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_45; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_46; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_47; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_48; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_49; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_50; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_51; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_52; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_53; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_54; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_55; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_56; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_57; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_58; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_59; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_60; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_61; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_62; // @[ipsa.scala 62:25]
  wire [5:0] proc_2_io_mod_mat_mod_table_mod_sram_id_table_63; // @[ipsa.scala 62:25]
  wire [6:0] proc_2_io_mod_mat_mod_table_mod_table_width; // @[ipsa.scala 62:25]
  wire [6:0] proc_2_io_mod_mat_mod_table_mod_table_depth; // @[ipsa.scala 62:25]
  wire  proc_2_io_mod_act_mod_en_0; // @[ipsa.scala 62:25]
  wire  proc_2_io_mod_act_mod_en_1; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mod_act_mod_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mod_act_mod_data_0; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mod_act_mod_data_1; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_0_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_0_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_0_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_1_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_1_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_1_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_2_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_2_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_2_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_3_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_3_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_3_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_4_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_4_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_4_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_5_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_5_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_5_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_6_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_6_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_6_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_7_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_7_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_7_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_8_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_8_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_8_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_9_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_9_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_9_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_10_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_10_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_10_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_11_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_11_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_11_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_12_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_12_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_12_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_13_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_13_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_13_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_14_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_14_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_14_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_15_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_15_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_15_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_16_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_16_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_16_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_17_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_17_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_17_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_18_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_18_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_18_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_19_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_19_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_19_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_20_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_20_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_20_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_21_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_21_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_21_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_22_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_22_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_22_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_23_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_23_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_23_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_24_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_24_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_24_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_25_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_25_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_25_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_26_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_26_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_26_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_27_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_27_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_27_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_28_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_28_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_28_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_29_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_29_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_29_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_30_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_30_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_30_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_31_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_31_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_31_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_32_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_32_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_32_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_33_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_33_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_33_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_34_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_34_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_34_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_35_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_35_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_35_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_36_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_36_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_36_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_37_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_37_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_37_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_38_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_38_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_38_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_39_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_39_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_39_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_40_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_40_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_40_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_41_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_41_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_41_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_42_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_42_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_42_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_43_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_43_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_43_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_44_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_44_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_44_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_45_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_45_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_45_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_46_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_46_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_46_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_47_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_47_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_47_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_48_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_48_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_48_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_49_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_49_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_49_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_50_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_50_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_50_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_51_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_51_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_51_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_52_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_52_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_52_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_53_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_53_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_53_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_54_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_54_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_54_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_55_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_55_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_55_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_56_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_56_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_56_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_57_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_57_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_57_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_58_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_58_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_58_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_59_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_59_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_59_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_60_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_60_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_60_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_61_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_61_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_61_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_62_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_62_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_62_data; // @[ipsa.scala 62:25]
  wire  proc_2_io_mem_cluster_63_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_2_io_mem_cluster_63_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_2_io_mem_cluster_63_data; // @[ipsa.scala 62:25]
  wire  proc_3_clock; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_0; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_1; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_2; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_3; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_4; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_5; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_6; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_7; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_8; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_9; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_10; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_11; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_12; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_13; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_14; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_15; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_16; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_17; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_18; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_19; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_20; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_21; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_22; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_23; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_24; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_25; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_26; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_27; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_28; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_29; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_30; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_31; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_32; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_33; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_34; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_35; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_36; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_37; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_38; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_39; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_40; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_41; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_42; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_43; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_44; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_45; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_46; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_47; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_48; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_49; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_50; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_51; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_52; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_53; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_54; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_55; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_56; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_57; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_58; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_59; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_60; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_61; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_62; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_63; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_64; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_65; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_66; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_67; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_68; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_69; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_70; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_71; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_72; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_73; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_74; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_75; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_76; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_77; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_78; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_79; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_80; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_81; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_82; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_83; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_84; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_85; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_86; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_87; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_88; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_89; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_90; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_91; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_92; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_93; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_94; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_95; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_96; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_97; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_98; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_99; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_100; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_101; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_102; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_103; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_104; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_105; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_106; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_107; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_108; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_109; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_110; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_111; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_112; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_113; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_114; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_115; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_116; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_117; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_118; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_119; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_120; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_121; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_122; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_123; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_124; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_125; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_126; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_127; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_128; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_129; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_130; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_131; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_132; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_133; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_134; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_135; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_136; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_137; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_138; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_139; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_140; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_141; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_142; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_143; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_144; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_145; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_146; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_147; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_148; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_149; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_150; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_151; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_152; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_153; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_154; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_155; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_156; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_157; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_158; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_159; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_160; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_161; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_162; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_163; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_164; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_165; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_166; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_167; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_168; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_169; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_170; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_171; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_172; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_173; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_174; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_175; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_176; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_177; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_178; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_179; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_180; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_181; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_182; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_183; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_184; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_185; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_186; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_187; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_188; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_189; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_190; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_191; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_192; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_193; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_194; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_195; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_196; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_197; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_198; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_199; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_200; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_201; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_202; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_203; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_204; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_205; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_206; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_207; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_208; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_209; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_210; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_211; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_212; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_213; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_214; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_215; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_216; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_217; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_218; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_219; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_220; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_221; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_222; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_223; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_224; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_225; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_226; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_227; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_228; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_229; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_230; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_231; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_232; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_233; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_234; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_235; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_236; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_237; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_238; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_239; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_240; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_241; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_242; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_243; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_244; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_245; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_246; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_247; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_248; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_249; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_250; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_251; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_252; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_253; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_254; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_255; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_0; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_1; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_2; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_3; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_4; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_5; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_6; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_7; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_8; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_9; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_10; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_11; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_12; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_13; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_14; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_in_header_15; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 62:25]
  wire [1:0] proc_3_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 62:25]
  wire  proc_3_io_pipe_phv_in_next_config_id; // @[ipsa.scala 62:25]
  wire  proc_3_io_pipe_phv_in_is_valid_processor; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_0; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_1; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_2; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_3; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_4; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_5; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_6; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_7; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_8; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_9; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_10; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_11; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_12; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_13; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_14; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_15; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_16; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_17; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_18; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_19; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_20; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_21; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_22; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_23; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_24; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_25; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_26; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_27; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_28; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_29; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_30; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_31; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_32; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_33; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_34; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_35; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_36; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_37; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_38; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_39; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_40; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_41; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_42; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_43; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_44; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_45; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_46; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_47; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_48; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_49; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_50; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_51; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_52; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_53; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_54; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_55; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_56; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_57; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_58; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_59; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_60; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_61; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_62; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_63; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_64; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_65; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_66; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_67; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_68; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_69; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_70; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_71; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_72; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_73; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_74; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_75; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_76; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_77; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_78; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_79; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_80; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_81; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_82; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_83; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_84; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_85; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_86; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_87; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_88; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_89; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_90; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_91; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_92; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_93; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_94; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_95; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_96; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_97; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_98; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_99; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_100; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_101; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_102; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_103; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_104; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_105; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_106; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_107; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_108; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_109; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_110; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_111; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_112; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_113; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_114; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_115; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_116; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_117; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_118; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_119; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_120; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_121; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_122; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_123; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_124; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_125; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_126; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_127; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_128; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_129; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_130; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_131; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_132; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_133; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_134; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_135; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_136; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_137; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_138; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_139; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_140; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_141; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_142; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_143; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_144; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_145; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_146; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_147; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_148; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_149; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_150; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_151; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_152; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_153; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_154; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_155; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_156; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_157; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_158; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_159; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_160; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_161; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_162; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_163; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_164; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_165; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_166; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_167; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_168; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_169; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_170; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_171; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_172; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_173; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_174; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_175; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_176; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_177; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_178; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_179; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_180; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_181; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_182; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_183; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_184; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_185; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_186; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_187; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_188; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_189; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_190; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_191; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_192; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_193; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_194; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_195; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_196; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_197; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_198; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_199; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_200; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_201; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_202; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_203; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_204; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_205; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_206; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_207; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_208; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_209; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_210; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_211; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_212; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_213; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_214; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_215; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_216; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_217; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_218; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_219; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_220; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_221; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_222; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_223; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_224; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_225; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_226; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_227; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_228; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_229; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_230; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_231; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_232; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_233; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_234; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_235; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_236; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_237; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_238; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_239; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_240; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_241; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_242; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_243; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_244; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_245; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_246; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_247; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_248; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_249; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_250; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_251; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_252; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_253; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_254; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_255; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_0; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_1; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_2; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_3; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_4; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_5; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_6; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_7; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_8; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_9; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_10; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_11; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_12; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_13; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_14; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_out_header_15; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 62:25]
  wire [15:0] proc_3_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 62:25]
  wire [1:0] proc_3_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 62:25]
  wire  proc_3_io_pipe_phv_out_next_config_id; // @[ipsa.scala 62:25]
  wire  proc_3_io_mod_par_mod_en; // @[ipsa.scala 62:25]
  wire  proc_3_io_mod_par_mod_last_mau_id_mod; // @[ipsa.scala 62:25]
  wire [1:0] proc_3_io_mod_par_mod_last_mau_id; // @[ipsa.scala 62:25]
  wire [1:0] proc_3_io_mod_par_mod_cs; // @[ipsa.scala 62:25]
  wire  proc_3_io_mod_par_mod_module_mod_state_id_mod; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mod_par_mod_module_mod_state_id; // @[ipsa.scala 62:25]
  wire  proc_3_io_mod_par_mod_module_mod_sram_w_cs; // @[ipsa.scala 62:25]
  wire  proc_3_io_mod_par_mod_module_mod_sram_w_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mod_par_mod_module_mod_sram_w_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mod_par_mod_module_mod_sram_w_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mod_mat_mod_en; // @[ipsa.scala 62:25]
  wire  proc_3_io_mod_mat_mod_config_id; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mod_mat_mod_key_mod_header_id; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mod_mat_mod_key_mod_internal_offset; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mod_mat_mod_key_mod_key_length; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_0; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_1; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_2; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_3; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_4; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_5; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_6; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_7; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_8; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_9; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_10; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_11; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_12; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_13; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_14; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_15; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_16; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_17; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_18; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_19; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_20; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_21; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_22; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_23; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_24; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_25; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_26; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_27; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_28; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_29; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_30; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_31; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_32; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_33; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_34; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_35; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_36; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_37; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_38; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_39; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_40; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_41; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_42; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_43; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_44; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_45; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_46; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_47; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_48; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_49; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_50; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_51; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_52; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_53; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_54; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_55; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_56; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_57; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_58; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_59; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_60; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_61; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_62; // @[ipsa.scala 62:25]
  wire [5:0] proc_3_io_mod_mat_mod_table_mod_sram_id_table_63; // @[ipsa.scala 62:25]
  wire [6:0] proc_3_io_mod_mat_mod_table_mod_table_width; // @[ipsa.scala 62:25]
  wire [6:0] proc_3_io_mod_mat_mod_table_mod_table_depth; // @[ipsa.scala 62:25]
  wire  proc_3_io_mod_act_mod_en_0; // @[ipsa.scala 62:25]
  wire  proc_3_io_mod_act_mod_en_1; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mod_act_mod_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mod_act_mod_data_0; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mod_act_mod_data_1; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_0_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_0_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_0_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_1_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_1_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_1_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_2_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_2_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_2_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_3_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_3_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_3_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_4_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_4_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_4_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_5_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_5_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_5_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_6_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_6_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_6_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_7_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_7_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_7_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_8_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_8_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_8_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_9_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_9_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_9_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_10_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_10_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_10_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_11_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_11_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_11_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_12_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_12_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_12_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_13_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_13_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_13_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_14_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_14_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_14_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_15_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_15_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_15_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_16_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_16_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_16_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_17_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_17_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_17_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_18_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_18_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_18_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_19_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_19_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_19_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_20_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_20_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_20_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_21_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_21_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_21_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_22_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_22_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_22_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_23_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_23_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_23_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_24_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_24_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_24_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_25_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_25_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_25_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_26_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_26_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_26_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_27_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_27_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_27_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_28_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_28_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_28_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_29_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_29_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_29_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_30_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_30_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_30_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_31_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_31_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_31_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_32_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_32_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_32_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_33_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_33_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_33_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_34_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_34_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_34_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_35_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_35_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_35_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_36_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_36_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_36_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_37_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_37_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_37_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_38_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_38_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_38_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_39_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_39_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_39_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_40_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_40_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_40_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_41_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_41_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_41_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_42_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_42_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_42_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_43_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_43_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_43_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_44_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_44_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_44_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_45_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_45_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_45_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_46_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_46_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_46_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_47_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_47_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_47_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_48_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_48_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_48_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_49_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_49_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_49_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_50_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_50_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_50_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_51_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_51_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_51_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_52_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_52_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_52_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_53_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_53_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_53_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_54_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_54_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_54_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_55_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_55_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_55_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_56_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_56_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_56_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_57_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_57_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_57_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_58_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_58_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_58_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_59_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_59_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_59_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_60_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_60_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_60_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_61_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_61_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_61_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_62_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_62_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_62_data; // @[ipsa.scala 62:25]
  wire  proc_3_io_mem_cluster_63_en; // @[ipsa.scala 62:25]
  wire [7:0] proc_3_io_mem_cluster_63_addr; // @[ipsa.scala 62:25]
  wire [63:0] proc_3_io_mem_cluster_63_data; // @[ipsa.scala 62:25]
  wire  sram_cluster_0_clock; // @[ipsa.scala 68:25]
  wire [5:0] sram_cluster_0_io_w_wcs; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_w_w_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_w_w_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_w_w_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_0_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_0_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_0_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_1_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_1_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_1_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_2_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_2_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_2_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_3_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_3_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_3_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_4_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_4_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_4_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_5_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_5_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_5_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_6_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_6_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_6_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_7_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_7_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_7_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_8_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_8_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_8_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_9_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_9_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_9_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_10_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_10_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_10_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_11_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_11_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_11_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_12_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_12_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_12_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_13_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_13_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_13_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_14_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_14_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_14_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_15_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_15_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_15_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_16_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_16_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_16_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_17_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_17_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_17_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_18_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_18_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_18_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_19_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_19_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_19_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_20_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_20_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_20_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_21_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_21_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_21_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_22_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_22_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_22_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_23_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_23_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_23_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_24_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_24_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_24_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_25_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_25_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_25_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_26_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_26_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_26_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_27_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_27_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_27_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_28_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_28_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_28_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_29_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_29_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_29_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_30_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_30_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_30_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_31_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_31_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_31_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_32_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_32_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_32_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_33_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_33_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_33_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_34_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_34_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_34_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_35_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_35_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_35_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_36_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_36_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_36_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_37_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_37_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_37_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_38_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_38_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_38_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_39_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_39_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_39_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_40_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_40_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_40_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_41_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_41_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_41_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_42_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_42_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_42_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_43_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_43_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_43_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_44_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_44_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_44_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_45_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_45_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_45_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_46_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_46_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_46_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_47_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_47_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_47_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_48_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_48_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_48_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_49_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_49_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_49_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_50_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_50_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_50_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_51_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_51_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_51_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_52_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_52_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_52_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_53_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_53_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_53_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_54_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_54_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_54_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_55_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_55_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_55_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_56_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_56_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_56_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_57_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_57_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_57_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_58_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_58_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_58_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_59_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_59_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_59_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_60_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_60_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_60_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_61_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_61_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_61_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_62_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_62_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_62_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_0_cluster_63_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_0_cluster_63_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_0_cluster_63_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_0_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_0_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_0_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_1_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_1_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_1_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_2_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_2_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_2_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_3_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_3_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_3_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_4_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_4_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_4_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_5_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_5_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_5_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_6_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_6_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_6_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_7_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_7_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_7_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_8_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_8_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_8_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_9_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_9_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_9_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_10_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_10_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_10_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_11_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_11_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_11_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_12_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_12_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_12_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_13_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_13_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_13_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_14_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_14_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_14_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_15_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_15_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_15_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_16_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_16_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_16_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_17_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_17_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_17_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_18_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_18_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_18_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_19_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_19_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_19_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_20_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_20_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_20_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_21_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_21_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_21_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_22_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_22_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_22_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_23_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_23_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_23_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_24_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_24_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_24_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_25_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_25_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_25_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_26_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_26_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_26_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_27_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_27_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_27_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_28_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_28_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_28_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_29_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_29_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_29_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_30_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_30_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_30_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_31_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_31_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_31_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_32_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_32_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_32_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_33_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_33_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_33_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_34_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_34_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_34_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_35_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_35_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_35_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_36_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_36_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_36_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_37_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_37_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_37_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_38_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_38_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_38_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_39_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_39_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_39_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_40_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_40_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_40_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_41_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_41_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_41_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_42_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_42_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_42_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_43_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_43_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_43_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_44_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_44_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_44_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_45_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_45_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_45_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_46_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_46_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_46_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_47_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_47_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_47_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_48_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_48_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_48_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_49_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_49_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_49_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_50_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_50_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_50_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_51_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_51_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_51_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_52_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_52_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_52_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_53_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_53_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_53_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_54_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_54_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_54_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_55_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_55_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_55_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_56_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_56_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_56_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_57_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_57_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_57_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_58_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_58_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_58_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_59_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_59_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_59_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_60_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_60_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_60_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_61_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_61_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_61_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_62_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_62_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_62_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_1_cluster_63_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_1_cluster_63_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_1_cluster_63_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_0_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_0_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_0_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_1_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_1_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_1_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_2_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_2_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_2_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_3_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_3_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_3_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_4_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_4_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_4_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_5_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_5_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_5_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_6_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_6_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_6_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_7_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_7_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_7_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_8_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_8_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_8_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_9_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_9_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_9_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_10_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_10_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_10_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_11_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_11_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_11_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_12_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_12_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_12_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_13_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_13_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_13_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_14_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_14_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_14_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_15_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_15_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_15_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_16_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_16_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_16_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_17_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_17_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_17_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_18_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_18_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_18_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_19_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_19_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_19_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_20_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_20_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_20_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_21_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_21_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_21_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_22_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_22_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_22_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_23_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_23_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_23_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_24_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_24_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_24_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_25_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_25_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_25_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_26_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_26_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_26_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_27_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_27_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_27_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_28_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_28_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_28_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_29_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_29_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_29_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_30_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_30_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_30_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_31_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_31_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_31_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_32_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_32_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_32_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_33_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_33_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_33_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_34_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_34_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_34_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_35_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_35_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_35_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_36_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_36_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_36_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_37_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_37_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_37_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_38_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_38_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_38_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_39_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_39_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_39_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_40_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_40_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_40_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_41_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_41_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_41_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_42_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_42_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_42_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_43_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_43_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_43_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_44_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_44_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_44_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_45_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_45_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_45_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_46_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_46_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_46_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_47_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_47_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_47_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_48_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_48_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_48_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_49_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_49_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_49_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_50_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_50_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_50_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_51_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_51_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_51_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_52_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_52_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_52_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_53_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_53_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_53_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_54_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_54_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_54_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_55_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_55_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_55_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_56_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_56_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_56_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_57_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_57_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_57_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_58_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_58_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_58_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_59_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_59_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_59_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_60_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_60_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_60_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_61_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_61_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_61_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_62_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_62_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_62_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_2_cluster_63_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_2_cluster_63_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_2_cluster_63_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_0_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_0_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_0_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_1_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_1_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_1_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_2_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_2_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_2_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_3_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_3_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_3_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_4_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_4_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_4_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_5_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_5_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_5_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_6_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_6_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_6_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_7_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_7_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_7_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_8_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_8_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_8_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_9_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_9_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_9_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_10_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_10_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_10_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_11_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_11_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_11_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_12_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_12_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_12_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_13_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_13_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_13_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_14_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_14_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_14_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_15_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_15_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_15_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_16_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_16_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_16_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_17_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_17_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_17_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_18_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_18_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_18_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_19_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_19_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_19_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_20_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_20_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_20_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_21_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_21_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_21_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_22_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_22_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_22_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_23_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_23_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_23_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_24_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_24_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_24_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_25_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_25_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_25_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_26_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_26_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_26_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_27_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_27_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_27_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_28_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_28_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_28_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_29_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_29_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_29_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_30_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_30_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_30_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_31_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_31_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_31_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_32_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_32_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_32_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_33_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_33_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_33_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_34_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_34_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_34_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_35_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_35_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_35_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_36_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_36_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_36_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_37_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_37_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_37_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_38_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_38_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_38_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_39_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_39_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_39_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_40_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_40_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_40_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_41_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_41_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_41_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_42_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_42_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_42_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_43_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_43_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_43_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_44_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_44_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_44_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_45_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_45_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_45_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_46_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_46_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_46_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_47_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_47_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_47_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_48_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_48_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_48_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_49_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_49_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_49_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_50_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_50_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_50_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_51_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_51_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_51_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_52_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_52_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_52_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_53_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_53_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_53_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_54_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_54_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_54_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_55_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_55_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_55_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_56_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_56_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_56_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_57_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_57_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_57_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_58_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_58_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_58_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_59_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_59_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_59_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_60_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_60_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_60_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_61_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_61_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_61_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_62_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_62_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_62_data; // @[ipsa.scala 68:25]
  wire  sram_cluster_0_io_r_3_cluster_63_en; // @[ipsa.scala 68:25]
  wire [7:0] sram_cluster_0_io_r_3_cluster_63_addr; // @[ipsa.scala 68:25]
  wire [63:0] sram_cluster_0_io_r_3_cluster_63_data; // @[ipsa.scala 68:25]
  wire  init_clock; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_0; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_1; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_2; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_3; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_4; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_5; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_6; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_7; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_8; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_9; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_10; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_11; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_12; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_13; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_14; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_15; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_16; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_17; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_18; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_19; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_20; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_21; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_22; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_23; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_24; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_25; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_26; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_27; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_28; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_29; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_30; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_31; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_32; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_33; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_34; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_35; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_36; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_37; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_38; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_39; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_40; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_41; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_42; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_43; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_44; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_45; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_46; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_47; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_48; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_49; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_50; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_51; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_52; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_53; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_54; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_55; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_56; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_57; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_58; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_59; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_60; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_61; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_62; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_63; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_64; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_65; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_66; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_67; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_68; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_69; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_70; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_71; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_72; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_73; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_74; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_75; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_76; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_77; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_78; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_79; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_80; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_81; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_82; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_83; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_84; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_85; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_86; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_87; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_88; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_89; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_90; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_91; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_92; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_93; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_94; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_95; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_96; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_97; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_98; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_99; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_100; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_101; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_102; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_103; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_104; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_105; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_106; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_107; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_108; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_109; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_110; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_111; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_112; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_113; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_114; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_115; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_116; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_117; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_118; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_119; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_120; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_121; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_122; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_123; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_124; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_125; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_126; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_127; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_128; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_129; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_130; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_131; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_132; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_133; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_134; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_135; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_136; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_137; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_138; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_139; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_140; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_141; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_142; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_143; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_144; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_145; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_146; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_147; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_148; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_149; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_150; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_151; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_152; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_153; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_154; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_155; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_156; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_157; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_158; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_159; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_160; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_161; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_162; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_163; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_164; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_165; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_166; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_167; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_168; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_169; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_170; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_171; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_172; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_173; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_174; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_175; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_176; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_177; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_178; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_179; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_180; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_181; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_182; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_183; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_184; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_185; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_186; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_187; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_188; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_189; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_190; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_in_data_191; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_0; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_1; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_2; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_3; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_4; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_5; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_6; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_7; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_8; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_9; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_10; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_11; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_12; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_13; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_14; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_15; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_16; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_17; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_18; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_19; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_20; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_21; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_22; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_23; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_24; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_25; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_26; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_27; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_28; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_29; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_30; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_31; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_32; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_33; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_34; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_35; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_36; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_37; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_38; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_39; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_40; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_41; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_42; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_43; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_44; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_45; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_46; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_47; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_48; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_49; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_50; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_51; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_52; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_53; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_54; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_55; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_56; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_57; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_58; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_59; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_60; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_61; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_62; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_63; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_64; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_65; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_66; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_67; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_68; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_69; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_70; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_71; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_72; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_73; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_74; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_75; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_76; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_77; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_78; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_79; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_80; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_81; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_82; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_83; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_84; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_85; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_86; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_87; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_88; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_89; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_90; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_91; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_92; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_93; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_94; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_95; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_96; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_97; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_98; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_99; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_100; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_101; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_102; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_103; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_104; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_105; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_106; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_107; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_108; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_109; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_110; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_111; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_112; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_113; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_114; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_115; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_116; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_117; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_118; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_119; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_120; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_121; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_122; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_123; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_124; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_125; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_126; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_127; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_128; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_129; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_130; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_131; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_132; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_133; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_134; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_135; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_136; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_137; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_138; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_139; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_140; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_141; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_142; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_143; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_144; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_145; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_146; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_147; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_148; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_149; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_150; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_151; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_152; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_153; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_154; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_155; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_156; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_157; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_158; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_159; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_160; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_161; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_162; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_163; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_164; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_165; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_166; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_167; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_168; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_169; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_170; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_171; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_172; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_173; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_174; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_175; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_176; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_177; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_178; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_179; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_180; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_181; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_182; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_183; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_184; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_185; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_186; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_187; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_188; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_189; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_190; // @[ipsa.scala 80:22]
  wire [7:0] init_io_pipe_phv_out_data_191; // @[ipsa.scala 80:22]
  wire [1:0] init_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 80:22]
  wire [1:0] init_io_first_proc_id; // @[ipsa.scala 80:22]
  wire  trans_0_clock; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_0; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_1; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_2; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_3; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_4; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_5; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_6; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_7; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_8; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_9; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_10; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_11; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_12; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_13; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_14; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_15; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_16; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_17; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_18; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_19; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_20; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_21; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_22; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_23; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_24; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_25; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_26; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_27; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_28; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_29; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_30; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_31; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_32; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_33; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_34; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_35; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_36; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_37; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_38; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_39; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_40; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_41; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_42; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_43; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_44; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_45; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_46; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_47; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_48; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_49; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_50; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_51; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_52; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_53; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_54; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_55; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_56; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_57; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_58; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_59; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_60; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_61; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_62; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_63; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_64; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_65; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_66; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_67; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_68; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_69; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_70; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_71; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_72; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_73; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_74; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_75; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_76; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_77; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_78; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_79; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_80; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_81; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_82; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_83; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_84; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_85; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_86; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_87; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_88; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_89; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_90; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_91; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_92; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_93; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_94; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_95; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_96; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_97; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_98; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_99; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_100; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_101; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_102; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_103; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_104; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_105; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_106; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_107; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_108; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_109; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_110; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_111; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_112; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_113; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_114; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_115; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_116; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_117; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_118; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_119; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_120; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_121; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_122; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_123; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_124; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_125; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_126; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_127; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_128; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_129; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_130; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_131; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_132; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_133; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_134; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_135; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_136; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_137; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_138; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_139; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_140; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_141; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_142; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_143; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_144; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_145; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_146; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_147; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_148; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_149; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_150; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_151; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_152; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_153; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_154; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_155; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_156; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_157; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_158; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_159; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_160; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_161; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_162; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_163; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_164; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_165; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_166; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_167; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_168; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_169; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_170; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_171; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_172; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_173; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_174; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_175; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_176; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_177; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_178; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_179; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_180; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_181; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_182; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_183; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_184; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_185; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_186; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_187; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_188; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_189; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_190; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_191; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_192; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_193; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_194; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_195; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_196; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_197; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_198; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_199; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_200; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_201; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_202; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_203; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_204; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_205; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_206; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_207; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_208; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_209; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_210; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_211; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_212; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_213; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_214; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_215; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_216; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_217; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_218; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_219; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_220; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_221; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_222; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_223; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_224; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_225; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_226; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_227; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_228; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_229; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_230; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_231; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_232; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_233; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_234; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_235; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_236; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_237; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_238; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_239; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_240; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_241; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_242; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_243; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_244; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_245; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_246; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_247; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_248; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_249; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_250; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_251; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_252; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_253; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_254; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_data_255; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_0; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_1; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_2; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_3; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_4; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_5; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_6; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_7; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_8; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_9; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_10; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_11; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_12; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_13; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_14; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_in_header_15; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 85:25]
  wire [1:0] trans_0_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 85:25]
  wire  trans_0_io_pipe_phv_in_next_config_id; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_0; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_1; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_2; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_3; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_4; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_5; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_6; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_7; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_8; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_9; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_10; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_11; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_12; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_13; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_14; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_15; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_16; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_17; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_18; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_19; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_20; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_21; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_22; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_23; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_24; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_25; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_26; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_27; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_28; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_29; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_30; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_31; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_32; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_33; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_34; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_35; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_36; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_37; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_38; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_39; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_40; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_41; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_42; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_43; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_44; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_45; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_46; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_47; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_48; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_49; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_50; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_51; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_52; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_53; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_54; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_55; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_56; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_57; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_58; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_59; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_60; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_61; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_62; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_63; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_64; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_65; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_66; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_67; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_68; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_69; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_70; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_71; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_72; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_73; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_74; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_75; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_76; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_77; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_78; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_79; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_80; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_81; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_82; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_83; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_84; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_85; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_86; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_87; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_88; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_89; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_90; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_91; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_92; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_93; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_94; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_95; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_96; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_97; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_98; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_99; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_100; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_101; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_102; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_103; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_104; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_105; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_106; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_107; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_108; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_109; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_110; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_111; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_112; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_113; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_114; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_115; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_116; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_117; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_118; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_119; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_120; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_121; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_122; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_123; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_124; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_125; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_126; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_127; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_128; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_129; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_130; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_131; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_132; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_133; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_134; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_135; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_136; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_137; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_138; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_139; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_140; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_141; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_142; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_143; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_144; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_145; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_146; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_147; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_148; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_149; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_150; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_151; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_152; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_153; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_154; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_155; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_156; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_157; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_158; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_159; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_160; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_161; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_162; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_163; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_164; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_165; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_166; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_167; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_168; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_169; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_170; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_171; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_172; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_173; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_174; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_175; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_176; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_177; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_178; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_179; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_180; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_181; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_182; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_183; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_184; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_185; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_186; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_187; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_188; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_189; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_190; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_191; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_192; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_193; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_194; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_195; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_196; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_197; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_198; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_199; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_200; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_201; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_202; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_203; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_204; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_205; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_206; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_207; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_208; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_209; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_210; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_211; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_212; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_213; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_214; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_215; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_216; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_217; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_218; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_219; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_220; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_221; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_222; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_223; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_224; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_225; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_226; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_227; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_228; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_229; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_230; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_231; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_232; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_233; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_234; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_235; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_236; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_237; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_238; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_239; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_240; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_241; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_242; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_243; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_244; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_245; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_246; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_247; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_248; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_249; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_250; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_251; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_252; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_253; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_254; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_data_255; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_0; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_1; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_2; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_3; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_4; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_5; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_6; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_7; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_8; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_9; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_10; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_11; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_12; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_13; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_14; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_out_header_15; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 85:25]
  wire [7:0] trans_0_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 85:25]
  wire [15:0] trans_0_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 85:25]
  wire [1:0] trans_0_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 85:25]
  wire  trans_0_io_pipe_phv_out_next_config_id; // @[ipsa.scala 85:25]
  wire  trans_0_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 85:25]
  wire  trans_0_io_next_proc_exist; // @[ipsa.scala 85:25]
  wire [1:0] trans_0_io_next_proc_id_in; // @[ipsa.scala 85:25]
  wire [1:0] trans_0_io_next_proc_id_out; // @[ipsa.scala 85:25]
  wire  trans_1_clock; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_0; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_1; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_2; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_3; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_4; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_5; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_6; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_7; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_8; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_9; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_10; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_11; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_12; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_13; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_14; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_15; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_16; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_17; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_18; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_19; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_20; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_21; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_22; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_23; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_24; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_25; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_26; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_27; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_28; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_29; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_30; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_31; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_32; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_33; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_34; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_35; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_36; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_37; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_38; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_39; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_40; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_41; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_42; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_43; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_44; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_45; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_46; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_47; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_48; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_49; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_50; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_51; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_52; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_53; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_54; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_55; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_56; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_57; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_58; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_59; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_60; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_61; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_62; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_63; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_64; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_65; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_66; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_67; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_68; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_69; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_70; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_71; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_72; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_73; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_74; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_75; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_76; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_77; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_78; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_79; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_80; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_81; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_82; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_83; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_84; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_85; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_86; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_87; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_88; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_89; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_90; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_91; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_92; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_93; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_94; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_95; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_96; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_97; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_98; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_99; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_100; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_101; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_102; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_103; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_104; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_105; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_106; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_107; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_108; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_109; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_110; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_111; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_112; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_113; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_114; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_115; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_116; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_117; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_118; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_119; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_120; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_121; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_122; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_123; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_124; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_125; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_126; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_127; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_128; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_129; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_130; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_131; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_132; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_133; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_134; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_135; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_136; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_137; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_138; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_139; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_140; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_141; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_142; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_143; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_144; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_145; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_146; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_147; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_148; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_149; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_150; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_151; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_152; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_153; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_154; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_155; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_156; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_157; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_158; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_159; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_160; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_161; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_162; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_163; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_164; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_165; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_166; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_167; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_168; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_169; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_170; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_171; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_172; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_173; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_174; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_175; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_176; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_177; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_178; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_179; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_180; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_181; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_182; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_183; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_184; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_185; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_186; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_187; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_188; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_189; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_190; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_191; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_192; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_193; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_194; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_195; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_196; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_197; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_198; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_199; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_200; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_201; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_202; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_203; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_204; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_205; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_206; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_207; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_208; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_209; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_210; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_211; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_212; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_213; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_214; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_215; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_216; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_217; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_218; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_219; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_220; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_221; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_222; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_223; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_224; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_225; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_226; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_227; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_228; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_229; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_230; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_231; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_232; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_233; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_234; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_235; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_236; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_237; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_238; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_239; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_240; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_241; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_242; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_243; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_244; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_245; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_246; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_247; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_248; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_249; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_250; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_251; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_252; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_253; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_254; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_data_255; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_0; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_1; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_2; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_3; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_4; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_5; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_6; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_7; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_8; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_9; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_10; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_11; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_12; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_13; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_14; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_in_header_15; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 85:25]
  wire [1:0] trans_1_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 85:25]
  wire  trans_1_io_pipe_phv_in_next_config_id; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_0; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_1; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_2; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_3; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_4; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_5; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_6; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_7; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_8; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_9; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_10; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_11; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_12; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_13; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_14; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_15; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_16; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_17; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_18; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_19; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_20; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_21; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_22; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_23; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_24; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_25; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_26; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_27; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_28; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_29; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_30; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_31; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_32; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_33; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_34; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_35; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_36; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_37; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_38; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_39; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_40; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_41; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_42; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_43; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_44; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_45; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_46; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_47; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_48; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_49; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_50; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_51; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_52; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_53; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_54; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_55; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_56; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_57; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_58; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_59; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_60; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_61; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_62; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_63; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_64; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_65; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_66; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_67; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_68; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_69; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_70; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_71; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_72; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_73; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_74; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_75; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_76; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_77; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_78; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_79; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_80; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_81; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_82; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_83; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_84; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_85; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_86; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_87; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_88; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_89; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_90; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_91; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_92; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_93; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_94; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_95; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_96; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_97; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_98; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_99; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_100; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_101; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_102; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_103; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_104; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_105; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_106; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_107; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_108; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_109; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_110; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_111; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_112; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_113; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_114; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_115; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_116; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_117; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_118; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_119; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_120; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_121; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_122; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_123; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_124; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_125; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_126; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_127; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_128; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_129; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_130; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_131; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_132; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_133; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_134; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_135; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_136; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_137; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_138; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_139; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_140; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_141; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_142; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_143; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_144; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_145; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_146; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_147; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_148; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_149; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_150; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_151; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_152; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_153; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_154; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_155; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_156; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_157; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_158; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_159; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_160; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_161; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_162; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_163; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_164; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_165; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_166; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_167; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_168; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_169; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_170; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_171; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_172; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_173; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_174; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_175; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_176; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_177; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_178; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_179; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_180; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_181; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_182; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_183; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_184; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_185; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_186; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_187; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_188; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_189; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_190; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_191; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_192; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_193; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_194; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_195; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_196; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_197; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_198; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_199; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_200; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_201; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_202; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_203; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_204; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_205; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_206; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_207; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_208; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_209; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_210; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_211; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_212; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_213; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_214; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_215; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_216; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_217; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_218; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_219; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_220; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_221; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_222; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_223; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_224; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_225; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_226; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_227; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_228; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_229; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_230; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_231; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_232; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_233; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_234; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_235; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_236; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_237; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_238; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_239; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_240; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_241; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_242; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_243; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_244; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_245; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_246; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_247; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_248; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_249; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_250; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_251; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_252; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_253; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_254; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_data_255; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_0; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_1; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_2; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_3; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_4; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_5; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_6; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_7; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_8; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_9; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_10; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_11; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_12; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_13; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_14; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_out_header_15; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 85:25]
  wire [7:0] trans_1_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 85:25]
  wire [15:0] trans_1_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 85:25]
  wire [1:0] trans_1_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 85:25]
  wire  trans_1_io_pipe_phv_out_next_config_id; // @[ipsa.scala 85:25]
  wire  trans_1_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 85:25]
  wire  trans_1_io_next_proc_exist; // @[ipsa.scala 85:25]
  wire [1:0] trans_1_io_next_proc_id_in; // @[ipsa.scala 85:25]
  wire [1:0] trans_1_io_next_proc_id_out; // @[ipsa.scala 85:25]
  wire  trans_2_clock; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_0; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_1; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_2; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_3; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_4; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_5; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_6; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_7; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_8; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_9; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_10; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_11; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_12; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_13; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_14; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_15; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_16; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_17; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_18; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_19; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_20; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_21; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_22; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_23; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_24; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_25; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_26; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_27; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_28; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_29; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_30; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_31; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_32; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_33; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_34; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_35; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_36; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_37; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_38; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_39; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_40; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_41; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_42; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_43; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_44; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_45; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_46; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_47; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_48; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_49; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_50; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_51; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_52; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_53; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_54; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_55; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_56; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_57; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_58; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_59; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_60; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_61; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_62; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_63; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_64; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_65; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_66; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_67; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_68; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_69; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_70; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_71; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_72; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_73; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_74; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_75; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_76; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_77; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_78; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_79; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_80; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_81; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_82; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_83; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_84; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_85; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_86; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_87; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_88; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_89; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_90; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_91; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_92; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_93; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_94; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_95; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_96; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_97; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_98; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_99; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_100; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_101; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_102; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_103; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_104; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_105; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_106; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_107; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_108; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_109; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_110; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_111; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_112; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_113; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_114; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_115; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_116; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_117; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_118; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_119; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_120; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_121; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_122; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_123; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_124; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_125; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_126; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_127; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_128; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_129; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_130; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_131; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_132; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_133; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_134; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_135; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_136; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_137; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_138; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_139; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_140; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_141; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_142; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_143; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_144; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_145; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_146; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_147; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_148; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_149; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_150; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_151; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_152; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_153; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_154; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_155; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_156; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_157; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_158; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_159; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_160; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_161; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_162; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_163; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_164; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_165; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_166; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_167; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_168; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_169; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_170; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_171; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_172; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_173; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_174; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_175; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_176; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_177; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_178; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_179; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_180; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_181; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_182; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_183; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_184; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_185; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_186; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_187; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_188; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_189; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_190; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_191; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_192; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_193; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_194; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_195; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_196; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_197; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_198; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_199; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_200; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_201; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_202; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_203; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_204; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_205; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_206; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_207; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_208; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_209; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_210; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_211; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_212; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_213; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_214; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_215; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_216; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_217; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_218; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_219; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_220; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_221; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_222; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_223; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_224; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_225; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_226; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_227; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_228; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_229; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_230; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_231; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_232; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_233; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_234; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_235; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_236; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_237; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_238; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_239; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_240; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_241; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_242; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_243; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_244; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_245; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_246; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_247; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_248; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_249; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_250; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_251; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_252; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_253; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_254; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_data_255; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_0; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_1; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_2; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_3; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_4; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_5; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_6; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_7; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_8; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_9; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_10; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_11; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_12; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_13; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_14; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_in_header_15; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 85:25]
  wire [1:0] trans_2_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 85:25]
  wire  trans_2_io_pipe_phv_in_next_config_id; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_0; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_1; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_2; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_3; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_4; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_5; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_6; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_7; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_8; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_9; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_10; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_11; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_12; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_13; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_14; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_15; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_16; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_17; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_18; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_19; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_20; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_21; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_22; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_23; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_24; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_25; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_26; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_27; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_28; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_29; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_30; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_31; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_32; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_33; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_34; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_35; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_36; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_37; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_38; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_39; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_40; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_41; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_42; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_43; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_44; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_45; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_46; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_47; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_48; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_49; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_50; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_51; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_52; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_53; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_54; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_55; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_56; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_57; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_58; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_59; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_60; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_61; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_62; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_63; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_64; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_65; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_66; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_67; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_68; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_69; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_70; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_71; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_72; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_73; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_74; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_75; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_76; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_77; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_78; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_79; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_80; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_81; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_82; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_83; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_84; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_85; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_86; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_87; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_88; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_89; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_90; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_91; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_92; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_93; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_94; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_95; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_96; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_97; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_98; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_99; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_100; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_101; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_102; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_103; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_104; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_105; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_106; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_107; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_108; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_109; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_110; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_111; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_112; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_113; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_114; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_115; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_116; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_117; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_118; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_119; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_120; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_121; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_122; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_123; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_124; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_125; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_126; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_127; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_128; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_129; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_130; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_131; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_132; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_133; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_134; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_135; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_136; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_137; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_138; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_139; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_140; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_141; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_142; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_143; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_144; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_145; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_146; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_147; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_148; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_149; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_150; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_151; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_152; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_153; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_154; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_155; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_156; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_157; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_158; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_159; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_160; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_161; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_162; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_163; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_164; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_165; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_166; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_167; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_168; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_169; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_170; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_171; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_172; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_173; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_174; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_175; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_176; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_177; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_178; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_179; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_180; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_181; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_182; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_183; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_184; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_185; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_186; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_187; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_188; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_189; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_190; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_191; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_192; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_193; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_194; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_195; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_196; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_197; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_198; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_199; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_200; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_201; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_202; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_203; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_204; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_205; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_206; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_207; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_208; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_209; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_210; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_211; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_212; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_213; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_214; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_215; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_216; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_217; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_218; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_219; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_220; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_221; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_222; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_223; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_224; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_225; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_226; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_227; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_228; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_229; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_230; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_231; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_232; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_233; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_234; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_235; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_236; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_237; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_238; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_239; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_240; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_241; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_242; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_243; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_244; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_245; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_246; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_247; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_248; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_249; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_250; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_251; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_252; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_253; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_254; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_data_255; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_0; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_1; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_2; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_3; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_4; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_5; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_6; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_7; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_8; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_9; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_10; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_11; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_12; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_13; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_14; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_out_header_15; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 85:25]
  wire [7:0] trans_2_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 85:25]
  wire [15:0] trans_2_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 85:25]
  wire [1:0] trans_2_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 85:25]
  wire  trans_2_io_pipe_phv_out_next_config_id; // @[ipsa.scala 85:25]
  wire  trans_2_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 85:25]
  wire  trans_2_io_next_proc_exist; // @[ipsa.scala 85:25]
  wire [1:0] trans_2_io_next_proc_id_in; // @[ipsa.scala 85:25]
  wire [1:0] trans_2_io_next_proc_id_out; // @[ipsa.scala 85:25]
  wire  trans_3_clock; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_0; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_1; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_2; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_3; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_4; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_5; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_6; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_7; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_8; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_9; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_10; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_11; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_12; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_13; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_14; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_15; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_16; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_17; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_18; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_19; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_20; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_21; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_22; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_23; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_24; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_25; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_26; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_27; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_28; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_29; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_30; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_31; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_32; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_33; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_34; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_35; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_36; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_37; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_38; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_39; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_40; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_41; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_42; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_43; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_44; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_45; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_46; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_47; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_48; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_49; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_50; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_51; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_52; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_53; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_54; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_55; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_56; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_57; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_58; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_59; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_60; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_61; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_62; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_63; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_64; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_65; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_66; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_67; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_68; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_69; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_70; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_71; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_72; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_73; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_74; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_75; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_76; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_77; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_78; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_79; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_80; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_81; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_82; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_83; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_84; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_85; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_86; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_87; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_88; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_89; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_90; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_91; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_92; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_93; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_94; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_95; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_96; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_97; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_98; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_99; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_100; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_101; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_102; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_103; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_104; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_105; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_106; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_107; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_108; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_109; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_110; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_111; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_112; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_113; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_114; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_115; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_116; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_117; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_118; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_119; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_120; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_121; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_122; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_123; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_124; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_125; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_126; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_127; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_128; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_129; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_130; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_131; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_132; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_133; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_134; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_135; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_136; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_137; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_138; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_139; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_140; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_141; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_142; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_143; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_144; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_145; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_146; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_147; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_148; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_149; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_150; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_151; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_152; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_153; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_154; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_155; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_156; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_157; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_158; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_159; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_160; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_161; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_162; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_163; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_164; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_165; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_166; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_167; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_168; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_169; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_170; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_171; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_172; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_173; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_174; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_175; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_176; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_177; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_178; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_179; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_180; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_181; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_182; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_183; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_184; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_185; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_186; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_187; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_188; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_189; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_190; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_191; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_192; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_193; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_194; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_195; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_196; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_197; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_198; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_199; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_200; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_201; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_202; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_203; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_204; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_205; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_206; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_207; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_208; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_209; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_210; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_211; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_212; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_213; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_214; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_215; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_216; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_217; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_218; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_219; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_220; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_221; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_222; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_223; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_224; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_225; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_226; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_227; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_228; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_229; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_230; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_231; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_232; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_233; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_234; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_235; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_236; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_237; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_238; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_239; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_240; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_241; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_242; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_243; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_244; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_245; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_246; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_247; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_248; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_249; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_250; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_251; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_252; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_253; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_254; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_data_255; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_0; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_1; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_2; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_3; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_4; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_5; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_6; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_7; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_8; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_9; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_10; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_11; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_12; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_13; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_14; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_in_header_15; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_parse_current_state; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_in_parse_current_offset; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_in_parse_transition_field; // @[ipsa.scala 85:25]
  wire [1:0] trans_3_io_pipe_phv_in_next_processor_id; // @[ipsa.scala 85:25]
  wire  trans_3_io_pipe_phv_in_next_config_id; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_0; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_1; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_2; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_3; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_4; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_5; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_6; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_7; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_8; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_9; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_10; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_11; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_12; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_13; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_14; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_15; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_16; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_17; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_18; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_19; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_20; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_21; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_22; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_23; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_24; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_25; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_26; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_27; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_28; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_29; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_30; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_31; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_32; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_33; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_34; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_35; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_36; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_37; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_38; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_39; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_40; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_41; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_42; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_43; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_44; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_45; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_46; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_47; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_48; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_49; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_50; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_51; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_52; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_53; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_54; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_55; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_56; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_57; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_58; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_59; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_60; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_61; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_62; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_63; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_64; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_65; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_66; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_67; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_68; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_69; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_70; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_71; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_72; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_73; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_74; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_75; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_76; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_77; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_78; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_79; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_80; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_81; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_82; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_83; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_84; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_85; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_86; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_87; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_88; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_89; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_90; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_91; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_92; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_93; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_94; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_95; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_96; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_97; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_98; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_99; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_100; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_101; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_102; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_103; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_104; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_105; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_106; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_107; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_108; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_109; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_110; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_111; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_112; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_113; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_114; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_115; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_116; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_117; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_118; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_119; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_120; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_121; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_122; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_123; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_124; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_125; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_126; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_127; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_128; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_129; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_130; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_131; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_132; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_133; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_134; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_135; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_136; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_137; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_138; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_139; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_140; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_141; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_142; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_143; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_144; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_145; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_146; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_147; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_148; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_149; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_150; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_151; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_152; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_153; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_154; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_155; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_156; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_157; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_158; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_159; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_160; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_161; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_162; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_163; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_164; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_165; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_166; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_167; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_168; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_169; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_170; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_171; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_172; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_173; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_174; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_175; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_176; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_177; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_178; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_179; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_180; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_181; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_182; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_183; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_184; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_185; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_186; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_187; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_188; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_189; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_190; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_191; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_192; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_193; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_194; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_195; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_196; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_197; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_198; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_199; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_200; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_201; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_202; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_203; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_204; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_205; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_206; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_207; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_208; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_209; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_210; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_211; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_212; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_213; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_214; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_215; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_216; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_217; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_218; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_219; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_220; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_221; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_222; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_223; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_224; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_225; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_226; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_227; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_228; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_229; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_230; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_231; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_232; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_233; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_234; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_235; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_236; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_237; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_238; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_239; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_240; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_241; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_242; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_243; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_244; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_245; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_246; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_247; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_248; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_249; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_250; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_251; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_252; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_253; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_254; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_data_255; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_0; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_1; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_2; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_3; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_4; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_5; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_6; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_7; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_8; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_9; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_10; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_11; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_12; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_13; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_14; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_out_header_15; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 85:25]
  wire [7:0] trans_3_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 85:25]
  wire [15:0] trans_3_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 85:25]
  wire [1:0] trans_3_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 85:25]
  wire  trans_3_io_pipe_phv_out_next_config_id; // @[ipsa.scala 85:25]
  wire  trans_3_io_pipe_phv_out_is_valid_processor; // @[ipsa.scala 85:25]
  wire  trans_3_io_next_proc_exist; // @[ipsa.scala 85:25]
  wire [1:0] trans_3_io_next_proc_id_in; // @[ipsa.scala 85:25]
  wire [1:0] trans_3_io_next_proc_id_out; // @[ipsa.scala 85:25]
  reg [1:0] first_proc_id; // @[ipsa.scala 48:28]
  reg [1:0] last_proc_id; // @[ipsa.scala 49:28]
  reg [1:0] next_proc_id_0; // @[ipsa.scala 50:28]
  reg [1:0] next_proc_id_1; // @[ipsa.scala 50:28]
  reg [1:0] next_proc_id_2; // @[ipsa.scala 50:28]
  reg [1:0] next_proc_id_3; // @[ipsa.scala 50:28]
  reg [7:0] recv_0_data_0; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_1; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_2; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_3; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_4; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_5; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_6; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_7; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_8; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_9; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_10; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_11; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_12; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_13; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_14; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_15; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_16; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_17; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_18; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_19; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_20; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_21; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_22; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_23; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_24; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_25; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_26; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_27; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_28; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_29; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_30; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_31; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_32; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_33; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_34; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_35; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_36; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_37; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_38; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_39; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_40; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_41; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_42; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_43; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_44; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_45; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_46; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_47; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_48; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_49; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_50; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_51; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_52; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_53; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_54; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_55; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_56; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_57; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_58; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_59; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_60; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_61; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_62; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_63; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_64; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_65; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_66; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_67; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_68; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_69; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_70; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_71; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_72; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_73; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_74; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_75; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_76; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_77; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_78; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_79; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_80; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_81; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_82; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_83; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_84; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_85; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_86; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_87; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_88; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_89; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_90; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_91; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_92; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_93; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_94; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_95; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_96; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_97; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_98; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_99; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_100; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_101; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_102; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_103; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_104; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_105; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_106; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_107; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_108; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_109; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_110; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_111; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_112; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_113; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_114; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_115; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_116; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_117; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_118; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_119; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_120; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_121; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_122; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_123; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_124; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_125; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_126; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_127; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_128; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_129; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_130; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_131; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_132; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_133; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_134; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_135; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_136; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_137; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_138; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_139; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_140; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_141; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_142; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_143; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_144; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_145; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_146; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_147; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_148; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_149; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_150; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_151; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_152; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_153; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_154; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_155; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_156; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_157; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_158; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_159; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_160; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_161; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_162; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_163; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_164; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_165; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_166; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_167; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_168; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_169; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_170; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_171; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_172; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_173; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_174; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_175; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_176; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_177; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_178; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_179; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_180; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_181; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_182; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_183; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_184; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_185; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_186; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_187; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_188; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_189; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_190; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_191; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_192; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_193; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_194; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_195; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_196; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_197; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_198; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_199; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_200; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_201; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_202; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_203; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_204; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_205; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_206; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_207; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_208; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_209; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_210; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_211; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_212; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_213; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_214; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_215; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_216; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_217; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_218; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_219; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_220; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_221; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_222; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_223; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_224; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_225; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_226; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_227; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_228; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_229; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_230; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_231; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_232; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_233; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_234; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_235; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_236; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_237; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_238; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_239; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_240; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_241; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_242; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_243; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_244; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_245; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_246; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_247; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_248; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_249; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_250; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_251; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_252; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_253; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_254; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_data_255; // @[ipsa.scala 60:19]
  reg [15:0] recv_0_header_0; // @[ipsa.scala 60:19]
  reg [15:0] recv_0_header_1; // @[ipsa.scala 60:19]
  reg [15:0] recv_0_header_2; // @[ipsa.scala 60:19]
  reg [15:0] recv_0_header_3; // @[ipsa.scala 60:19]
  reg [15:0] recv_0_header_4; // @[ipsa.scala 60:19]
  reg [15:0] recv_0_header_5; // @[ipsa.scala 60:19]
  reg [15:0] recv_0_header_6; // @[ipsa.scala 60:19]
  reg [15:0] recv_0_header_7; // @[ipsa.scala 60:19]
  reg [15:0] recv_0_header_8; // @[ipsa.scala 60:19]
  reg [15:0] recv_0_header_9; // @[ipsa.scala 60:19]
  reg [15:0] recv_0_header_10; // @[ipsa.scala 60:19]
  reg [15:0] recv_0_header_11; // @[ipsa.scala 60:19]
  reg [15:0] recv_0_header_12; // @[ipsa.scala 60:19]
  reg [15:0] recv_0_header_13; // @[ipsa.scala 60:19]
  reg [15:0] recv_0_header_14; // @[ipsa.scala 60:19]
  reg [15:0] recv_0_header_15; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_parse_current_state; // @[ipsa.scala 60:19]
  reg [7:0] recv_0_parse_current_offset; // @[ipsa.scala 60:19]
  reg [15:0] recv_0_parse_transition_field; // @[ipsa.scala 60:19]
  reg [1:0] recv_0_next_processor_id; // @[ipsa.scala 60:19]
  reg  recv_0_next_config_id; // @[ipsa.scala 60:19]
  reg  recv_0_is_valid_processor; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_0; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_1; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_2; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_3; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_4; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_5; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_6; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_7; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_8; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_9; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_10; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_11; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_12; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_13; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_14; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_15; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_16; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_17; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_18; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_19; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_20; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_21; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_22; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_23; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_24; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_25; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_26; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_27; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_28; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_29; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_30; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_31; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_32; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_33; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_34; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_35; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_36; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_37; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_38; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_39; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_40; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_41; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_42; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_43; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_44; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_45; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_46; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_47; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_48; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_49; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_50; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_51; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_52; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_53; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_54; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_55; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_56; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_57; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_58; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_59; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_60; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_61; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_62; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_63; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_64; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_65; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_66; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_67; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_68; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_69; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_70; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_71; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_72; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_73; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_74; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_75; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_76; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_77; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_78; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_79; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_80; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_81; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_82; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_83; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_84; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_85; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_86; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_87; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_88; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_89; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_90; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_91; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_92; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_93; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_94; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_95; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_96; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_97; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_98; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_99; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_100; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_101; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_102; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_103; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_104; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_105; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_106; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_107; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_108; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_109; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_110; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_111; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_112; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_113; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_114; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_115; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_116; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_117; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_118; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_119; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_120; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_121; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_122; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_123; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_124; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_125; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_126; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_127; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_128; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_129; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_130; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_131; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_132; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_133; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_134; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_135; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_136; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_137; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_138; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_139; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_140; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_141; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_142; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_143; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_144; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_145; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_146; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_147; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_148; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_149; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_150; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_151; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_152; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_153; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_154; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_155; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_156; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_157; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_158; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_159; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_160; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_161; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_162; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_163; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_164; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_165; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_166; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_167; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_168; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_169; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_170; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_171; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_172; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_173; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_174; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_175; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_176; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_177; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_178; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_179; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_180; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_181; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_182; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_183; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_184; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_185; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_186; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_187; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_188; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_189; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_190; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_191; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_192; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_193; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_194; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_195; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_196; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_197; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_198; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_199; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_200; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_201; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_202; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_203; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_204; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_205; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_206; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_207; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_208; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_209; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_210; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_211; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_212; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_213; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_214; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_215; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_216; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_217; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_218; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_219; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_220; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_221; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_222; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_223; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_224; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_225; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_226; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_227; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_228; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_229; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_230; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_231; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_232; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_233; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_234; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_235; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_236; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_237; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_238; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_239; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_240; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_241; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_242; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_243; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_244; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_245; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_246; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_247; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_248; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_249; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_250; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_251; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_252; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_253; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_254; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_data_255; // @[ipsa.scala 60:19]
  reg [15:0] recv_1_header_0; // @[ipsa.scala 60:19]
  reg [15:0] recv_1_header_1; // @[ipsa.scala 60:19]
  reg [15:0] recv_1_header_2; // @[ipsa.scala 60:19]
  reg [15:0] recv_1_header_3; // @[ipsa.scala 60:19]
  reg [15:0] recv_1_header_4; // @[ipsa.scala 60:19]
  reg [15:0] recv_1_header_5; // @[ipsa.scala 60:19]
  reg [15:0] recv_1_header_6; // @[ipsa.scala 60:19]
  reg [15:0] recv_1_header_7; // @[ipsa.scala 60:19]
  reg [15:0] recv_1_header_8; // @[ipsa.scala 60:19]
  reg [15:0] recv_1_header_9; // @[ipsa.scala 60:19]
  reg [15:0] recv_1_header_10; // @[ipsa.scala 60:19]
  reg [15:0] recv_1_header_11; // @[ipsa.scala 60:19]
  reg [15:0] recv_1_header_12; // @[ipsa.scala 60:19]
  reg [15:0] recv_1_header_13; // @[ipsa.scala 60:19]
  reg [15:0] recv_1_header_14; // @[ipsa.scala 60:19]
  reg [15:0] recv_1_header_15; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_parse_current_state; // @[ipsa.scala 60:19]
  reg [7:0] recv_1_parse_current_offset; // @[ipsa.scala 60:19]
  reg [15:0] recv_1_parse_transition_field; // @[ipsa.scala 60:19]
  reg [1:0] recv_1_next_processor_id; // @[ipsa.scala 60:19]
  reg  recv_1_next_config_id; // @[ipsa.scala 60:19]
  reg  recv_1_is_valid_processor; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_0; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_1; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_2; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_3; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_4; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_5; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_6; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_7; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_8; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_9; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_10; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_11; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_12; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_13; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_14; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_15; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_16; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_17; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_18; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_19; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_20; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_21; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_22; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_23; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_24; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_25; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_26; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_27; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_28; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_29; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_30; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_31; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_32; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_33; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_34; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_35; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_36; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_37; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_38; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_39; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_40; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_41; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_42; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_43; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_44; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_45; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_46; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_47; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_48; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_49; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_50; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_51; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_52; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_53; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_54; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_55; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_56; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_57; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_58; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_59; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_60; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_61; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_62; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_63; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_64; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_65; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_66; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_67; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_68; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_69; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_70; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_71; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_72; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_73; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_74; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_75; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_76; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_77; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_78; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_79; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_80; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_81; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_82; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_83; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_84; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_85; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_86; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_87; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_88; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_89; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_90; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_91; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_92; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_93; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_94; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_95; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_96; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_97; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_98; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_99; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_100; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_101; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_102; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_103; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_104; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_105; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_106; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_107; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_108; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_109; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_110; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_111; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_112; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_113; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_114; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_115; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_116; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_117; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_118; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_119; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_120; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_121; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_122; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_123; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_124; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_125; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_126; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_127; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_128; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_129; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_130; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_131; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_132; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_133; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_134; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_135; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_136; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_137; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_138; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_139; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_140; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_141; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_142; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_143; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_144; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_145; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_146; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_147; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_148; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_149; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_150; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_151; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_152; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_153; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_154; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_155; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_156; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_157; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_158; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_159; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_160; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_161; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_162; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_163; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_164; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_165; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_166; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_167; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_168; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_169; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_170; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_171; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_172; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_173; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_174; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_175; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_176; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_177; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_178; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_179; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_180; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_181; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_182; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_183; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_184; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_185; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_186; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_187; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_188; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_189; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_190; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_191; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_192; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_193; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_194; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_195; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_196; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_197; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_198; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_199; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_200; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_201; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_202; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_203; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_204; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_205; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_206; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_207; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_208; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_209; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_210; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_211; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_212; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_213; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_214; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_215; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_216; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_217; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_218; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_219; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_220; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_221; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_222; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_223; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_224; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_225; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_226; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_227; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_228; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_229; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_230; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_231; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_232; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_233; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_234; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_235; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_236; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_237; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_238; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_239; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_240; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_241; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_242; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_243; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_244; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_245; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_246; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_247; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_248; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_249; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_250; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_251; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_252; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_253; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_254; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_data_255; // @[ipsa.scala 60:19]
  reg [15:0] recv_2_header_0; // @[ipsa.scala 60:19]
  reg [15:0] recv_2_header_1; // @[ipsa.scala 60:19]
  reg [15:0] recv_2_header_2; // @[ipsa.scala 60:19]
  reg [15:0] recv_2_header_3; // @[ipsa.scala 60:19]
  reg [15:0] recv_2_header_4; // @[ipsa.scala 60:19]
  reg [15:0] recv_2_header_5; // @[ipsa.scala 60:19]
  reg [15:0] recv_2_header_6; // @[ipsa.scala 60:19]
  reg [15:0] recv_2_header_7; // @[ipsa.scala 60:19]
  reg [15:0] recv_2_header_8; // @[ipsa.scala 60:19]
  reg [15:0] recv_2_header_9; // @[ipsa.scala 60:19]
  reg [15:0] recv_2_header_10; // @[ipsa.scala 60:19]
  reg [15:0] recv_2_header_11; // @[ipsa.scala 60:19]
  reg [15:0] recv_2_header_12; // @[ipsa.scala 60:19]
  reg [15:0] recv_2_header_13; // @[ipsa.scala 60:19]
  reg [15:0] recv_2_header_14; // @[ipsa.scala 60:19]
  reg [15:0] recv_2_header_15; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_parse_current_state; // @[ipsa.scala 60:19]
  reg [7:0] recv_2_parse_current_offset; // @[ipsa.scala 60:19]
  reg [15:0] recv_2_parse_transition_field; // @[ipsa.scala 60:19]
  reg [1:0] recv_2_next_processor_id; // @[ipsa.scala 60:19]
  reg  recv_2_next_config_id; // @[ipsa.scala 60:19]
  reg  recv_2_is_valid_processor; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_0; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_1; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_2; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_3; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_4; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_5; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_6; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_7; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_8; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_9; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_10; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_11; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_12; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_13; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_14; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_15; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_16; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_17; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_18; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_19; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_20; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_21; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_22; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_23; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_24; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_25; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_26; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_27; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_28; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_29; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_30; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_31; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_32; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_33; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_34; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_35; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_36; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_37; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_38; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_39; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_40; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_41; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_42; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_43; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_44; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_45; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_46; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_47; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_48; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_49; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_50; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_51; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_52; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_53; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_54; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_55; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_56; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_57; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_58; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_59; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_60; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_61; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_62; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_63; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_64; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_65; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_66; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_67; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_68; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_69; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_70; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_71; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_72; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_73; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_74; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_75; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_76; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_77; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_78; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_79; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_80; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_81; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_82; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_83; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_84; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_85; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_86; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_87; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_88; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_89; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_90; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_91; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_92; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_93; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_94; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_95; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_96; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_97; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_98; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_99; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_100; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_101; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_102; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_103; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_104; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_105; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_106; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_107; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_108; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_109; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_110; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_111; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_112; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_113; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_114; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_115; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_116; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_117; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_118; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_119; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_120; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_121; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_122; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_123; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_124; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_125; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_126; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_127; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_128; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_129; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_130; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_131; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_132; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_133; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_134; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_135; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_136; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_137; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_138; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_139; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_140; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_141; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_142; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_143; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_144; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_145; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_146; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_147; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_148; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_149; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_150; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_151; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_152; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_153; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_154; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_155; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_156; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_157; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_158; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_159; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_160; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_161; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_162; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_163; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_164; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_165; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_166; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_167; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_168; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_169; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_170; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_171; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_172; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_173; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_174; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_175; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_176; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_177; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_178; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_179; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_180; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_181; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_182; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_183; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_184; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_185; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_186; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_187; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_188; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_189; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_190; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_191; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_192; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_193; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_194; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_195; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_196; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_197; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_198; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_199; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_200; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_201; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_202; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_203; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_204; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_205; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_206; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_207; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_208; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_209; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_210; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_211; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_212; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_213; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_214; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_215; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_216; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_217; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_218; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_219; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_220; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_221; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_222; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_223; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_224; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_225; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_226; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_227; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_228; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_229; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_230; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_231; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_232; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_233; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_234; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_235; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_236; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_237; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_238; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_239; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_240; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_241; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_242; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_243; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_244; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_245; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_246; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_247; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_248; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_249; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_250; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_251; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_252; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_253; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_254; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_data_255; // @[ipsa.scala 60:19]
  reg [15:0] recv_3_header_0; // @[ipsa.scala 60:19]
  reg [15:0] recv_3_header_1; // @[ipsa.scala 60:19]
  reg [15:0] recv_3_header_2; // @[ipsa.scala 60:19]
  reg [15:0] recv_3_header_3; // @[ipsa.scala 60:19]
  reg [15:0] recv_3_header_4; // @[ipsa.scala 60:19]
  reg [15:0] recv_3_header_5; // @[ipsa.scala 60:19]
  reg [15:0] recv_3_header_6; // @[ipsa.scala 60:19]
  reg [15:0] recv_3_header_7; // @[ipsa.scala 60:19]
  reg [15:0] recv_3_header_8; // @[ipsa.scala 60:19]
  reg [15:0] recv_3_header_9; // @[ipsa.scala 60:19]
  reg [15:0] recv_3_header_10; // @[ipsa.scala 60:19]
  reg [15:0] recv_3_header_11; // @[ipsa.scala 60:19]
  reg [15:0] recv_3_header_12; // @[ipsa.scala 60:19]
  reg [15:0] recv_3_header_13; // @[ipsa.scala 60:19]
  reg [15:0] recv_3_header_14; // @[ipsa.scala 60:19]
  reg [15:0] recv_3_header_15; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_parse_current_state; // @[ipsa.scala 60:19]
  reg [7:0] recv_3_parse_current_offset; // @[ipsa.scala 60:19]
  reg [15:0] recv_3_parse_transition_field; // @[ipsa.scala 60:19]
  reg [1:0] recv_3_next_processor_id; // @[ipsa.scala 60:19]
  reg  recv_3_next_config_id; // @[ipsa.scala 60:19]
  reg  recv_3_is_valid_processor; // @[ipsa.scala 60:19]
  wire [7:0] _GEN_28 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_0 : io_pipe_phv_in_data_0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_29 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_1 : io_pipe_phv_in_data_1; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_30 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_2 : io_pipe_phv_in_data_2; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_31 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_3 : io_pipe_phv_in_data_3; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_32 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_4 : io_pipe_phv_in_data_4; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_33 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_5 : io_pipe_phv_in_data_5; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_34 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_6 : io_pipe_phv_in_data_6; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_35 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_7 : io_pipe_phv_in_data_7; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_36 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_8 : io_pipe_phv_in_data_8; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_37 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_9 : io_pipe_phv_in_data_9; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_38 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_10 : io_pipe_phv_in_data_10; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_39 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_11 : io_pipe_phv_in_data_11; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_40 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_12 : io_pipe_phv_in_data_12; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_41 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_13 : io_pipe_phv_in_data_13; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_42 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_14 : io_pipe_phv_in_data_14; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_43 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_15 : io_pipe_phv_in_data_15; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_44 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_16 : io_pipe_phv_in_data_16; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_45 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_17 : io_pipe_phv_in_data_17; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_46 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_18 : io_pipe_phv_in_data_18; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_47 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_19 : io_pipe_phv_in_data_19; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_48 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_20 : io_pipe_phv_in_data_20; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_49 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_21 : io_pipe_phv_in_data_21; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_50 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_22 : io_pipe_phv_in_data_22; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_51 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_23 : io_pipe_phv_in_data_23; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_52 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_24 : io_pipe_phv_in_data_24; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_53 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_25 : io_pipe_phv_in_data_25; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_54 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_26 : io_pipe_phv_in_data_26; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_55 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_27 : io_pipe_phv_in_data_27; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_56 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_28 : io_pipe_phv_in_data_28; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_57 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_29 : io_pipe_phv_in_data_29; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_58 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_30 : io_pipe_phv_in_data_30; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_59 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_31 : io_pipe_phv_in_data_31; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_60 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_32 : io_pipe_phv_in_data_32; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_61 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_33 : io_pipe_phv_in_data_33; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_62 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_34 : io_pipe_phv_in_data_34; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_63 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_35 : io_pipe_phv_in_data_35; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_64 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_36 : io_pipe_phv_in_data_36; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_65 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_37 : io_pipe_phv_in_data_37; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_66 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_38 : io_pipe_phv_in_data_38; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_67 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_39 : io_pipe_phv_in_data_39; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_68 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_40 : io_pipe_phv_in_data_40; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_69 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_41 : io_pipe_phv_in_data_41; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_70 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_42 : io_pipe_phv_in_data_42; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_71 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_43 : io_pipe_phv_in_data_43; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_72 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_44 : io_pipe_phv_in_data_44; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_73 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_45 : io_pipe_phv_in_data_45; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_74 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_46 : io_pipe_phv_in_data_46; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_75 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_47 : io_pipe_phv_in_data_47; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_76 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_48 : io_pipe_phv_in_data_48; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_77 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_49 : io_pipe_phv_in_data_49; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_78 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_50 : io_pipe_phv_in_data_50; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_79 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_51 : io_pipe_phv_in_data_51; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_80 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_52 : io_pipe_phv_in_data_52; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_81 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_53 : io_pipe_phv_in_data_53; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_82 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_54 : io_pipe_phv_in_data_54; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_83 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_55 : io_pipe_phv_in_data_55; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_84 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_56 : io_pipe_phv_in_data_56; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_85 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_57 : io_pipe_phv_in_data_57; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_86 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_58 : io_pipe_phv_in_data_58; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_87 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_59 : io_pipe_phv_in_data_59; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_88 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_60 : io_pipe_phv_in_data_60; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_89 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_61 : io_pipe_phv_in_data_61; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_90 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_62 : io_pipe_phv_in_data_62; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_91 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_63 : io_pipe_phv_in_data_63; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_92 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_64 : io_pipe_phv_in_data_64; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_93 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_65 : io_pipe_phv_in_data_65; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_94 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_66 : io_pipe_phv_in_data_66; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_95 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_67 : io_pipe_phv_in_data_67; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_96 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_68 : io_pipe_phv_in_data_68; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_97 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_69 : io_pipe_phv_in_data_69; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_98 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_70 : io_pipe_phv_in_data_70; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_99 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_71 : io_pipe_phv_in_data_71; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_100 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_72 : io_pipe_phv_in_data_72; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_101 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_73 : io_pipe_phv_in_data_73; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_102 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_74 : io_pipe_phv_in_data_74; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_103 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_75 : io_pipe_phv_in_data_75; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_104 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_76 : io_pipe_phv_in_data_76; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_105 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_77 : io_pipe_phv_in_data_77; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_106 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_78 : io_pipe_phv_in_data_78; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_107 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_79 : io_pipe_phv_in_data_79; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_108 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_80 : io_pipe_phv_in_data_80; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_109 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_81 : io_pipe_phv_in_data_81; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_110 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_82 : io_pipe_phv_in_data_82; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_111 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_83 : io_pipe_phv_in_data_83; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_112 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_84 : io_pipe_phv_in_data_84; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_113 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_85 : io_pipe_phv_in_data_85; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_114 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_86 : io_pipe_phv_in_data_86; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_115 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_87 : io_pipe_phv_in_data_87; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_116 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_88 : io_pipe_phv_in_data_88; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_117 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_89 : io_pipe_phv_in_data_89; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_118 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_90 : io_pipe_phv_in_data_90; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_119 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_91 : io_pipe_phv_in_data_91; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_120 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_92 : io_pipe_phv_in_data_92; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_121 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_93 : io_pipe_phv_in_data_93; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_122 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_94 : io_pipe_phv_in_data_94; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_123 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_95 : io_pipe_phv_in_data_95; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_124 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_96 : io_pipe_phv_in_data_96; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_125 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_97 : io_pipe_phv_in_data_97; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_126 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_98 : io_pipe_phv_in_data_98; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_127 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_99 : io_pipe_phv_in_data_99; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_128 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_100 : io_pipe_phv_in_data_100; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_129 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_101 : io_pipe_phv_in_data_101; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_130 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_102 : io_pipe_phv_in_data_102; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_131 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_103 : io_pipe_phv_in_data_103; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_132 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_104 : io_pipe_phv_in_data_104; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_133 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_105 : io_pipe_phv_in_data_105; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_134 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_106 : io_pipe_phv_in_data_106; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_135 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_107 : io_pipe_phv_in_data_107; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_136 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_108 : io_pipe_phv_in_data_108; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_137 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_109 : io_pipe_phv_in_data_109; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_138 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_110 : io_pipe_phv_in_data_110; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_139 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_111 : io_pipe_phv_in_data_111; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_140 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_112 : io_pipe_phv_in_data_112; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_141 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_113 : io_pipe_phv_in_data_113; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_142 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_114 : io_pipe_phv_in_data_114; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_143 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_115 : io_pipe_phv_in_data_115; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_144 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_116 : io_pipe_phv_in_data_116; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_145 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_117 : io_pipe_phv_in_data_117; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_146 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_118 : io_pipe_phv_in_data_118; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_147 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_119 : io_pipe_phv_in_data_119; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_148 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_120 : io_pipe_phv_in_data_120; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_149 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_121 : io_pipe_phv_in_data_121; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_150 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_122 : io_pipe_phv_in_data_122; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_151 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_123 : io_pipe_phv_in_data_123; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_152 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_124 : io_pipe_phv_in_data_124; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_153 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_125 : io_pipe_phv_in_data_125; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_154 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_126 : io_pipe_phv_in_data_126; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_155 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_127 : io_pipe_phv_in_data_127; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_156 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_128 : io_pipe_phv_in_data_128; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_157 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_129 : io_pipe_phv_in_data_129; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_158 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_130 : io_pipe_phv_in_data_130; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_159 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_131 : io_pipe_phv_in_data_131; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_160 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_132 : io_pipe_phv_in_data_132; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_161 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_133 : io_pipe_phv_in_data_133; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_162 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_134 : io_pipe_phv_in_data_134; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_163 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_135 : io_pipe_phv_in_data_135; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_164 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_136 : io_pipe_phv_in_data_136; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_165 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_137 : io_pipe_phv_in_data_137; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_166 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_138 : io_pipe_phv_in_data_138; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_167 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_139 : io_pipe_phv_in_data_139; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_168 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_140 : io_pipe_phv_in_data_140; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_169 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_141 : io_pipe_phv_in_data_141; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_170 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_142 : io_pipe_phv_in_data_142; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_171 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_143 : io_pipe_phv_in_data_143; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_172 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_144 : io_pipe_phv_in_data_144; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_173 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_145 : io_pipe_phv_in_data_145; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_174 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_146 : io_pipe_phv_in_data_146; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_175 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_147 : io_pipe_phv_in_data_147; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_176 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_148 : io_pipe_phv_in_data_148; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_177 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_149 : io_pipe_phv_in_data_149; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_178 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_150 : io_pipe_phv_in_data_150; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_179 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_151 : io_pipe_phv_in_data_151; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_180 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_152 : io_pipe_phv_in_data_152; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_181 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_153 : io_pipe_phv_in_data_153; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_182 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_154 : io_pipe_phv_in_data_154; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_183 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_155 : io_pipe_phv_in_data_155; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_184 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_156 : io_pipe_phv_in_data_156; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_185 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_157 : io_pipe_phv_in_data_157; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_186 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_158 : io_pipe_phv_in_data_158; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_187 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_159 : io_pipe_phv_in_data_159; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_188 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_160 : io_pipe_phv_in_data_160; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_189 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_161 : io_pipe_phv_in_data_161; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_190 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_162 : io_pipe_phv_in_data_162; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_191 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_163 : io_pipe_phv_in_data_163; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_192 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_164 : io_pipe_phv_in_data_164; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_193 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_165 : io_pipe_phv_in_data_165; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_194 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_166 : io_pipe_phv_in_data_166; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_195 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_167 : io_pipe_phv_in_data_167; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_196 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_168 : io_pipe_phv_in_data_168; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_197 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_169 : io_pipe_phv_in_data_169; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_198 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_170 : io_pipe_phv_in_data_170; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_199 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_171 : io_pipe_phv_in_data_171; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_200 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_172 : io_pipe_phv_in_data_172; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_201 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_173 : io_pipe_phv_in_data_173; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_202 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_174 : io_pipe_phv_in_data_174; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_203 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_175 : io_pipe_phv_in_data_175; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_204 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_176 : io_pipe_phv_in_data_176; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_205 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_177 : io_pipe_phv_in_data_177; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_206 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_178 : io_pipe_phv_in_data_178; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_207 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_179 : io_pipe_phv_in_data_179; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_208 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_180 : io_pipe_phv_in_data_180; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_209 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_181 : io_pipe_phv_in_data_181; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_210 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_182 : io_pipe_phv_in_data_182; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_211 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_183 : io_pipe_phv_in_data_183; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_212 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_184 : io_pipe_phv_in_data_184; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_213 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_185 : io_pipe_phv_in_data_185; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_214 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_186 : io_pipe_phv_in_data_186; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_215 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_187 : io_pipe_phv_in_data_187; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_216 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_188 : io_pipe_phv_in_data_188; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_217 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_189 : io_pipe_phv_in_data_189; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_218 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_190 : io_pipe_phv_in_data_190; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_219 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_191 : io_pipe_phv_in_data_191; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_220 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_192 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_221 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_193 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_222 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_194 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_223 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_195 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_224 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_196 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_225 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_197 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_226 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_198 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_227 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_199 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_228 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_200 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_229 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_201 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_230 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_202 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_231 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_203 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_232 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_204 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_233 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_205 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_234 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_206 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_235 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_207 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_236 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_208 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_237 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_209 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_238 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_210 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_239 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_211 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_240 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_212 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_241 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_213 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_242 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_214 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_243 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_215 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_244 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_216 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_245 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_217 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_246 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_218 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_247 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_219 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_248 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_220 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_249 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_221 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_250 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_222 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_251 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_223 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_252 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_224 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_253 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_225 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_254 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_226 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_255 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_227 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_256 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_228 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_257 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_229 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_258 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_230 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_259 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_231 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_260 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_232 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_261 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_233 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_262 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_234 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_263 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_235 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_264 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_236 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_265 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_237 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_266 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_238 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_267 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_239 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_268 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_240 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_269 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_241 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_270 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_242 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_271 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_243 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_272 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_244 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_273 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_245 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_274 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_246 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_275 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_247 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_276 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_248 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_277 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_249 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_278 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_250 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_279 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_251 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_280 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_252 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_281 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_253 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_282 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_254 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_283 = 2'h0 == last_proc_id ? trans_0_io_pipe_phv_out_data_255 : 8'h0; // @[ipsa.scala 96:65 ipsa.scala 97:29 ipsa.scala 92:21]
  wire [7:0] _GEN_306 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_0 : _GEN_28; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_307 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_1 : _GEN_29; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_308 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_2 : _GEN_30; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_309 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_3 : _GEN_31; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_310 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_4 : _GEN_32; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_311 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_5 : _GEN_33; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_312 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_6 : _GEN_34; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_313 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_7 : _GEN_35; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_314 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_8 : _GEN_36; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_315 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_9 : _GEN_37; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_316 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_10 : _GEN_38; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_317 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_11 : _GEN_39; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_318 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_12 : _GEN_40; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_319 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_13 : _GEN_41; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_320 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_14 : _GEN_42; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_321 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_15 : _GEN_43; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_322 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_16 : _GEN_44; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_323 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_17 : _GEN_45; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_324 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_18 : _GEN_46; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_325 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_19 : _GEN_47; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_326 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_20 : _GEN_48; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_327 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_21 : _GEN_49; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_328 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_22 : _GEN_50; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_329 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_23 : _GEN_51; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_330 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_24 : _GEN_52; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_331 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_25 : _GEN_53; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_332 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_26 : _GEN_54; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_333 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_27 : _GEN_55; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_334 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_28 : _GEN_56; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_335 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_29 : _GEN_57; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_336 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_30 : _GEN_58; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_337 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_31 : _GEN_59; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_338 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_32 : _GEN_60; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_339 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_33 : _GEN_61; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_340 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_34 : _GEN_62; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_341 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_35 : _GEN_63; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_342 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_36 : _GEN_64; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_343 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_37 : _GEN_65; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_344 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_38 : _GEN_66; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_345 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_39 : _GEN_67; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_346 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_40 : _GEN_68; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_347 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_41 : _GEN_69; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_348 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_42 : _GEN_70; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_349 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_43 : _GEN_71; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_350 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_44 : _GEN_72; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_351 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_45 : _GEN_73; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_352 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_46 : _GEN_74; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_353 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_47 : _GEN_75; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_354 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_48 : _GEN_76; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_355 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_49 : _GEN_77; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_356 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_50 : _GEN_78; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_357 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_51 : _GEN_79; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_358 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_52 : _GEN_80; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_359 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_53 : _GEN_81; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_360 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_54 : _GEN_82; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_361 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_55 : _GEN_83; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_362 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_56 : _GEN_84; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_363 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_57 : _GEN_85; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_364 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_58 : _GEN_86; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_365 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_59 : _GEN_87; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_366 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_60 : _GEN_88; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_367 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_61 : _GEN_89; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_368 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_62 : _GEN_90; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_369 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_63 : _GEN_91; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_370 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_64 : _GEN_92; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_371 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_65 : _GEN_93; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_372 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_66 : _GEN_94; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_373 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_67 : _GEN_95; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_374 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_68 : _GEN_96; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_375 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_69 : _GEN_97; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_376 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_70 : _GEN_98; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_377 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_71 : _GEN_99; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_378 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_72 : _GEN_100; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_379 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_73 : _GEN_101; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_380 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_74 : _GEN_102; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_381 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_75 : _GEN_103; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_382 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_76 : _GEN_104; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_383 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_77 : _GEN_105; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_384 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_78 : _GEN_106; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_385 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_79 : _GEN_107; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_386 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_80 : _GEN_108; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_387 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_81 : _GEN_109; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_388 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_82 : _GEN_110; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_389 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_83 : _GEN_111; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_390 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_84 : _GEN_112; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_391 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_85 : _GEN_113; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_392 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_86 : _GEN_114; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_393 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_87 : _GEN_115; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_394 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_88 : _GEN_116; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_395 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_89 : _GEN_117; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_396 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_90 : _GEN_118; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_397 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_91 : _GEN_119; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_398 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_92 : _GEN_120; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_399 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_93 : _GEN_121; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_400 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_94 : _GEN_122; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_401 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_95 : _GEN_123; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_402 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_96 : _GEN_124; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_403 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_97 : _GEN_125; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_404 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_98 : _GEN_126; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_405 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_99 : _GEN_127; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_406 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_100 : _GEN_128; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_407 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_101 : _GEN_129; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_408 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_102 : _GEN_130; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_409 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_103 : _GEN_131; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_410 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_104 : _GEN_132; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_411 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_105 : _GEN_133; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_412 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_106 : _GEN_134; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_413 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_107 : _GEN_135; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_414 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_108 : _GEN_136; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_415 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_109 : _GEN_137; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_416 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_110 : _GEN_138; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_417 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_111 : _GEN_139; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_418 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_112 : _GEN_140; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_419 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_113 : _GEN_141; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_420 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_114 : _GEN_142; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_421 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_115 : _GEN_143; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_422 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_116 : _GEN_144; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_423 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_117 : _GEN_145; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_424 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_118 : _GEN_146; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_425 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_119 : _GEN_147; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_426 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_120 : _GEN_148; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_427 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_121 : _GEN_149; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_428 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_122 : _GEN_150; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_429 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_123 : _GEN_151; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_430 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_124 : _GEN_152; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_431 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_125 : _GEN_153; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_432 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_126 : _GEN_154; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_433 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_127 : _GEN_155; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_434 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_128 : _GEN_156; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_435 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_129 : _GEN_157; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_436 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_130 : _GEN_158; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_437 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_131 : _GEN_159; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_438 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_132 : _GEN_160; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_439 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_133 : _GEN_161; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_440 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_134 : _GEN_162; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_441 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_135 : _GEN_163; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_442 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_136 : _GEN_164; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_443 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_137 : _GEN_165; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_444 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_138 : _GEN_166; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_445 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_139 : _GEN_167; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_446 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_140 : _GEN_168; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_447 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_141 : _GEN_169; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_448 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_142 : _GEN_170; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_449 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_143 : _GEN_171; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_450 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_144 : _GEN_172; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_451 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_145 : _GEN_173; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_452 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_146 : _GEN_174; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_453 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_147 : _GEN_175; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_454 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_148 : _GEN_176; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_455 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_149 : _GEN_177; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_456 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_150 : _GEN_178; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_457 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_151 : _GEN_179; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_458 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_152 : _GEN_180; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_459 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_153 : _GEN_181; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_460 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_154 : _GEN_182; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_461 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_155 : _GEN_183; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_462 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_156 : _GEN_184; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_463 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_157 : _GEN_185; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_464 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_158 : _GEN_186; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_465 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_159 : _GEN_187; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_466 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_160 : _GEN_188; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_467 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_161 : _GEN_189; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_468 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_162 : _GEN_190; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_469 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_163 : _GEN_191; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_470 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_164 : _GEN_192; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_471 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_165 : _GEN_193; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_472 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_166 : _GEN_194; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_473 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_167 : _GEN_195; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_474 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_168 : _GEN_196; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_475 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_169 : _GEN_197; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_476 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_170 : _GEN_198; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_477 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_171 : _GEN_199; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_478 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_172 : _GEN_200; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_479 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_173 : _GEN_201; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_480 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_174 : _GEN_202; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_481 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_175 : _GEN_203; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_482 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_176 : _GEN_204; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_483 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_177 : _GEN_205; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_484 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_178 : _GEN_206; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_485 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_179 : _GEN_207; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_486 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_180 : _GEN_208; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_487 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_181 : _GEN_209; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_488 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_182 : _GEN_210; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_489 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_183 : _GEN_211; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_490 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_184 : _GEN_212; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_491 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_185 : _GEN_213; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_492 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_186 : _GEN_214; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_493 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_187 : _GEN_215; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_494 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_188 : _GEN_216; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_495 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_189 : _GEN_217; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_496 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_190 : _GEN_218; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_497 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_191 : _GEN_219; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_498 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_192 : _GEN_220; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_499 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_193 : _GEN_221; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_500 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_194 : _GEN_222; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_501 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_195 : _GEN_223; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_502 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_196 : _GEN_224; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_503 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_197 : _GEN_225; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_504 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_198 : _GEN_226; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_505 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_199 : _GEN_227; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_506 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_200 : _GEN_228; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_507 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_201 : _GEN_229; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_508 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_202 : _GEN_230; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_509 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_203 : _GEN_231; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_510 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_204 : _GEN_232; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_511 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_205 : _GEN_233; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_512 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_206 : _GEN_234; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_513 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_207 : _GEN_235; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_514 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_208 : _GEN_236; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_515 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_209 : _GEN_237; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_516 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_210 : _GEN_238; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_517 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_211 : _GEN_239; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_518 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_212 : _GEN_240; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_519 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_213 : _GEN_241; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_520 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_214 : _GEN_242; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_521 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_215 : _GEN_243; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_522 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_216 : _GEN_244; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_523 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_217 : _GEN_245; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_524 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_218 : _GEN_246; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_525 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_219 : _GEN_247; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_526 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_220 : _GEN_248; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_527 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_221 : _GEN_249; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_528 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_222 : _GEN_250; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_529 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_223 : _GEN_251; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_530 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_224 : _GEN_252; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_531 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_225 : _GEN_253; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_532 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_226 : _GEN_254; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_533 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_227 : _GEN_255; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_534 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_228 : _GEN_256; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_535 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_229 : _GEN_257; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_536 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_230 : _GEN_258; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_537 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_231 : _GEN_259; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_538 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_232 : _GEN_260; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_539 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_233 : _GEN_261; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_540 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_234 : _GEN_262; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_541 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_235 : _GEN_263; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_542 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_236 : _GEN_264; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_543 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_237 : _GEN_265; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_544 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_238 : _GEN_266; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_545 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_239 : _GEN_267; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_546 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_240 : _GEN_268; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_547 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_241 : _GEN_269; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_548 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_242 : _GEN_270; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_549 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_243 : _GEN_271; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_550 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_244 : _GEN_272; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_551 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_245 : _GEN_273; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_552 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_246 : _GEN_274; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_553 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_247 : _GEN_275; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_554 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_248 : _GEN_276; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_555 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_249 : _GEN_277; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_556 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_250 : _GEN_278; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_557 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_251 : _GEN_279; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_558 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_252 : _GEN_280; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_559 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_253 : _GEN_281; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_560 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_254 : _GEN_282; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_561 = 2'h1 == last_proc_id ? trans_1_io_pipe_phv_out_data_255 : _GEN_283; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_584 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_0 : _GEN_306; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_585 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_1 : _GEN_307; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_586 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_2 : _GEN_308; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_587 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_3 : _GEN_309; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_588 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_4 : _GEN_310; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_589 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_5 : _GEN_311; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_590 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_6 : _GEN_312; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_591 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_7 : _GEN_313; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_592 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_8 : _GEN_314; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_593 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_9 : _GEN_315; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_594 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_10 : _GEN_316; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_595 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_11 : _GEN_317; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_596 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_12 : _GEN_318; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_597 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_13 : _GEN_319; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_598 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_14 : _GEN_320; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_599 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_15 : _GEN_321; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_600 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_16 : _GEN_322; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_601 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_17 : _GEN_323; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_602 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_18 : _GEN_324; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_603 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_19 : _GEN_325; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_604 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_20 : _GEN_326; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_605 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_21 : _GEN_327; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_606 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_22 : _GEN_328; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_607 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_23 : _GEN_329; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_608 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_24 : _GEN_330; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_609 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_25 : _GEN_331; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_610 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_26 : _GEN_332; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_611 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_27 : _GEN_333; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_612 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_28 : _GEN_334; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_613 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_29 : _GEN_335; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_614 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_30 : _GEN_336; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_615 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_31 : _GEN_337; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_616 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_32 : _GEN_338; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_617 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_33 : _GEN_339; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_618 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_34 : _GEN_340; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_619 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_35 : _GEN_341; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_620 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_36 : _GEN_342; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_621 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_37 : _GEN_343; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_622 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_38 : _GEN_344; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_623 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_39 : _GEN_345; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_624 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_40 : _GEN_346; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_625 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_41 : _GEN_347; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_626 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_42 : _GEN_348; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_627 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_43 : _GEN_349; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_628 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_44 : _GEN_350; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_629 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_45 : _GEN_351; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_630 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_46 : _GEN_352; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_631 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_47 : _GEN_353; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_632 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_48 : _GEN_354; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_633 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_49 : _GEN_355; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_634 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_50 : _GEN_356; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_635 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_51 : _GEN_357; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_636 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_52 : _GEN_358; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_637 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_53 : _GEN_359; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_638 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_54 : _GEN_360; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_639 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_55 : _GEN_361; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_640 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_56 : _GEN_362; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_641 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_57 : _GEN_363; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_642 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_58 : _GEN_364; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_643 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_59 : _GEN_365; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_644 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_60 : _GEN_366; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_645 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_61 : _GEN_367; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_646 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_62 : _GEN_368; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_647 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_63 : _GEN_369; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_648 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_64 : _GEN_370; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_649 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_65 : _GEN_371; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_650 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_66 : _GEN_372; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_651 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_67 : _GEN_373; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_652 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_68 : _GEN_374; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_653 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_69 : _GEN_375; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_654 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_70 : _GEN_376; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_655 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_71 : _GEN_377; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_656 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_72 : _GEN_378; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_657 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_73 : _GEN_379; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_658 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_74 : _GEN_380; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_659 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_75 : _GEN_381; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_660 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_76 : _GEN_382; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_661 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_77 : _GEN_383; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_662 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_78 : _GEN_384; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_663 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_79 : _GEN_385; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_664 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_80 : _GEN_386; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_665 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_81 : _GEN_387; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_666 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_82 : _GEN_388; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_667 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_83 : _GEN_389; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_668 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_84 : _GEN_390; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_669 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_85 : _GEN_391; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_670 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_86 : _GEN_392; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_671 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_87 : _GEN_393; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_672 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_88 : _GEN_394; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_673 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_89 : _GEN_395; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_674 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_90 : _GEN_396; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_675 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_91 : _GEN_397; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_676 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_92 : _GEN_398; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_677 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_93 : _GEN_399; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_678 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_94 : _GEN_400; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_679 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_95 : _GEN_401; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_680 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_96 : _GEN_402; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_681 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_97 : _GEN_403; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_682 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_98 : _GEN_404; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_683 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_99 : _GEN_405; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_684 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_100 : _GEN_406; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_685 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_101 : _GEN_407; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_686 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_102 : _GEN_408; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_687 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_103 : _GEN_409; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_688 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_104 : _GEN_410; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_689 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_105 : _GEN_411; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_690 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_106 : _GEN_412; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_691 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_107 : _GEN_413; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_692 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_108 : _GEN_414; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_693 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_109 : _GEN_415; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_694 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_110 : _GEN_416; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_695 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_111 : _GEN_417; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_696 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_112 : _GEN_418; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_697 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_113 : _GEN_419; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_698 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_114 : _GEN_420; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_699 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_115 : _GEN_421; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_700 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_116 : _GEN_422; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_701 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_117 : _GEN_423; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_702 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_118 : _GEN_424; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_703 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_119 : _GEN_425; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_704 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_120 : _GEN_426; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_705 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_121 : _GEN_427; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_706 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_122 : _GEN_428; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_707 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_123 : _GEN_429; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_708 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_124 : _GEN_430; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_709 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_125 : _GEN_431; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_710 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_126 : _GEN_432; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_711 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_127 : _GEN_433; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_712 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_128 : _GEN_434; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_713 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_129 : _GEN_435; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_714 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_130 : _GEN_436; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_715 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_131 : _GEN_437; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_716 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_132 : _GEN_438; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_717 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_133 : _GEN_439; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_718 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_134 : _GEN_440; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_719 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_135 : _GEN_441; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_720 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_136 : _GEN_442; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_721 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_137 : _GEN_443; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_722 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_138 : _GEN_444; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_723 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_139 : _GEN_445; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_724 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_140 : _GEN_446; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_725 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_141 : _GEN_447; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_726 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_142 : _GEN_448; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_727 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_143 : _GEN_449; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_728 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_144 : _GEN_450; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_729 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_145 : _GEN_451; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_730 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_146 : _GEN_452; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_731 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_147 : _GEN_453; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_732 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_148 : _GEN_454; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_733 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_149 : _GEN_455; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_734 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_150 : _GEN_456; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_735 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_151 : _GEN_457; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_736 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_152 : _GEN_458; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_737 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_153 : _GEN_459; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_738 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_154 : _GEN_460; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_739 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_155 : _GEN_461; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_740 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_156 : _GEN_462; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_741 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_157 : _GEN_463; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_742 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_158 : _GEN_464; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_743 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_159 : _GEN_465; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_744 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_160 : _GEN_466; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_745 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_161 : _GEN_467; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_746 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_162 : _GEN_468; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_747 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_163 : _GEN_469; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_748 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_164 : _GEN_470; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_749 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_165 : _GEN_471; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_750 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_166 : _GEN_472; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_751 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_167 : _GEN_473; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_752 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_168 : _GEN_474; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_753 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_169 : _GEN_475; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_754 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_170 : _GEN_476; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_755 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_171 : _GEN_477; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_756 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_172 : _GEN_478; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_757 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_173 : _GEN_479; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_758 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_174 : _GEN_480; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_759 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_175 : _GEN_481; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_760 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_176 : _GEN_482; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_761 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_177 : _GEN_483; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_762 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_178 : _GEN_484; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_763 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_179 : _GEN_485; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_764 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_180 : _GEN_486; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_765 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_181 : _GEN_487; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_766 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_182 : _GEN_488; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_767 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_183 : _GEN_489; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_768 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_184 : _GEN_490; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_769 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_185 : _GEN_491; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_770 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_186 : _GEN_492; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_771 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_187 : _GEN_493; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_772 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_188 : _GEN_494; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_773 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_189 : _GEN_495; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_774 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_190 : _GEN_496; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_775 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_191 : _GEN_497; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_776 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_192 : _GEN_498; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_777 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_193 : _GEN_499; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_778 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_194 : _GEN_500; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_779 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_195 : _GEN_501; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_780 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_196 : _GEN_502; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_781 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_197 : _GEN_503; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_782 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_198 : _GEN_504; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_783 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_199 : _GEN_505; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_784 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_200 : _GEN_506; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_785 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_201 : _GEN_507; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_786 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_202 : _GEN_508; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_787 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_203 : _GEN_509; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_788 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_204 : _GEN_510; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_789 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_205 : _GEN_511; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_790 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_206 : _GEN_512; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_791 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_207 : _GEN_513; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_792 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_208 : _GEN_514; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_793 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_209 : _GEN_515; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_794 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_210 : _GEN_516; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_795 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_211 : _GEN_517; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_796 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_212 : _GEN_518; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_797 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_213 : _GEN_519; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_798 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_214 : _GEN_520; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_799 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_215 : _GEN_521; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_800 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_216 : _GEN_522; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_801 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_217 : _GEN_523; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_802 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_218 : _GEN_524; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_803 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_219 : _GEN_525; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_804 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_220 : _GEN_526; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_805 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_221 : _GEN_527; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_806 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_222 : _GEN_528; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_807 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_223 : _GEN_529; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_808 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_224 : _GEN_530; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_809 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_225 : _GEN_531; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_810 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_226 : _GEN_532; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_811 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_227 : _GEN_533; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_812 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_228 : _GEN_534; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_813 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_229 : _GEN_535; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_814 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_230 : _GEN_536; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_815 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_231 : _GEN_537; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_816 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_232 : _GEN_538; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_817 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_233 : _GEN_539; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_818 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_234 : _GEN_540; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_819 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_235 : _GEN_541; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_820 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_236 : _GEN_542; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_821 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_237 : _GEN_543; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_822 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_238 : _GEN_544; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_823 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_239 : _GEN_545; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_824 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_240 : _GEN_546; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_825 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_241 : _GEN_547; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_826 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_242 : _GEN_548; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_827 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_243 : _GEN_549; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_828 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_244 : _GEN_550; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_829 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_245 : _GEN_551; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_830 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_246 : _GEN_552; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_831 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_247 : _GEN_553; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_832 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_248 : _GEN_554; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_833 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_249 : _GEN_555; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_834 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_250 : _GEN_556; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_835 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_251 : _GEN_557; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_836 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_252 : _GEN_558; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_837 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_253 : _GEN_559; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_838 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_254 : _GEN_560; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  wire [7:0] _GEN_839 = 2'h2 == last_proc_id ? trans_2_io_pipe_phv_out_data_255 : _GEN_561; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  reg [7:0] amplifier_0_0_data_0; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_1; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_2; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_3; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_4; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_5; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_6; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_7; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_8; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_9; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_10; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_11; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_12; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_13; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_14; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_15; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_16; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_17; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_18; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_19; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_20; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_21; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_22; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_23; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_24; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_25; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_26; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_27; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_28; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_29; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_30; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_31; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_32; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_33; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_34; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_35; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_36; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_37; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_38; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_39; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_40; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_41; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_42; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_43; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_44; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_45; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_46; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_47; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_48; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_49; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_50; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_51; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_52; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_53; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_54; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_55; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_56; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_57; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_58; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_59; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_60; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_61; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_62; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_63; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_64; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_65; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_66; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_67; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_68; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_69; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_70; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_71; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_72; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_73; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_74; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_75; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_76; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_77; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_78; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_79; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_80; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_81; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_82; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_83; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_84; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_85; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_86; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_87; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_88; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_89; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_90; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_91; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_92; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_93; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_94; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_95; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_96; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_97; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_98; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_99; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_100; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_101; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_102; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_103; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_104; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_105; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_106; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_107; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_108; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_109; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_110; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_111; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_112; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_113; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_114; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_115; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_116; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_117; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_118; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_119; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_120; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_121; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_122; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_123; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_124; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_125; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_126; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_127; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_128; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_129; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_130; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_131; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_132; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_133; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_134; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_135; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_136; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_137; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_138; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_139; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_140; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_141; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_142; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_143; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_144; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_145; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_146; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_147; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_148; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_149; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_150; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_151; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_152; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_153; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_154; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_155; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_156; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_157; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_158; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_159; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_160; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_161; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_162; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_163; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_164; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_165; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_166; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_167; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_168; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_169; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_170; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_171; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_172; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_173; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_174; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_175; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_176; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_177; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_178; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_179; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_180; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_181; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_182; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_183; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_184; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_185; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_186; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_187; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_188; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_189; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_190; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_191; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_192; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_193; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_194; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_195; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_196; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_197; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_198; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_199; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_200; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_201; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_202; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_203; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_204; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_205; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_206; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_207; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_208; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_209; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_210; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_211; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_212; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_213; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_214; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_215; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_216; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_217; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_218; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_219; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_220; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_221; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_222; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_223; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_224; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_225; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_226; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_227; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_228; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_229; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_230; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_231; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_232; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_233; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_234; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_235; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_236; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_237; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_238; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_239; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_240; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_241; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_242; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_243; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_244; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_245; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_246; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_247; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_248; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_249; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_250; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_251; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_252; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_253; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_254; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_data_255; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_0_header_0; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_0_header_1; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_0_header_2; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_0_header_3; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_0_header_4; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_0_header_5; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_0_header_6; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_0_header_7; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_0_header_8; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_0_header_9; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_0_header_10; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_0_header_11; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_0_header_12; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_0_header_13; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_0_header_14; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_0_header_15; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_parse_current_state; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_0_parse_current_offset; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_0_parse_transition_field; // @[ipsa.scala 103:24]
  reg [1:0] amplifier_0_0_next_processor_id; // @[ipsa.scala 103:24]
  reg  amplifier_0_0_next_config_id; // @[ipsa.scala 103:24]
  reg  amplifier_0_0_is_valid_processor; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_0; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_1; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_2; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_3; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_4; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_5; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_6; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_7; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_8; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_9; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_10; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_11; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_12; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_13; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_14; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_15; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_16; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_17; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_18; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_19; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_20; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_21; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_22; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_23; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_24; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_25; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_26; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_27; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_28; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_29; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_30; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_31; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_32; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_33; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_34; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_35; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_36; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_37; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_38; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_39; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_40; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_41; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_42; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_43; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_44; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_45; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_46; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_47; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_48; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_49; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_50; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_51; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_52; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_53; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_54; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_55; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_56; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_57; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_58; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_59; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_60; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_61; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_62; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_63; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_64; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_65; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_66; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_67; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_68; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_69; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_70; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_71; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_72; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_73; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_74; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_75; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_76; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_77; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_78; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_79; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_80; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_81; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_82; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_83; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_84; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_85; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_86; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_87; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_88; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_89; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_90; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_91; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_92; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_93; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_94; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_95; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_96; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_97; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_98; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_99; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_100; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_101; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_102; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_103; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_104; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_105; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_106; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_107; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_108; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_109; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_110; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_111; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_112; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_113; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_114; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_115; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_116; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_117; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_118; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_119; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_120; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_121; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_122; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_123; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_124; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_125; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_126; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_127; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_128; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_129; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_130; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_131; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_132; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_133; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_134; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_135; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_136; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_137; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_138; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_139; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_140; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_141; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_142; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_143; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_144; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_145; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_146; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_147; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_148; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_149; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_150; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_151; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_152; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_153; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_154; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_155; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_156; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_157; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_158; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_159; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_160; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_161; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_162; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_163; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_164; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_165; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_166; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_167; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_168; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_169; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_170; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_171; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_172; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_173; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_174; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_175; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_176; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_177; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_178; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_179; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_180; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_181; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_182; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_183; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_184; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_185; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_186; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_187; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_188; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_189; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_190; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_191; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_192; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_193; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_194; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_195; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_196; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_197; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_198; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_199; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_200; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_201; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_202; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_203; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_204; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_205; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_206; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_207; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_208; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_209; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_210; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_211; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_212; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_213; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_214; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_215; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_216; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_217; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_218; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_219; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_220; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_221; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_222; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_223; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_224; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_225; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_226; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_227; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_228; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_229; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_230; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_231; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_232; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_233; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_234; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_235; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_236; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_237; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_238; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_239; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_240; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_241; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_242; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_243; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_244; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_245; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_246; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_247; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_248; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_249; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_250; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_251; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_252; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_253; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_254; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_data_255; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_1_header_0; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_1_header_1; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_1_header_2; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_1_header_3; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_1_header_4; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_1_header_5; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_1_header_6; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_1_header_7; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_1_header_8; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_1_header_9; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_1_header_10; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_1_header_11; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_1_header_12; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_1_header_13; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_1_header_14; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_1_header_15; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_parse_current_state; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_1_parse_current_offset; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_1_parse_transition_field; // @[ipsa.scala 103:24]
  reg [1:0] amplifier_0_1_next_processor_id; // @[ipsa.scala 103:24]
  reg  amplifier_0_1_next_config_id; // @[ipsa.scala 103:24]
  reg  amplifier_0_1_is_valid_processor; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_0; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_1; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_2; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_3; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_4; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_5; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_6; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_7; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_8; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_9; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_10; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_11; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_12; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_13; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_14; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_15; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_16; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_17; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_18; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_19; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_20; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_21; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_22; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_23; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_24; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_25; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_26; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_27; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_28; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_29; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_30; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_31; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_32; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_33; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_34; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_35; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_36; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_37; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_38; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_39; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_40; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_41; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_42; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_43; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_44; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_45; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_46; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_47; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_48; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_49; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_50; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_51; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_52; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_53; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_54; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_55; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_56; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_57; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_58; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_59; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_60; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_61; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_62; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_63; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_64; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_65; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_66; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_67; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_68; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_69; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_70; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_71; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_72; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_73; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_74; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_75; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_76; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_77; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_78; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_79; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_80; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_81; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_82; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_83; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_84; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_85; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_86; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_87; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_88; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_89; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_90; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_91; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_92; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_93; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_94; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_95; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_96; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_97; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_98; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_99; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_100; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_101; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_102; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_103; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_104; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_105; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_106; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_107; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_108; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_109; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_110; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_111; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_112; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_113; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_114; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_115; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_116; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_117; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_118; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_119; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_120; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_121; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_122; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_123; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_124; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_125; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_126; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_127; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_128; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_129; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_130; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_131; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_132; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_133; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_134; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_135; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_136; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_137; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_138; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_139; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_140; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_141; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_142; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_143; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_144; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_145; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_146; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_147; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_148; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_149; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_150; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_151; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_152; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_153; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_154; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_155; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_156; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_157; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_158; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_159; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_160; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_161; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_162; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_163; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_164; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_165; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_166; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_167; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_168; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_169; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_170; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_171; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_172; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_173; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_174; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_175; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_176; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_177; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_178; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_179; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_180; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_181; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_182; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_183; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_184; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_185; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_186; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_187; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_188; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_189; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_190; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_191; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_192; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_193; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_194; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_195; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_196; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_197; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_198; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_199; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_200; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_201; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_202; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_203; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_204; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_205; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_206; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_207; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_208; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_209; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_210; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_211; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_212; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_213; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_214; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_215; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_216; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_217; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_218; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_219; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_220; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_221; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_222; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_223; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_224; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_225; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_226; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_227; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_228; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_229; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_230; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_231; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_232; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_233; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_234; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_235; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_236; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_237; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_238; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_239; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_240; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_241; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_242; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_243; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_244; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_245; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_246; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_247; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_248; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_249; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_250; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_251; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_252; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_253; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_254; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_data_255; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_2_header_0; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_2_header_1; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_2_header_2; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_2_header_3; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_2_header_4; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_2_header_5; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_2_header_6; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_2_header_7; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_2_header_8; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_2_header_9; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_2_header_10; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_2_header_11; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_2_header_12; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_2_header_13; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_2_header_14; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_2_header_15; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_parse_current_state; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_2_parse_current_offset; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_2_parse_transition_field; // @[ipsa.scala 103:24]
  reg [1:0] amplifier_0_2_next_processor_id; // @[ipsa.scala 103:24]
  reg  amplifier_0_2_next_config_id; // @[ipsa.scala 103:24]
  reg  amplifier_0_2_is_valid_processor; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_0; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_1; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_2; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_3; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_4; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_5; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_6; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_7; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_8; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_9; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_10; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_11; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_12; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_13; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_14; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_15; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_16; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_17; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_18; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_19; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_20; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_21; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_22; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_23; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_24; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_25; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_26; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_27; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_28; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_29; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_30; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_31; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_32; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_33; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_34; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_35; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_36; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_37; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_38; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_39; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_40; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_41; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_42; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_43; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_44; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_45; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_46; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_47; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_48; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_49; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_50; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_51; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_52; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_53; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_54; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_55; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_56; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_57; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_58; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_59; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_60; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_61; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_62; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_63; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_64; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_65; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_66; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_67; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_68; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_69; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_70; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_71; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_72; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_73; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_74; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_75; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_76; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_77; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_78; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_79; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_80; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_81; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_82; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_83; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_84; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_85; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_86; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_87; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_88; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_89; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_90; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_91; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_92; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_93; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_94; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_95; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_96; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_97; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_98; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_99; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_100; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_101; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_102; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_103; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_104; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_105; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_106; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_107; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_108; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_109; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_110; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_111; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_112; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_113; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_114; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_115; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_116; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_117; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_118; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_119; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_120; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_121; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_122; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_123; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_124; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_125; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_126; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_127; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_128; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_129; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_130; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_131; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_132; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_133; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_134; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_135; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_136; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_137; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_138; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_139; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_140; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_141; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_142; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_143; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_144; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_145; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_146; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_147; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_148; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_149; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_150; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_151; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_152; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_153; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_154; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_155; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_156; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_157; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_158; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_159; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_160; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_161; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_162; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_163; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_164; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_165; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_166; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_167; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_168; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_169; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_170; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_171; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_172; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_173; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_174; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_175; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_176; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_177; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_178; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_179; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_180; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_181; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_182; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_183; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_184; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_185; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_186; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_187; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_188; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_189; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_190; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_191; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_192; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_193; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_194; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_195; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_196; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_197; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_198; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_199; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_200; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_201; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_202; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_203; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_204; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_205; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_206; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_207; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_208; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_209; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_210; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_211; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_212; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_213; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_214; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_215; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_216; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_217; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_218; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_219; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_220; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_221; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_222; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_223; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_224; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_225; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_226; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_227; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_228; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_229; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_230; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_231; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_232; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_233; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_234; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_235; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_236; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_237; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_238; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_239; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_240; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_241; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_242; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_243; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_244; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_245; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_246; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_247; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_248; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_249; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_250; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_251; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_252; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_253; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_254; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_data_255; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_3_header_0; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_3_header_1; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_3_header_2; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_3_header_3; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_3_header_4; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_3_header_5; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_3_header_6; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_3_header_7; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_3_header_8; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_3_header_9; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_3_header_10; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_3_header_11; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_3_header_12; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_3_header_13; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_3_header_14; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_3_header_15; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_parse_current_state; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_0_3_parse_current_offset; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_0_3_parse_transition_field; // @[ipsa.scala 103:24]
  reg [1:0] amplifier_0_3_next_processor_id; // @[ipsa.scala 103:24]
  reg  amplifier_0_3_next_config_id; // @[ipsa.scala 103:24]
  reg  amplifier_0_3_is_valid_processor; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_0; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_1; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_2; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_3; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_4; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_5; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_6; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_7; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_8; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_9; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_10; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_11; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_12; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_13; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_14; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_15; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_16; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_17; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_18; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_19; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_20; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_21; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_22; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_23; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_24; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_25; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_26; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_27; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_28; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_29; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_30; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_31; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_32; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_33; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_34; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_35; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_36; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_37; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_38; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_39; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_40; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_41; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_42; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_43; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_44; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_45; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_46; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_47; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_48; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_49; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_50; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_51; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_52; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_53; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_54; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_55; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_56; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_57; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_58; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_59; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_60; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_61; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_62; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_63; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_64; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_65; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_66; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_67; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_68; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_69; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_70; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_71; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_72; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_73; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_74; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_75; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_76; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_77; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_78; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_79; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_80; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_81; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_82; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_83; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_84; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_85; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_86; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_87; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_88; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_89; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_90; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_91; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_92; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_93; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_94; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_95; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_96; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_97; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_98; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_99; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_100; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_101; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_102; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_103; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_104; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_105; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_106; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_107; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_108; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_109; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_110; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_111; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_112; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_113; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_114; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_115; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_116; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_117; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_118; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_119; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_120; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_121; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_122; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_123; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_124; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_125; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_126; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_127; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_128; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_129; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_130; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_131; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_132; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_133; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_134; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_135; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_136; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_137; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_138; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_139; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_140; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_141; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_142; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_143; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_144; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_145; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_146; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_147; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_148; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_149; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_150; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_151; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_152; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_153; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_154; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_155; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_156; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_157; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_158; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_159; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_160; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_161; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_162; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_163; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_164; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_165; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_166; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_167; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_168; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_169; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_170; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_171; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_172; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_173; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_174; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_175; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_176; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_177; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_178; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_179; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_180; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_181; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_182; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_183; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_184; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_185; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_186; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_187; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_188; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_189; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_190; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_191; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_192; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_193; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_194; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_195; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_196; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_197; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_198; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_199; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_200; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_201; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_202; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_203; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_204; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_205; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_206; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_207; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_208; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_209; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_210; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_211; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_212; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_213; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_214; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_215; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_216; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_217; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_218; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_219; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_220; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_221; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_222; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_223; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_224; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_225; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_226; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_227; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_228; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_229; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_230; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_231; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_232; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_233; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_234; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_235; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_236; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_237; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_238; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_239; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_240; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_241; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_242; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_243; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_244; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_245; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_246; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_247; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_248; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_249; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_250; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_251; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_252; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_253; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_254; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_data_255; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_0_header_0; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_0_header_1; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_0_header_2; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_0_header_3; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_0_header_4; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_0_header_5; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_0_header_6; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_0_header_7; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_0_header_8; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_0_header_9; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_0_header_10; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_0_header_11; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_0_header_12; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_0_header_13; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_0_header_14; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_0_header_15; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_parse_current_state; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_0_parse_current_offset; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_0_parse_transition_field; // @[ipsa.scala 103:24]
  reg [1:0] amplifier_1_0_next_processor_id; // @[ipsa.scala 103:24]
  reg  amplifier_1_0_next_config_id; // @[ipsa.scala 103:24]
  reg  amplifier_1_0_is_valid_processor; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_0; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_1; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_2; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_3; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_4; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_5; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_6; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_7; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_8; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_9; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_10; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_11; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_12; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_13; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_14; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_15; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_16; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_17; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_18; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_19; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_20; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_21; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_22; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_23; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_24; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_25; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_26; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_27; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_28; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_29; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_30; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_31; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_32; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_33; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_34; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_35; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_36; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_37; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_38; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_39; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_40; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_41; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_42; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_43; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_44; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_45; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_46; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_47; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_48; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_49; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_50; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_51; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_52; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_53; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_54; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_55; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_56; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_57; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_58; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_59; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_60; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_61; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_62; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_63; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_64; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_65; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_66; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_67; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_68; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_69; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_70; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_71; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_72; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_73; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_74; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_75; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_76; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_77; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_78; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_79; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_80; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_81; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_82; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_83; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_84; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_85; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_86; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_87; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_88; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_89; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_90; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_91; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_92; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_93; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_94; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_95; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_96; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_97; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_98; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_99; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_100; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_101; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_102; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_103; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_104; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_105; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_106; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_107; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_108; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_109; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_110; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_111; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_112; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_113; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_114; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_115; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_116; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_117; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_118; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_119; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_120; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_121; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_122; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_123; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_124; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_125; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_126; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_127; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_128; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_129; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_130; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_131; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_132; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_133; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_134; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_135; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_136; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_137; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_138; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_139; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_140; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_141; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_142; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_143; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_144; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_145; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_146; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_147; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_148; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_149; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_150; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_151; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_152; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_153; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_154; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_155; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_156; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_157; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_158; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_159; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_160; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_161; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_162; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_163; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_164; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_165; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_166; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_167; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_168; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_169; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_170; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_171; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_172; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_173; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_174; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_175; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_176; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_177; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_178; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_179; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_180; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_181; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_182; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_183; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_184; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_185; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_186; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_187; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_188; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_189; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_190; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_191; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_192; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_193; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_194; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_195; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_196; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_197; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_198; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_199; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_200; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_201; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_202; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_203; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_204; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_205; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_206; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_207; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_208; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_209; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_210; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_211; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_212; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_213; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_214; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_215; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_216; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_217; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_218; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_219; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_220; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_221; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_222; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_223; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_224; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_225; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_226; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_227; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_228; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_229; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_230; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_231; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_232; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_233; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_234; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_235; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_236; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_237; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_238; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_239; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_240; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_241; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_242; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_243; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_244; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_245; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_246; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_247; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_248; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_249; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_250; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_251; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_252; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_253; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_254; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_data_255; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_1_header_0; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_1_header_1; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_1_header_2; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_1_header_3; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_1_header_4; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_1_header_5; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_1_header_6; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_1_header_7; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_1_header_8; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_1_header_9; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_1_header_10; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_1_header_11; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_1_header_12; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_1_header_13; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_1_header_14; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_1_header_15; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_parse_current_state; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_1_parse_current_offset; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_1_parse_transition_field; // @[ipsa.scala 103:24]
  reg [1:0] amplifier_1_1_next_processor_id; // @[ipsa.scala 103:24]
  reg  amplifier_1_1_next_config_id; // @[ipsa.scala 103:24]
  reg  amplifier_1_1_is_valid_processor; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_0; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_1; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_2; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_3; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_4; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_5; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_6; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_7; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_8; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_9; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_10; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_11; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_12; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_13; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_14; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_15; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_16; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_17; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_18; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_19; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_20; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_21; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_22; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_23; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_24; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_25; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_26; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_27; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_28; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_29; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_30; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_31; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_32; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_33; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_34; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_35; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_36; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_37; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_38; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_39; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_40; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_41; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_42; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_43; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_44; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_45; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_46; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_47; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_48; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_49; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_50; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_51; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_52; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_53; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_54; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_55; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_56; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_57; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_58; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_59; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_60; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_61; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_62; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_63; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_64; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_65; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_66; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_67; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_68; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_69; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_70; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_71; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_72; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_73; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_74; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_75; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_76; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_77; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_78; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_79; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_80; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_81; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_82; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_83; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_84; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_85; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_86; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_87; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_88; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_89; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_90; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_91; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_92; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_93; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_94; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_95; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_96; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_97; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_98; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_99; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_100; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_101; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_102; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_103; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_104; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_105; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_106; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_107; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_108; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_109; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_110; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_111; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_112; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_113; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_114; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_115; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_116; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_117; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_118; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_119; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_120; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_121; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_122; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_123; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_124; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_125; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_126; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_127; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_128; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_129; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_130; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_131; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_132; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_133; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_134; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_135; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_136; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_137; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_138; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_139; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_140; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_141; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_142; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_143; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_144; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_145; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_146; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_147; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_148; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_149; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_150; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_151; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_152; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_153; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_154; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_155; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_156; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_157; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_158; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_159; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_160; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_161; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_162; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_163; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_164; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_165; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_166; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_167; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_168; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_169; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_170; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_171; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_172; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_173; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_174; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_175; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_176; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_177; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_178; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_179; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_180; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_181; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_182; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_183; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_184; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_185; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_186; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_187; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_188; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_189; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_190; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_191; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_192; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_193; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_194; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_195; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_196; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_197; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_198; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_199; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_200; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_201; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_202; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_203; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_204; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_205; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_206; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_207; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_208; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_209; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_210; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_211; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_212; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_213; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_214; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_215; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_216; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_217; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_218; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_219; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_220; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_221; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_222; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_223; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_224; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_225; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_226; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_227; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_228; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_229; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_230; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_231; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_232; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_233; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_234; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_235; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_236; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_237; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_238; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_239; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_240; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_241; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_242; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_243; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_244; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_245; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_246; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_247; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_248; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_249; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_250; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_251; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_252; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_253; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_254; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_data_255; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_2_header_0; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_2_header_1; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_2_header_2; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_2_header_3; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_2_header_4; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_2_header_5; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_2_header_6; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_2_header_7; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_2_header_8; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_2_header_9; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_2_header_10; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_2_header_11; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_2_header_12; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_2_header_13; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_2_header_14; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_2_header_15; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_parse_current_state; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_2_parse_current_offset; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_2_parse_transition_field; // @[ipsa.scala 103:24]
  reg [1:0] amplifier_1_2_next_processor_id; // @[ipsa.scala 103:24]
  reg  amplifier_1_2_next_config_id; // @[ipsa.scala 103:24]
  reg  amplifier_1_2_is_valid_processor; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_0; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_1; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_2; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_3; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_4; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_5; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_6; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_7; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_8; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_9; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_10; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_11; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_12; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_13; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_14; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_15; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_16; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_17; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_18; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_19; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_20; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_21; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_22; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_23; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_24; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_25; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_26; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_27; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_28; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_29; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_30; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_31; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_32; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_33; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_34; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_35; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_36; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_37; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_38; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_39; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_40; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_41; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_42; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_43; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_44; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_45; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_46; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_47; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_48; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_49; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_50; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_51; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_52; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_53; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_54; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_55; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_56; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_57; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_58; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_59; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_60; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_61; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_62; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_63; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_64; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_65; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_66; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_67; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_68; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_69; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_70; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_71; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_72; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_73; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_74; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_75; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_76; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_77; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_78; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_79; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_80; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_81; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_82; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_83; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_84; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_85; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_86; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_87; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_88; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_89; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_90; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_91; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_92; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_93; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_94; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_95; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_96; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_97; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_98; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_99; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_100; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_101; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_102; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_103; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_104; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_105; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_106; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_107; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_108; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_109; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_110; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_111; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_112; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_113; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_114; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_115; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_116; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_117; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_118; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_119; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_120; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_121; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_122; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_123; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_124; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_125; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_126; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_127; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_128; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_129; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_130; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_131; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_132; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_133; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_134; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_135; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_136; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_137; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_138; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_139; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_140; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_141; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_142; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_143; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_144; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_145; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_146; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_147; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_148; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_149; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_150; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_151; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_152; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_153; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_154; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_155; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_156; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_157; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_158; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_159; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_160; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_161; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_162; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_163; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_164; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_165; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_166; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_167; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_168; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_169; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_170; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_171; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_172; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_173; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_174; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_175; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_176; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_177; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_178; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_179; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_180; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_181; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_182; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_183; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_184; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_185; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_186; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_187; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_188; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_189; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_190; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_191; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_192; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_193; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_194; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_195; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_196; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_197; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_198; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_199; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_200; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_201; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_202; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_203; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_204; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_205; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_206; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_207; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_208; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_209; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_210; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_211; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_212; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_213; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_214; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_215; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_216; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_217; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_218; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_219; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_220; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_221; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_222; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_223; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_224; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_225; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_226; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_227; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_228; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_229; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_230; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_231; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_232; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_233; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_234; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_235; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_236; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_237; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_238; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_239; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_240; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_241; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_242; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_243; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_244; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_245; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_246; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_247; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_248; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_249; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_250; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_251; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_252; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_253; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_254; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_data_255; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_3_header_0; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_3_header_1; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_3_header_2; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_3_header_3; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_3_header_4; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_3_header_5; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_3_header_6; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_3_header_7; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_3_header_8; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_3_header_9; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_3_header_10; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_3_header_11; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_3_header_12; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_3_header_13; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_3_header_14; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_3_header_15; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_parse_current_state; // @[ipsa.scala 103:24]
  reg [7:0] amplifier_1_3_parse_current_offset; // @[ipsa.scala 103:24]
  reg [15:0] amplifier_1_3_parse_transition_field; // @[ipsa.scala 103:24]
  reg [1:0] amplifier_1_3_next_processor_id; // @[ipsa.scala 103:24]
  reg  amplifier_1_3_next_config_id; // @[ipsa.scala 103:24]
  reg  amplifier_1_3_is_valid_processor; // @[ipsa.scala 103:24]
  reg [1:0] next_proc_id_buf_0_0; // @[ipsa.scala 104:31]
  reg [1:0] next_proc_id_buf_0_1; // @[ipsa.scala 104:31]
  reg [1:0] next_proc_id_buf_0_2; // @[ipsa.scala 104:31]
  reg [1:0] next_proc_id_buf_0_3; // @[ipsa.scala 104:31]
  reg [1:0] next_proc_id_buf_1_0; // @[ipsa.scala 104:31]
  reg [1:0] next_proc_id_buf_1_1; // @[ipsa.scala 104:31]
  reg [1:0] next_proc_id_buf_1_2; // @[ipsa.scala 104:31]
  reg [1:0] next_proc_id_buf_1_3; // @[ipsa.scala 104:31]
  wire  _amplifier_0_0_T = trans_1_io_next_proc_id_out == 2'h0; // @[ipsa.scala 110:42]
  wire  _amplifier_0_1_T = trans_0_io_next_proc_id_out == 2'h1; // @[ipsa.scala 117:42]
  wire  _amplifier_0_2_T = trans_3_io_next_proc_id_out == 2'h2; // @[ipsa.scala 110:42]
  wire  _amplifier_0_3_T = trans_2_io_next_proc_id_out == 2'h3; // @[ipsa.scala 117:42]
  wire  _amplifier_1_0_T = next_proc_id_buf_0_2 == 2'h0; // @[ipsa.scala 136:36]
  wire  _amplifier_1_2_T = next_proc_id_buf_0_0 == 2'h2; // @[ipsa.scala 142:36]
  wire  _amplifier_1_1_T = next_proc_id_buf_0_3 == 2'h1; // @[ipsa.scala 136:36]
  wire  _amplifier_1_3_T = next_proc_id_buf_0_1 == 2'h3; // @[ipsa.scala 142:36]
  wire  _recv_0_T = next_proc_id_buf_1_3 == 2'h0; // @[ipsa.scala 153:36]
  wire  _recv_3_T = next_proc_id_buf_1_0 == 2'h3; // @[ipsa.scala 156:36]
  wire  _recv_1_T = next_proc_id_buf_1_2 == 2'h1; // @[ipsa.scala 153:36]
  wire  _recv_2_T = next_proc_id_buf_1_1 == 2'h2; // @[ipsa.scala 156:36]
  Processor proc_0 ( // @[ipsa.scala 62:25]
    .clock(proc_0_clock),
    .io_pipe_phv_in_data_0(proc_0_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_0_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_0_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_0_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_0_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_0_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_0_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_0_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_0_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_0_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_0_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_0_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_0_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_0_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_0_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_0_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_0_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_0_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_0_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_0_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_0_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_0_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_0_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_0_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_0_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_0_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_0_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_0_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_0_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_0_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_0_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_0_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_0_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_0_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_0_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_0_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_0_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_0_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_0_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_0_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_0_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_0_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_0_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_0_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_0_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_0_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_0_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_0_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_0_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_0_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_0_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_0_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_0_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_0_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_0_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_0_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_0_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_0_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_0_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_0_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_0_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_0_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_0_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_0_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_0_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_0_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_0_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_0_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_0_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_0_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_0_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_0_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_0_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_0_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_0_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_0_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_0_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_0_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_0_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_0_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_0_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_0_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_0_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_0_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_0_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_0_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_0_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_0_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_0_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_0_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_0_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_0_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_0_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_0_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_0_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_0_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_0_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_0_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_0_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_0_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_0_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_0_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_0_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_0_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_0_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_0_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_0_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_0_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_0_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_0_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_0_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_0_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_0_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_0_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_0_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_0_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_0_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_0_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_0_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_0_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_0_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_0_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_0_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_0_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_0_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_0_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_0_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_0_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_0_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_0_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_0_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_0_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_0_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_0_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_0_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_0_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_0_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_0_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_0_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_0_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_0_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_0_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_0_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_0_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_0_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_0_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_0_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_0_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_0_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_0_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_0_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_0_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_0_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_0_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_0_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_0_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_0_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_0_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_0_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_0_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(proc_0_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(proc_0_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(proc_0_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(proc_0_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(proc_0_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(proc_0_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(proc_0_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(proc_0_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(proc_0_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(proc_0_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(proc_0_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(proc_0_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(proc_0_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(proc_0_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(proc_0_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(proc_0_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(proc_0_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(proc_0_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(proc_0_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(proc_0_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(proc_0_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(proc_0_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(proc_0_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(proc_0_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(proc_0_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(proc_0_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(proc_0_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(proc_0_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(proc_0_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(proc_0_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(proc_0_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(proc_0_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(proc_0_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(proc_0_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(proc_0_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(proc_0_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(proc_0_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(proc_0_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(proc_0_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(proc_0_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(proc_0_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(proc_0_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(proc_0_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(proc_0_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(proc_0_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(proc_0_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(proc_0_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(proc_0_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(proc_0_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(proc_0_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(proc_0_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(proc_0_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(proc_0_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(proc_0_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(proc_0_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(proc_0_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(proc_0_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(proc_0_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(proc_0_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(proc_0_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(proc_0_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(proc_0_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(proc_0_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(proc_0_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(proc_0_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(proc_0_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(proc_0_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(proc_0_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(proc_0_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(proc_0_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(proc_0_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(proc_0_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(proc_0_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(proc_0_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(proc_0_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(proc_0_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(proc_0_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(proc_0_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(proc_0_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(proc_0_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(proc_0_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(proc_0_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(proc_0_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(proc_0_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(proc_0_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(proc_0_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(proc_0_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(proc_0_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(proc_0_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(proc_0_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(proc_0_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(proc_0_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(proc_0_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(proc_0_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(proc_0_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(proc_0_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(proc_0_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_0_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_0_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_0_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_0_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_0_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_0_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_0_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_0_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_0_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_0_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_0_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_0_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_0_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_0_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_0_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_0_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_0_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_0_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_0_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_0_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_0_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_0_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_0_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_0_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_0_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_0_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_0_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_0_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_0_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_0_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_0_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_0_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_0_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_0_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_0_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_0_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_0_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_0_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_0_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_0_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_0_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_0_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_0_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_0_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_0_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_0_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_0_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_0_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_0_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_0_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_0_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_0_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_0_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_0_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_0_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_0_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_0_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_0_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_0_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_0_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_0_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_0_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_0_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_0_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_0_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_0_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_0_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_0_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_0_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_0_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_0_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_0_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_0_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_0_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_0_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_0_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_0_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_0_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_0_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_0_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_0_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_0_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_0_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_0_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_0_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_0_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_0_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_0_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_0_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_0_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_0_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_0_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_0_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_0_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_0_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_0_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_0_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_0_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_0_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_0_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_0_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_0_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_0_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_0_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_0_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_0_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_0_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_0_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_0_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_0_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_0_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_0_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_0_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_0_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_0_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_0_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_0_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_0_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_0_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_0_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_0_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_0_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_0_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_0_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_0_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_0_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_0_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_0_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_0_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_0_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_0_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_0_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_0_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_0_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_0_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_0_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_0_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_0_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_0_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_0_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_0_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_0_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_0_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_0_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_0_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_0_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_0_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_0_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_0_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_0_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_0_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_0_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_0_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_0_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_0_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_0_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_0_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_0_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_0_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_0_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_0_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_0_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_0_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_0_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_0_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_0_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_0_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_0_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_0_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_0_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_0_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_0_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_0_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_0_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_0_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_0_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_0_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_0_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_0_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_0_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_0_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(proc_0_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(proc_0_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(proc_0_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(proc_0_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(proc_0_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(proc_0_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(proc_0_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(proc_0_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(proc_0_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(proc_0_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(proc_0_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(proc_0_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(proc_0_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(proc_0_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(proc_0_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(proc_0_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(proc_0_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(proc_0_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(proc_0_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(proc_0_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(proc_0_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(proc_0_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(proc_0_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(proc_0_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(proc_0_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(proc_0_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(proc_0_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(proc_0_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(proc_0_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(proc_0_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(proc_0_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(proc_0_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(proc_0_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(proc_0_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(proc_0_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(proc_0_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(proc_0_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(proc_0_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(proc_0_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(proc_0_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(proc_0_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(proc_0_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(proc_0_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(proc_0_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(proc_0_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(proc_0_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(proc_0_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(proc_0_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(proc_0_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(proc_0_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(proc_0_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(proc_0_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(proc_0_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(proc_0_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(proc_0_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(proc_0_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(proc_0_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(proc_0_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(proc_0_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(proc_0_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(proc_0_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(proc_0_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(proc_0_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(proc_0_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(proc_0_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(proc_0_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(proc_0_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(proc_0_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(proc_0_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(proc_0_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(proc_0_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(proc_0_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(proc_0_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(proc_0_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(proc_0_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(proc_0_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(proc_0_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(proc_0_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(proc_0_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(proc_0_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(proc_0_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(proc_0_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(proc_0_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(proc_0_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(proc_0_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(proc_0_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(proc_0_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(proc_0_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(proc_0_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(proc_0_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(proc_0_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(proc_0_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(proc_0_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(proc_0_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(proc_0_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(proc_0_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(proc_0_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_0_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_0_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_0_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_0_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_0_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_0_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_0_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_0_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_0_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_0_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_0_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_0_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_0_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_0_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_0_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_0_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_0_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_0_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_0_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_0_io_pipe_phv_out_next_config_id),
    .io_mod_par_mod_en(proc_0_io_mod_par_mod_en),
    .io_mod_par_mod_last_mau_id_mod(proc_0_io_mod_par_mod_last_mau_id_mod),
    .io_mod_par_mod_last_mau_id(proc_0_io_mod_par_mod_last_mau_id),
    .io_mod_par_mod_cs(proc_0_io_mod_par_mod_cs),
    .io_mod_par_mod_module_mod_state_id_mod(proc_0_io_mod_par_mod_module_mod_state_id_mod),
    .io_mod_par_mod_module_mod_state_id(proc_0_io_mod_par_mod_module_mod_state_id),
    .io_mod_par_mod_module_mod_sram_w_cs(proc_0_io_mod_par_mod_module_mod_sram_w_cs),
    .io_mod_par_mod_module_mod_sram_w_en(proc_0_io_mod_par_mod_module_mod_sram_w_en),
    .io_mod_par_mod_module_mod_sram_w_addr(proc_0_io_mod_par_mod_module_mod_sram_w_addr),
    .io_mod_par_mod_module_mod_sram_w_data(proc_0_io_mod_par_mod_module_mod_sram_w_data),
    .io_mod_mat_mod_en(proc_0_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_0_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_header_id(proc_0_io_mod_mat_mod_key_mod_header_id),
    .io_mod_mat_mod_key_mod_internal_offset(proc_0_io_mod_mat_mod_key_mod_internal_offset),
    .io_mod_mat_mod_key_mod_key_length(proc_0_io_mod_mat_mod_key_mod_key_length),
    .io_mod_mat_mod_table_mod_sram_id_table_0(proc_0_io_mod_mat_mod_table_mod_sram_id_table_0),
    .io_mod_mat_mod_table_mod_sram_id_table_1(proc_0_io_mod_mat_mod_table_mod_sram_id_table_1),
    .io_mod_mat_mod_table_mod_sram_id_table_2(proc_0_io_mod_mat_mod_table_mod_sram_id_table_2),
    .io_mod_mat_mod_table_mod_sram_id_table_3(proc_0_io_mod_mat_mod_table_mod_sram_id_table_3),
    .io_mod_mat_mod_table_mod_sram_id_table_4(proc_0_io_mod_mat_mod_table_mod_sram_id_table_4),
    .io_mod_mat_mod_table_mod_sram_id_table_5(proc_0_io_mod_mat_mod_table_mod_sram_id_table_5),
    .io_mod_mat_mod_table_mod_sram_id_table_6(proc_0_io_mod_mat_mod_table_mod_sram_id_table_6),
    .io_mod_mat_mod_table_mod_sram_id_table_7(proc_0_io_mod_mat_mod_table_mod_sram_id_table_7),
    .io_mod_mat_mod_table_mod_sram_id_table_8(proc_0_io_mod_mat_mod_table_mod_sram_id_table_8),
    .io_mod_mat_mod_table_mod_sram_id_table_9(proc_0_io_mod_mat_mod_table_mod_sram_id_table_9),
    .io_mod_mat_mod_table_mod_sram_id_table_10(proc_0_io_mod_mat_mod_table_mod_sram_id_table_10),
    .io_mod_mat_mod_table_mod_sram_id_table_11(proc_0_io_mod_mat_mod_table_mod_sram_id_table_11),
    .io_mod_mat_mod_table_mod_sram_id_table_12(proc_0_io_mod_mat_mod_table_mod_sram_id_table_12),
    .io_mod_mat_mod_table_mod_sram_id_table_13(proc_0_io_mod_mat_mod_table_mod_sram_id_table_13),
    .io_mod_mat_mod_table_mod_sram_id_table_14(proc_0_io_mod_mat_mod_table_mod_sram_id_table_14),
    .io_mod_mat_mod_table_mod_sram_id_table_15(proc_0_io_mod_mat_mod_table_mod_sram_id_table_15),
    .io_mod_mat_mod_table_mod_sram_id_table_16(proc_0_io_mod_mat_mod_table_mod_sram_id_table_16),
    .io_mod_mat_mod_table_mod_sram_id_table_17(proc_0_io_mod_mat_mod_table_mod_sram_id_table_17),
    .io_mod_mat_mod_table_mod_sram_id_table_18(proc_0_io_mod_mat_mod_table_mod_sram_id_table_18),
    .io_mod_mat_mod_table_mod_sram_id_table_19(proc_0_io_mod_mat_mod_table_mod_sram_id_table_19),
    .io_mod_mat_mod_table_mod_sram_id_table_20(proc_0_io_mod_mat_mod_table_mod_sram_id_table_20),
    .io_mod_mat_mod_table_mod_sram_id_table_21(proc_0_io_mod_mat_mod_table_mod_sram_id_table_21),
    .io_mod_mat_mod_table_mod_sram_id_table_22(proc_0_io_mod_mat_mod_table_mod_sram_id_table_22),
    .io_mod_mat_mod_table_mod_sram_id_table_23(proc_0_io_mod_mat_mod_table_mod_sram_id_table_23),
    .io_mod_mat_mod_table_mod_sram_id_table_24(proc_0_io_mod_mat_mod_table_mod_sram_id_table_24),
    .io_mod_mat_mod_table_mod_sram_id_table_25(proc_0_io_mod_mat_mod_table_mod_sram_id_table_25),
    .io_mod_mat_mod_table_mod_sram_id_table_26(proc_0_io_mod_mat_mod_table_mod_sram_id_table_26),
    .io_mod_mat_mod_table_mod_sram_id_table_27(proc_0_io_mod_mat_mod_table_mod_sram_id_table_27),
    .io_mod_mat_mod_table_mod_sram_id_table_28(proc_0_io_mod_mat_mod_table_mod_sram_id_table_28),
    .io_mod_mat_mod_table_mod_sram_id_table_29(proc_0_io_mod_mat_mod_table_mod_sram_id_table_29),
    .io_mod_mat_mod_table_mod_sram_id_table_30(proc_0_io_mod_mat_mod_table_mod_sram_id_table_30),
    .io_mod_mat_mod_table_mod_sram_id_table_31(proc_0_io_mod_mat_mod_table_mod_sram_id_table_31),
    .io_mod_mat_mod_table_mod_sram_id_table_32(proc_0_io_mod_mat_mod_table_mod_sram_id_table_32),
    .io_mod_mat_mod_table_mod_sram_id_table_33(proc_0_io_mod_mat_mod_table_mod_sram_id_table_33),
    .io_mod_mat_mod_table_mod_sram_id_table_34(proc_0_io_mod_mat_mod_table_mod_sram_id_table_34),
    .io_mod_mat_mod_table_mod_sram_id_table_35(proc_0_io_mod_mat_mod_table_mod_sram_id_table_35),
    .io_mod_mat_mod_table_mod_sram_id_table_36(proc_0_io_mod_mat_mod_table_mod_sram_id_table_36),
    .io_mod_mat_mod_table_mod_sram_id_table_37(proc_0_io_mod_mat_mod_table_mod_sram_id_table_37),
    .io_mod_mat_mod_table_mod_sram_id_table_38(proc_0_io_mod_mat_mod_table_mod_sram_id_table_38),
    .io_mod_mat_mod_table_mod_sram_id_table_39(proc_0_io_mod_mat_mod_table_mod_sram_id_table_39),
    .io_mod_mat_mod_table_mod_sram_id_table_40(proc_0_io_mod_mat_mod_table_mod_sram_id_table_40),
    .io_mod_mat_mod_table_mod_sram_id_table_41(proc_0_io_mod_mat_mod_table_mod_sram_id_table_41),
    .io_mod_mat_mod_table_mod_sram_id_table_42(proc_0_io_mod_mat_mod_table_mod_sram_id_table_42),
    .io_mod_mat_mod_table_mod_sram_id_table_43(proc_0_io_mod_mat_mod_table_mod_sram_id_table_43),
    .io_mod_mat_mod_table_mod_sram_id_table_44(proc_0_io_mod_mat_mod_table_mod_sram_id_table_44),
    .io_mod_mat_mod_table_mod_sram_id_table_45(proc_0_io_mod_mat_mod_table_mod_sram_id_table_45),
    .io_mod_mat_mod_table_mod_sram_id_table_46(proc_0_io_mod_mat_mod_table_mod_sram_id_table_46),
    .io_mod_mat_mod_table_mod_sram_id_table_47(proc_0_io_mod_mat_mod_table_mod_sram_id_table_47),
    .io_mod_mat_mod_table_mod_sram_id_table_48(proc_0_io_mod_mat_mod_table_mod_sram_id_table_48),
    .io_mod_mat_mod_table_mod_sram_id_table_49(proc_0_io_mod_mat_mod_table_mod_sram_id_table_49),
    .io_mod_mat_mod_table_mod_sram_id_table_50(proc_0_io_mod_mat_mod_table_mod_sram_id_table_50),
    .io_mod_mat_mod_table_mod_sram_id_table_51(proc_0_io_mod_mat_mod_table_mod_sram_id_table_51),
    .io_mod_mat_mod_table_mod_sram_id_table_52(proc_0_io_mod_mat_mod_table_mod_sram_id_table_52),
    .io_mod_mat_mod_table_mod_sram_id_table_53(proc_0_io_mod_mat_mod_table_mod_sram_id_table_53),
    .io_mod_mat_mod_table_mod_sram_id_table_54(proc_0_io_mod_mat_mod_table_mod_sram_id_table_54),
    .io_mod_mat_mod_table_mod_sram_id_table_55(proc_0_io_mod_mat_mod_table_mod_sram_id_table_55),
    .io_mod_mat_mod_table_mod_sram_id_table_56(proc_0_io_mod_mat_mod_table_mod_sram_id_table_56),
    .io_mod_mat_mod_table_mod_sram_id_table_57(proc_0_io_mod_mat_mod_table_mod_sram_id_table_57),
    .io_mod_mat_mod_table_mod_sram_id_table_58(proc_0_io_mod_mat_mod_table_mod_sram_id_table_58),
    .io_mod_mat_mod_table_mod_sram_id_table_59(proc_0_io_mod_mat_mod_table_mod_sram_id_table_59),
    .io_mod_mat_mod_table_mod_sram_id_table_60(proc_0_io_mod_mat_mod_table_mod_sram_id_table_60),
    .io_mod_mat_mod_table_mod_sram_id_table_61(proc_0_io_mod_mat_mod_table_mod_sram_id_table_61),
    .io_mod_mat_mod_table_mod_sram_id_table_62(proc_0_io_mod_mat_mod_table_mod_sram_id_table_62),
    .io_mod_mat_mod_table_mod_sram_id_table_63(proc_0_io_mod_mat_mod_table_mod_sram_id_table_63),
    .io_mod_mat_mod_table_mod_table_width(proc_0_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_table_mod_table_depth(proc_0_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_act_mod_en_0(proc_0_io_mod_act_mod_en_0),
    .io_mod_act_mod_en_1(proc_0_io_mod_act_mod_en_1),
    .io_mod_act_mod_addr(proc_0_io_mod_act_mod_addr),
    .io_mod_act_mod_data_0(proc_0_io_mod_act_mod_data_0),
    .io_mod_act_mod_data_1(proc_0_io_mod_act_mod_data_1),
    .io_mem_cluster_0_en(proc_0_io_mem_cluster_0_en),
    .io_mem_cluster_0_addr(proc_0_io_mem_cluster_0_addr),
    .io_mem_cluster_0_data(proc_0_io_mem_cluster_0_data),
    .io_mem_cluster_1_en(proc_0_io_mem_cluster_1_en),
    .io_mem_cluster_1_addr(proc_0_io_mem_cluster_1_addr),
    .io_mem_cluster_1_data(proc_0_io_mem_cluster_1_data),
    .io_mem_cluster_2_en(proc_0_io_mem_cluster_2_en),
    .io_mem_cluster_2_addr(proc_0_io_mem_cluster_2_addr),
    .io_mem_cluster_2_data(proc_0_io_mem_cluster_2_data),
    .io_mem_cluster_3_en(proc_0_io_mem_cluster_3_en),
    .io_mem_cluster_3_addr(proc_0_io_mem_cluster_3_addr),
    .io_mem_cluster_3_data(proc_0_io_mem_cluster_3_data),
    .io_mem_cluster_4_en(proc_0_io_mem_cluster_4_en),
    .io_mem_cluster_4_addr(proc_0_io_mem_cluster_4_addr),
    .io_mem_cluster_4_data(proc_0_io_mem_cluster_4_data),
    .io_mem_cluster_5_en(proc_0_io_mem_cluster_5_en),
    .io_mem_cluster_5_addr(proc_0_io_mem_cluster_5_addr),
    .io_mem_cluster_5_data(proc_0_io_mem_cluster_5_data),
    .io_mem_cluster_6_en(proc_0_io_mem_cluster_6_en),
    .io_mem_cluster_6_addr(proc_0_io_mem_cluster_6_addr),
    .io_mem_cluster_6_data(proc_0_io_mem_cluster_6_data),
    .io_mem_cluster_7_en(proc_0_io_mem_cluster_7_en),
    .io_mem_cluster_7_addr(proc_0_io_mem_cluster_7_addr),
    .io_mem_cluster_7_data(proc_0_io_mem_cluster_7_data),
    .io_mem_cluster_8_en(proc_0_io_mem_cluster_8_en),
    .io_mem_cluster_8_addr(proc_0_io_mem_cluster_8_addr),
    .io_mem_cluster_8_data(proc_0_io_mem_cluster_8_data),
    .io_mem_cluster_9_en(proc_0_io_mem_cluster_9_en),
    .io_mem_cluster_9_addr(proc_0_io_mem_cluster_9_addr),
    .io_mem_cluster_9_data(proc_0_io_mem_cluster_9_data),
    .io_mem_cluster_10_en(proc_0_io_mem_cluster_10_en),
    .io_mem_cluster_10_addr(proc_0_io_mem_cluster_10_addr),
    .io_mem_cluster_10_data(proc_0_io_mem_cluster_10_data),
    .io_mem_cluster_11_en(proc_0_io_mem_cluster_11_en),
    .io_mem_cluster_11_addr(proc_0_io_mem_cluster_11_addr),
    .io_mem_cluster_11_data(proc_0_io_mem_cluster_11_data),
    .io_mem_cluster_12_en(proc_0_io_mem_cluster_12_en),
    .io_mem_cluster_12_addr(proc_0_io_mem_cluster_12_addr),
    .io_mem_cluster_12_data(proc_0_io_mem_cluster_12_data),
    .io_mem_cluster_13_en(proc_0_io_mem_cluster_13_en),
    .io_mem_cluster_13_addr(proc_0_io_mem_cluster_13_addr),
    .io_mem_cluster_13_data(proc_0_io_mem_cluster_13_data),
    .io_mem_cluster_14_en(proc_0_io_mem_cluster_14_en),
    .io_mem_cluster_14_addr(proc_0_io_mem_cluster_14_addr),
    .io_mem_cluster_14_data(proc_0_io_mem_cluster_14_data),
    .io_mem_cluster_15_en(proc_0_io_mem_cluster_15_en),
    .io_mem_cluster_15_addr(proc_0_io_mem_cluster_15_addr),
    .io_mem_cluster_15_data(proc_0_io_mem_cluster_15_data),
    .io_mem_cluster_16_en(proc_0_io_mem_cluster_16_en),
    .io_mem_cluster_16_addr(proc_0_io_mem_cluster_16_addr),
    .io_mem_cluster_16_data(proc_0_io_mem_cluster_16_data),
    .io_mem_cluster_17_en(proc_0_io_mem_cluster_17_en),
    .io_mem_cluster_17_addr(proc_0_io_mem_cluster_17_addr),
    .io_mem_cluster_17_data(proc_0_io_mem_cluster_17_data),
    .io_mem_cluster_18_en(proc_0_io_mem_cluster_18_en),
    .io_mem_cluster_18_addr(proc_0_io_mem_cluster_18_addr),
    .io_mem_cluster_18_data(proc_0_io_mem_cluster_18_data),
    .io_mem_cluster_19_en(proc_0_io_mem_cluster_19_en),
    .io_mem_cluster_19_addr(proc_0_io_mem_cluster_19_addr),
    .io_mem_cluster_19_data(proc_0_io_mem_cluster_19_data),
    .io_mem_cluster_20_en(proc_0_io_mem_cluster_20_en),
    .io_mem_cluster_20_addr(proc_0_io_mem_cluster_20_addr),
    .io_mem_cluster_20_data(proc_0_io_mem_cluster_20_data),
    .io_mem_cluster_21_en(proc_0_io_mem_cluster_21_en),
    .io_mem_cluster_21_addr(proc_0_io_mem_cluster_21_addr),
    .io_mem_cluster_21_data(proc_0_io_mem_cluster_21_data),
    .io_mem_cluster_22_en(proc_0_io_mem_cluster_22_en),
    .io_mem_cluster_22_addr(proc_0_io_mem_cluster_22_addr),
    .io_mem_cluster_22_data(proc_0_io_mem_cluster_22_data),
    .io_mem_cluster_23_en(proc_0_io_mem_cluster_23_en),
    .io_mem_cluster_23_addr(proc_0_io_mem_cluster_23_addr),
    .io_mem_cluster_23_data(proc_0_io_mem_cluster_23_data),
    .io_mem_cluster_24_en(proc_0_io_mem_cluster_24_en),
    .io_mem_cluster_24_addr(proc_0_io_mem_cluster_24_addr),
    .io_mem_cluster_24_data(proc_0_io_mem_cluster_24_data),
    .io_mem_cluster_25_en(proc_0_io_mem_cluster_25_en),
    .io_mem_cluster_25_addr(proc_0_io_mem_cluster_25_addr),
    .io_mem_cluster_25_data(proc_0_io_mem_cluster_25_data),
    .io_mem_cluster_26_en(proc_0_io_mem_cluster_26_en),
    .io_mem_cluster_26_addr(proc_0_io_mem_cluster_26_addr),
    .io_mem_cluster_26_data(proc_0_io_mem_cluster_26_data),
    .io_mem_cluster_27_en(proc_0_io_mem_cluster_27_en),
    .io_mem_cluster_27_addr(proc_0_io_mem_cluster_27_addr),
    .io_mem_cluster_27_data(proc_0_io_mem_cluster_27_data),
    .io_mem_cluster_28_en(proc_0_io_mem_cluster_28_en),
    .io_mem_cluster_28_addr(proc_0_io_mem_cluster_28_addr),
    .io_mem_cluster_28_data(proc_0_io_mem_cluster_28_data),
    .io_mem_cluster_29_en(proc_0_io_mem_cluster_29_en),
    .io_mem_cluster_29_addr(proc_0_io_mem_cluster_29_addr),
    .io_mem_cluster_29_data(proc_0_io_mem_cluster_29_data),
    .io_mem_cluster_30_en(proc_0_io_mem_cluster_30_en),
    .io_mem_cluster_30_addr(proc_0_io_mem_cluster_30_addr),
    .io_mem_cluster_30_data(proc_0_io_mem_cluster_30_data),
    .io_mem_cluster_31_en(proc_0_io_mem_cluster_31_en),
    .io_mem_cluster_31_addr(proc_0_io_mem_cluster_31_addr),
    .io_mem_cluster_31_data(proc_0_io_mem_cluster_31_data),
    .io_mem_cluster_32_en(proc_0_io_mem_cluster_32_en),
    .io_mem_cluster_32_addr(proc_0_io_mem_cluster_32_addr),
    .io_mem_cluster_32_data(proc_0_io_mem_cluster_32_data),
    .io_mem_cluster_33_en(proc_0_io_mem_cluster_33_en),
    .io_mem_cluster_33_addr(proc_0_io_mem_cluster_33_addr),
    .io_mem_cluster_33_data(proc_0_io_mem_cluster_33_data),
    .io_mem_cluster_34_en(proc_0_io_mem_cluster_34_en),
    .io_mem_cluster_34_addr(proc_0_io_mem_cluster_34_addr),
    .io_mem_cluster_34_data(proc_0_io_mem_cluster_34_data),
    .io_mem_cluster_35_en(proc_0_io_mem_cluster_35_en),
    .io_mem_cluster_35_addr(proc_0_io_mem_cluster_35_addr),
    .io_mem_cluster_35_data(proc_0_io_mem_cluster_35_data),
    .io_mem_cluster_36_en(proc_0_io_mem_cluster_36_en),
    .io_mem_cluster_36_addr(proc_0_io_mem_cluster_36_addr),
    .io_mem_cluster_36_data(proc_0_io_mem_cluster_36_data),
    .io_mem_cluster_37_en(proc_0_io_mem_cluster_37_en),
    .io_mem_cluster_37_addr(proc_0_io_mem_cluster_37_addr),
    .io_mem_cluster_37_data(proc_0_io_mem_cluster_37_data),
    .io_mem_cluster_38_en(proc_0_io_mem_cluster_38_en),
    .io_mem_cluster_38_addr(proc_0_io_mem_cluster_38_addr),
    .io_mem_cluster_38_data(proc_0_io_mem_cluster_38_data),
    .io_mem_cluster_39_en(proc_0_io_mem_cluster_39_en),
    .io_mem_cluster_39_addr(proc_0_io_mem_cluster_39_addr),
    .io_mem_cluster_39_data(proc_0_io_mem_cluster_39_data),
    .io_mem_cluster_40_en(proc_0_io_mem_cluster_40_en),
    .io_mem_cluster_40_addr(proc_0_io_mem_cluster_40_addr),
    .io_mem_cluster_40_data(proc_0_io_mem_cluster_40_data),
    .io_mem_cluster_41_en(proc_0_io_mem_cluster_41_en),
    .io_mem_cluster_41_addr(proc_0_io_mem_cluster_41_addr),
    .io_mem_cluster_41_data(proc_0_io_mem_cluster_41_data),
    .io_mem_cluster_42_en(proc_0_io_mem_cluster_42_en),
    .io_mem_cluster_42_addr(proc_0_io_mem_cluster_42_addr),
    .io_mem_cluster_42_data(proc_0_io_mem_cluster_42_data),
    .io_mem_cluster_43_en(proc_0_io_mem_cluster_43_en),
    .io_mem_cluster_43_addr(proc_0_io_mem_cluster_43_addr),
    .io_mem_cluster_43_data(proc_0_io_mem_cluster_43_data),
    .io_mem_cluster_44_en(proc_0_io_mem_cluster_44_en),
    .io_mem_cluster_44_addr(proc_0_io_mem_cluster_44_addr),
    .io_mem_cluster_44_data(proc_0_io_mem_cluster_44_data),
    .io_mem_cluster_45_en(proc_0_io_mem_cluster_45_en),
    .io_mem_cluster_45_addr(proc_0_io_mem_cluster_45_addr),
    .io_mem_cluster_45_data(proc_0_io_mem_cluster_45_data),
    .io_mem_cluster_46_en(proc_0_io_mem_cluster_46_en),
    .io_mem_cluster_46_addr(proc_0_io_mem_cluster_46_addr),
    .io_mem_cluster_46_data(proc_0_io_mem_cluster_46_data),
    .io_mem_cluster_47_en(proc_0_io_mem_cluster_47_en),
    .io_mem_cluster_47_addr(proc_0_io_mem_cluster_47_addr),
    .io_mem_cluster_47_data(proc_0_io_mem_cluster_47_data),
    .io_mem_cluster_48_en(proc_0_io_mem_cluster_48_en),
    .io_mem_cluster_48_addr(proc_0_io_mem_cluster_48_addr),
    .io_mem_cluster_48_data(proc_0_io_mem_cluster_48_data),
    .io_mem_cluster_49_en(proc_0_io_mem_cluster_49_en),
    .io_mem_cluster_49_addr(proc_0_io_mem_cluster_49_addr),
    .io_mem_cluster_49_data(proc_0_io_mem_cluster_49_data),
    .io_mem_cluster_50_en(proc_0_io_mem_cluster_50_en),
    .io_mem_cluster_50_addr(proc_0_io_mem_cluster_50_addr),
    .io_mem_cluster_50_data(proc_0_io_mem_cluster_50_data),
    .io_mem_cluster_51_en(proc_0_io_mem_cluster_51_en),
    .io_mem_cluster_51_addr(proc_0_io_mem_cluster_51_addr),
    .io_mem_cluster_51_data(proc_0_io_mem_cluster_51_data),
    .io_mem_cluster_52_en(proc_0_io_mem_cluster_52_en),
    .io_mem_cluster_52_addr(proc_0_io_mem_cluster_52_addr),
    .io_mem_cluster_52_data(proc_0_io_mem_cluster_52_data),
    .io_mem_cluster_53_en(proc_0_io_mem_cluster_53_en),
    .io_mem_cluster_53_addr(proc_0_io_mem_cluster_53_addr),
    .io_mem_cluster_53_data(proc_0_io_mem_cluster_53_data),
    .io_mem_cluster_54_en(proc_0_io_mem_cluster_54_en),
    .io_mem_cluster_54_addr(proc_0_io_mem_cluster_54_addr),
    .io_mem_cluster_54_data(proc_0_io_mem_cluster_54_data),
    .io_mem_cluster_55_en(proc_0_io_mem_cluster_55_en),
    .io_mem_cluster_55_addr(proc_0_io_mem_cluster_55_addr),
    .io_mem_cluster_55_data(proc_0_io_mem_cluster_55_data),
    .io_mem_cluster_56_en(proc_0_io_mem_cluster_56_en),
    .io_mem_cluster_56_addr(proc_0_io_mem_cluster_56_addr),
    .io_mem_cluster_56_data(proc_0_io_mem_cluster_56_data),
    .io_mem_cluster_57_en(proc_0_io_mem_cluster_57_en),
    .io_mem_cluster_57_addr(proc_0_io_mem_cluster_57_addr),
    .io_mem_cluster_57_data(proc_0_io_mem_cluster_57_data),
    .io_mem_cluster_58_en(proc_0_io_mem_cluster_58_en),
    .io_mem_cluster_58_addr(proc_0_io_mem_cluster_58_addr),
    .io_mem_cluster_58_data(proc_0_io_mem_cluster_58_data),
    .io_mem_cluster_59_en(proc_0_io_mem_cluster_59_en),
    .io_mem_cluster_59_addr(proc_0_io_mem_cluster_59_addr),
    .io_mem_cluster_59_data(proc_0_io_mem_cluster_59_data),
    .io_mem_cluster_60_en(proc_0_io_mem_cluster_60_en),
    .io_mem_cluster_60_addr(proc_0_io_mem_cluster_60_addr),
    .io_mem_cluster_60_data(proc_0_io_mem_cluster_60_data),
    .io_mem_cluster_61_en(proc_0_io_mem_cluster_61_en),
    .io_mem_cluster_61_addr(proc_0_io_mem_cluster_61_addr),
    .io_mem_cluster_61_data(proc_0_io_mem_cluster_61_data),
    .io_mem_cluster_62_en(proc_0_io_mem_cluster_62_en),
    .io_mem_cluster_62_addr(proc_0_io_mem_cluster_62_addr),
    .io_mem_cluster_62_data(proc_0_io_mem_cluster_62_data),
    .io_mem_cluster_63_en(proc_0_io_mem_cluster_63_en),
    .io_mem_cluster_63_addr(proc_0_io_mem_cluster_63_addr),
    .io_mem_cluster_63_data(proc_0_io_mem_cluster_63_data)
  );
  Processor proc_1 ( // @[ipsa.scala 62:25]
    .clock(proc_1_clock),
    .io_pipe_phv_in_data_0(proc_1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(proc_1_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(proc_1_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(proc_1_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(proc_1_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(proc_1_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(proc_1_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(proc_1_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(proc_1_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(proc_1_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(proc_1_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(proc_1_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(proc_1_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(proc_1_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(proc_1_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(proc_1_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(proc_1_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(proc_1_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(proc_1_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(proc_1_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(proc_1_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(proc_1_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(proc_1_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(proc_1_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(proc_1_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(proc_1_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(proc_1_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(proc_1_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(proc_1_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(proc_1_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(proc_1_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(proc_1_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(proc_1_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(proc_1_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(proc_1_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(proc_1_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(proc_1_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(proc_1_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(proc_1_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(proc_1_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(proc_1_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(proc_1_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(proc_1_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(proc_1_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(proc_1_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(proc_1_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(proc_1_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(proc_1_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(proc_1_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(proc_1_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(proc_1_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(proc_1_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(proc_1_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(proc_1_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(proc_1_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(proc_1_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(proc_1_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(proc_1_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(proc_1_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(proc_1_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(proc_1_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(proc_1_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(proc_1_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(proc_1_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(proc_1_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(proc_1_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(proc_1_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(proc_1_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(proc_1_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(proc_1_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(proc_1_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(proc_1_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(proc_1_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(proc_1_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(proc_1_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(proc_1_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(proc_1_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(proc_1_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(proc_1_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(proc_1_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(proc_1_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(proc_1_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(proc_1_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(proc_1_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(proc_1_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(proc_1_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(proc_1_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(proc_1_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(proc_1_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(proc_1_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(proc_1_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(proc_1_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(proc_1_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(proc_1_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(proc_1_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(proc_1_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(proc_1_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(proc_1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(proc_1_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(proc_1_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(proc_1_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(proc_1_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(proc_1_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(proc_1_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(proc_1_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(proc_1_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(proc_1_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(proc_1_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(proc_1_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(proc_1_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(proc_1_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(proc_1_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(proc_1_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(proc_1_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(proc_1_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(proc_1_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(proc_1_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(proc_1_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(proc_1_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(proc_1_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(proc_1_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(proc_1_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(proc_1_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(proc_1_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(proc_1_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(proc_1_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(proc_1_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(proc_1_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(proc_1_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(proc_1_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(proc_1_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(proc_1_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(proc_1_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(proc_1_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(proc_1_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(proc_1_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(proc_1_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(proc_1_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(proc_1_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(proc_1_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(proc_1_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(proc_1_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(proc_1_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(proc_1_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(proc_1_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(proc_1_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(proc_1_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(proc_1_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(proc_1_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(proc_1_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(proc_1_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(proc_1_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(proc_1_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(proc_1_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(proc_1_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(proc_1_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(proc_1_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(proc_1_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(proc_1_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(proc_1_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(proc_1_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(proc_1_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(proc_1_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(proc_1_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(proc_1_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(proc_1_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(proc_1_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(proc_1_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(proc_1_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(proc_1_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(proc_1_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(proc_1_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(proc_1_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(proc_1_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(proc_1_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(proc_1_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(proc_1_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(proc_1_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(proc_1_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(proc_1_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(proc_1_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(proc_1_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(proc_1_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(proc_1_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(proc_1_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(proc_1_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(proc_1_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(proc_1_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(proc_1_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(proc_1_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(proc_1_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(proc_1_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(proc_1_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(proc_1_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(proc_1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_1_io_pipe_phv_out_next_config_id),
    .io_mod_par_mod_en(proc_1_io_mod_par_mod_en),
    .io_mod_par_mod_last_mau_id_mod(proc_1_io_mod_par_mod_last_mau_id_mod),
    .io_mod_par_mod_last_mau_id(proc_1_io_mod_par_mod_last_mau_id),
    .io_mod_par_mod_cs(proc_1_io_mod_par_mod_cs),
    .io_mod_par_mod_module_mod_state_id_mod(proc_1_io_mod_par_mod_module_mod_state_id_mod),
    .io_mod_par_mod_module_mod_state_id(proc_1_io_mod_par_mod_module_mod_state_id),
    .io_mod_par_mod_module_mod_sram_w_cs(proc_1_io_mod_par_mod_module_mod_sram_w_cs),
    .io_mod_par_mod_module_mod_sram_w_en(proc_1_io_mod_par_mod_module_mod_sram_w_en),
    .io_mod_par_mod_module_mod_sram_w_addr(proc_1_io_mod_par_mod_module_mod_sram_w_addr),
    .io_mod_par_mod_module_mod_sram_w_data(proc_1_io_mod_par_mod_module_mod_sram_w_data),
    .io_mod_mat_mod_en(proc_1_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_1_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_header_id(proc_1_io_mod_mat_mod_key_mod_header_id),
    .io_mod_mat_mod_key_mod_internal_offset(proc_1_io_mod_mat_mod_key_mod_internal_offset),
    .io_mod_mat_mod_key_mod_key_length(proc_1_io_mod_mat_mod_key_mod_key_length),
    .io_mod_mat_mod_table_mod_sram_id_table_0(proc_1_io_mod_mat_mod_table_mod_sram_id_table_0),
    .io_mod_mat_mod_table_mod_sram_id_table_1(proc_1_io_mod_mat_mod_table_mod_sram_id_table_1),
    .io_mod_mat_mod_table_mod_sram_id_table_2(proc_1_io_mod_mat_mod_table_mod_sram_id_table_2),
    .io_mod_mat_mod_table_mod_sram_id_table_3(proc_1_io_mod_mat_mod_table_mod_sram_id_table_3),
    .io_mod_mat_mod_table_mod_sram_id_table_4(proc_1_io_mod_mat_mod_table_mod_sram_id_table_4),
    .io_mod_mat_mod_table_mod_sram_id_table_5(proc_1_io_mod_mat_mod_table_mod_sram_id_table_5),
    .io_mod_mat_mod_table_mod_sram_id_table_6(proc_1_io_mod_mat_mod_table_mod_sram_id_table_6),
    .io_mod_mat_mod_table_mod_sram_id_table_7(proc_1_io_mod_mat_mod_table_mod_sram_id_table_7),
    .io_mod_mat_mod_table_mod_sram_id_table_8(proc_1_io_mod_mat_mod_table_mod_sram_id_table_8),
    .io_mod_mat_mod_table_mod_sram_id_table_9(proc_1_io_mod_mat_mod_table_mod_sram_id_table_9),
    .io_mod_mat_mod_table_mod_sram_id_table_10(proc_1_io_mod_mat_mod_table_mod_sram_id_table_10),
    .io_mod_mat_mod_table_mod_sram_id_table_11(proc_1_io_mod_mat_mod_table_mod_sram_id_table_11),
    .io_mod_mat_mod_table_mod_sram_id_table_12(proc_1_io_mod_mat_mod_table_mod_sram_id_table_12),
    .io_mod_mat_mod_table_mod_sram_id_table_13(proc_1_io_mod_mat_mod_table_mod_sram_id_table_13),
    .io_mod_mat_mod_table_mod_sram_id_table_14(proc_1_io_mod_mat_mod_table_mod_sram_id_table_14),
    .io_mod_mat_mod_table_mod_sram_id_table_15(proc_1_io_mod_mat_mod_table_mod_sram_id_table_15),
    .io_mod_mat_mod_table_mod_sram_id_table_16(proc_1_io_mod_mat_mod_table_mod_sram_id_table_16),
    .io_mod_mat_mod_table_mod_sram_id_table_17(proc_1_io_mod_mat_mod_table_mod_sram_id_table_17),
    .io_mod_mat_mod_table_mod_sram_id_table_18(proc_1_io_mod_mat_mod_table_mod_sram_id_table_18),
    .io_mod_mat_mod_table_mod_sram_id_table_19(proc_1_io_mod_mat_mod_table_mod_sram_id_table_19),
    .io_mod_mat_mod_table_mod_sram_id_table_20(proc_1_io_mod_mat_mod_table_mod_sram_id_table_20),
    .io_mod_mat_mod_table_mod_sram_id_table_21(proc_1_io_mod_mat_mod_table_mod_sram_id_table_21),
    .io_mod_mat_mod_table_mod_sram_id_table_22(proc_1_io_mod_mat_mod_table_mod_sram_id_table_22),
    .io_mod_mat_mod_table_mod_sram_id_table_23(proc_1_io_mod_mat_mod_table_mod_sram_id_table_23),
    .io_mod_mat_mod_table_mod_sram_id_table_24(proc_1_io_mod_mat_mod_table_mod_sram_id_table_24),
    .io_mod_mat_mod_table_mod_sram_id_table_25(proc_1_io_mod_mat_mod_table_mod_sram_id_table_25),
    .io_mod_mat_mod_table_mod_sram_id_table_26(proc_1_io_mod_mat_mod_table_mod_sram_id_table_26),
    .io_mod_mat_mod_table_mod_sram_id_table_27(proc_1_io_mod_mat_mod_table_mod_sram_id_table_27),
    .io_mod_mat_mod_table_mod_sram_id_table_28(proc_1_io_mod_mat_mod_table_mod_sram_id_table_28),
    .io_mod_mat_mod_table_mod_sram_id_table_29(proc_1_io_mod_mat_mod_table_mod_sram_id_table_29),
    .io_mod_mat_mod_table_mod_sram_id_table_30(proc_1_io_mod_mat_mod_table_mod_sram_id_table_30),
    .io_mod_mat_mod_table_mod_sram_id_table_31(proc_1_io_mod_mat_mod_table_mod_sram_id_table_31),
    .io_mod_mat_mod_table_mod_sram_id_table_32(proc_1_io_mod_mat_mod_table_mod_sram_id_table_32),
    .io_mod_mat_mod_table_mod_sram_id_table_33(proc_1_io_mod_mat_mod_table_mod_sram_id_table_33),
    .io_mod_mat_mod_table_mod_sram_id_table_34(proc_1_io_mod_mat_mod_table_mod_sram_id_table_34),
    .io_mod_mat_mod_table_mod_sram_id_table_35(proc_1_io_mod_mat_mod_table_mod_sram_id_table_35),
    .io_mod_mat_mod_table_mod_sram_id_table_36(proc_1_io_mod_mat_mod_table_mod_sram_id_table_36),
    .io_mod_mat_mod_table_mod_sram_id_table_37(proc_1_io_mod_mat_mod_table_mod_sram_id_table_37),
    .io_mod_mat_mod_table_mod_sram_id_table_38(proc_1_io_mod_mat_mod_table_mod_sram_id_table_38),
    .io_mod_mat_mod_table_mod_sram_id_table_39(proc_1_io_mod_mat_mod_table_mod_sram_id_table_39),
    .io_mod_mat_mod_table_mod_sram_id_table_40(proc_1_io_mod_mat_mod_table_mod_sram_id_table_40),
    .io_mod_mat_mod_table_mod_sram_id_table_41(proc_1_io_mod_mat_mod_table_mod_sram_id_table_41),
    .io_mod_mat_mod_table_mod_sram_id_table_42(proc_1_io_mod_mat_mod_table_mod_sram_id_table_42),
    .io_mod_mat_mod_table_mod_sram_id_table_43(proc_1_io_mod_mat_mod_table_mod_sram_id_table_43),
    .io_mod_mat_mod_table_mod_sram_id_table_44(proc_1_io_mod_mat_mod_table_mod_sram_id_table_44),
    .io_mod_mat_mod_table_mod_sram_id_table_45(proc_1_io_mod_mat_mod_table_mod_sram_id_table_45),
    .io_mod_mat_mod_table_mod_sram_id_table_46(proc_1_io_mod_mat_mod_table_mod_sram_id_table_46),
    .io_mod_mat_mod_table_mod_sram_id_table_47(proc_1_io_mod_mat_mod_table_mod_sram_id_table_47),
    .io_mod_mat_mod_table_mod_sram_id_table_48(proc_1_io_mod_mat_mod_table_mod_sram_id_table_48),
    .io_mod_mat_mod_table_mod_sram_id_table_49(proc_1_io_mod_mat_mod_table_mod_sram_id_table_49),
    .io_mod_mat_mod_table_mod_sram_id_table_50(proc_1_io_mod_mat_mod_table_mod_sram_id_table_50),
    .io_mod_mat_mod_table_mod_sram_id_table_51(proc_1_io_mod_mat_mod_table_mod_sram_id_table_51),
    .io_mod_mat_mod_table_mod_sram_id_table_52(proc_1_io_mod_mat_mod_table_mod_sram_id_table_52),
    .io_mod_mat_mod_table_mod_sram_id_table_53(proc_1_io_mod_mat_mod_table_mod_sram_id_table_53),
    .io_mod_mat_mod_table_mod_sram_id_table_54(proc_1_io_mod_mat_mod_table_mod_sram_id_table_54),
    .io_mod_mat_mod_table_mod_sram_id_table_55(proc_1_io_mod_mat_mod_table_mod_sram_id_table_55),
    .io_mod_mat_mod_table_mod_sram_id_table_56(proc_1_io_mod_mat_mod_table_mod_sram_id_table_56),
    .io_mod_mat_mod_table_mod_sram_id_table_57(proc_1_io_mod_mat_mod_table_mod_sram_id_table_57),
    .io_mod_mat_mod_table_mod_sram_id_table_58(proc_1_io_mod_mat_mod_table_mod_sram_id_table_58),
    .io_mod_mat_mod_table_mod_sram_id_table_59(proc_1_io_mod_mat_mod_table_mod_sram_id_table_59),
    .io_mod_mat_mod_table_mod_sram_id_table_60(proc_1_io_mod_mat_mod_table_mod_sram_id_table_60),
    .io_mod_mat_mod_table_mod_sram_id_table_61(proc_1_io_mod_mat_mod_table_mod_sram_id_table_61),
    .io_mod_mat_mod_table_mod_sram_id_table_62(proc_1_io_mod_mat_mod_table_mod_sram_id_table_62),
    .io_mod_mat_mod_table_mod_sram_id_table_63(proc_1_io_mod_mat_mod_table_mod_sram_id_table_63),
    .io_mod_mat_mod_table_mod_table_width(proc_1_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_table_mod_table_depth(proc_1_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_act_mod_en_0(proc_1_io_mod_act_mod_en_0),
    .io_mod_act_mod_en_1(proc_1_io_mod_act_mod_en_1),
    .io_mod_act_mod_addr(proc_1_io_mod_act_mod_addr),
    .io_mod_act_mod_data_0(proc_1_io_mod_act_mod_data_0),
    .io_mod_act_mod_data_1(proc_1_io_mod_act_mod_data_1),
    .io_mem_cluster_0_en(proc_1_io_mem_cluster_0_en),
    .io_mem_cluster_0_addr(proc_1_io_mem_cluster_0_addr),
    .io_mem_cluster_0_data(proc_1_io_mem_cluster_0_data),
    .io_mem_cluster_1_en(proc_1_io_mem_cluster_1_en),
    .io_mem_cluster_1_addr(proc_1_io_mem_cluster_1_addr),
    .io_mem_cluster_1_data(proc_1_io_mem_cluster_1_data),
    .io_mem_cluster_2_en(proc_1_io_mem_cluster_2_en),
    .io_mem_cluster_2_addr(proc_1_io_mem_cluster_2_addr),
    .io_mem_cluster_2_data(proc_1_io_mem_cluster_2_data),
    .io_mem_cluster_3_en(proc_1_io_mem_cluster_3_en),
    .io_mem_cluster_3_addr(proc_1_io_mem_cluster_3_addr),
    .io_mem_cluster_3_data(proc_1_io_mem_cluster_3_data),
    .io_mem_cluster_4_en(proc_1_io_mem_cluster_4_en),
    .io_mem_cluster_4_addr(proc_1_io_mem_cluster_4_addr),
    .io_mem_cluster_4_data(proc_1_io_mem_cluster_4_data),
    .io_mem_cluster_5_en(proc_1_io_mem_cluster_5_en),
    .io_mem_cluster_5_addr(proc_1_io_mem_cluster_5_addr),
    .io_mem_cluster_5_data(proc_1_io_mem_cluster_5_data),
    .io_mem_cluster_6_en(proc_1_io_mem_cluster_6_en),
    .io_mem_cluster_6_addr(proc_1_io_mem_cluster_6_addr),
    .io_mem_cluster_6_data(proc_1_io_mem_cluster_6_data),
    .io_mem_cluster_7_en(proc_1_io_mem_cluster_7_en),
    .io_mem_cluster_7_addr(proc_1_io_mem_cluster_7_addr),
    .io_mem_cluster_7_data(proc_1_io_mem_cluster_7_data),
    .io_mem_cluster_8_en(proc_1_io_mem_cluster_8_en),
    .io_mem_cluster_8_addr(proc_1_io_mem_cluster_8_addr),
    .io_mem_cluster_8_data(proc_1_io_mem_cluster_8_data),
    .io_mem_cluster_9_en(proc_1_io_mem_cluster_9_en),
    .io_mem_cluster_9_addr(proc_1_io_mem_cluster_9_addr),
    .io_mem_cluster_9_data(proc_1_io_mem_cluster_9_data),
    .io_mem_cluster_10_en(proc_1_io_mem_cluster_10_en),
    .io_mem_cluster_10_addr(proc_1_io_mem_cluster_10_addr),
    .io_mem_cluster_10_data(proc_1_io_mem_cluster_10_data),
    .io_mem_cluster_11_en(proc_1_io_mem_cluster_11_en),
    .io_mem_cluster_11_addr(proc_1_io_mem_cluster_11_addr),
    .io_mem_cluster_11_data(proc_1_io_mem_cluster_11_data),
    .io_mem_cluster_12_en(proc_1_io_mem_cluster_12_en),
    .io_mem_cluster_12_addr(proc_1_io_mem_cluster_12_addr),
    .io_mem_cluster_12_data(proc_1_io_mem_cluster_12_data),
    .io_mem_cluster_13_en(proc_1_io_mem_cluster_13_en),
    .io_mem_cluster_13_addr(proc_1_io_mem_cluster_13_addr),
    .io_mem_cluster_13_data(proc_1_io_mem_cluster_13_data),
    .io_mem_cluster_14_en(proc_1_io_mem_cluster_14_en),
    .io_mem_cluster_14_addr(proc_1_io_mem_cluster_14_addr),
    .io_mem_cluster_14_data(proc_1_io_mem_cluster_14_data),
    .io_mem_cluster_15_en(proc_1_io_mem_cluster_15_en),
    .io_mem_cluster_15_addr(proc_1_io_mem_cluster_15_addr),
    .io_mem_cluster_15_data(proc_1_io_mem_cluster_15_data),
    .io_mem_cluster_16_en(proc_1_io_mem_cluster_16_en),
    .io_mem_cluster_16_addr(proc_1_io_mem_cluster_16_addr),
    .io_mem_cluster_16_data(proc_1_io_mem_cluster_16_data),
    .io_mem_cluster_17_en(proc_1_io_mem_cluster_17_en),
    .io_mem_cluster_17_addr(proc_1_io_mem_cluster_17_addr),
    .io_mem_cluster_17_data(proc_1_io_mem_cluster_17_data),
    .io_mem_cluster_18_en(proc_1_io_mem_cluster_18_en),
    .io_mem_cluster_18_addr(proc_1_io_mem_cluster_18_addr),
    .io_mem_cluster_18_data(proc_1_io_mem_cluster_18_data),
    .io_mem_cluster_19_en(proc_1_io_mem_cluster_19_en),
    .io_mem_cluster_19_addr(proc_1_io_mem_cluster_19_addr),
    .io_mem_cluster_19_data(proc_1_io_mem_cluster_19_data),
    .io_mem_cluster_20_en(proc_1_io_mem_cluster_20_en),
    .io_mem_cluster_20_addr(proc_1_io_mem_cluster_20_addr),
    .io_mem_cluster_20_data(proc_1_io_mem_cluster_20_data),
    .io_mem_cluster_21_en(proc_1_io_mem_cluster_21_en),
    .io_mem_cluster_21_addr(proc_1_io_mem_cluster_21_addr),
    .io_mem_cluster_21_data(proc_1_io_mem_cluster_21_data),
    .io_mem_cluster_22_en(proc_1_io_mem_cluster_22_en),
    .io_mem_cluster_22_addr(proc_1_io_mem_cluster_22_addr),
    .io_mem_cluster_22_data(proc_1_io_mem_cluster_22_data),
    .io_mem_cluster_23_en(proc_1_io_mem_cluster_23_en),
    .io_mem_cluster_23_addr(proc_1_io_mem_cluster_23_addr),
    .io_mem_cluster_23_data(proc_1_io_mem_cluster_23_data),
    .io_mem_cluster_24_en(proc_1_io_mem_cluster_24_en),
    .io_mem_cluster_24_addr(proc_1_io_mem_cluster_24_addr),
    .io_mem_cluster_24_data(proc_1_io_mem_cluster_24_data),
    .io_mem_cluster_25_en(proc_1_io_mem_cluster_25_en),
    .io_mem_cluster_25_addr(proc_1_io_mem_cluster_25_addr),
    .io_mem_cluster_25_data(proc_1_io_mem_cluster_25_data),
    .io_mem_cluster_26_en(proc_1_io_mem_cluster_26_en),
    .io_mem_cluster_26_addr(proc_1_io_mem_cluster_26_addr),
    .io_mem_cluster_26_data(proc_1_io_mem_cluster_26_data),
    .io_mem_cluster_27_en(proc_1_io_mem_cluster_27_en),
    .io_mem_cluster_27_addr(proc_1_io_mem_cluster_27_addr),
    .io_mem_cluster_27_data(proc_1_io_mem_cluster_27_data),
    .io_mem_cluster_28_en(proc_1_io_mem_cluster_28_en),
    .io_mem_cluster_28_addr(proc_1_io_mem_cluster_28_addr),
    .io_mem_cluster_28_data(proc_1_io_mem_cluster_28_data),
    .io_mem_cluster_29_en(proc_1_io_mem_cluster_29_en),
    .io_mem_cluster_29_addr(proc_1_io_mem_cluster_29_addr),
    .io_mem_cluster_29_data(proc_1_io_mem_cluster_29_data),
    .io_mem_cluster_30_en(proc_1_io_mem_cluster_30_en),
    .io_mem_cluster_30_addr(proc_1_io_mem_cluster_30_addr),
    .io_mem_cluster_30_data(proc_1_io_mem_cluster_30_data),
    .io_mem_cluster_31_en(proc_1_io_mem_cluster_31_en),
    .io_mem_cluster_31_addr(proc_1_io_mem_cluster_31_addr),
    .io_mem_cluster_31_data(proc_1_io_mem_cluster_31_data),
    .io_mem_cluster_32_en(proc_1_io_mem_cluster_32_en),
    .io_mem_cluster_32_addr(proc_1_io_mem_cluster_32_addr),
    .io_mem_cluster_32_data(proc_1_io_mem_cluster_32_data),
    .io_mem_cluster_33_en(proc_1_io_mem_cluster_33_en),
    .io_mem_cluster_33_addr(proc_1_io_mem_cluster_33_addr),
    .io_mem_cluster_33_data(proc_1_io_mem_cluster_33_data),
    .io_mem_cluster_34_en(proc_1_io_mem_cluster_34_en),
    .io_mem_cluster_34_addr(proc_1_io_mem_cluster_34_addr),
    .io_mem_cluster_34_data(proc_1_io_mem_cluster_34_data),
    .io_mem_cluster_35_en(proc_1_io_mem_cluster_35_en),
    .io_mem_cluster_35_addr(proc_1_io_mem_cluster_35_addr),
    .io_mem_cluster_35_data(proc_1_io_mem_cluster_35_data),
    .io_mem_cluster_36_en(proc_1_io_mem_cluster_36_en),
    .io_mem_cluster_36_addr(proc_1_io_mem_cluster_36_addr),
    .io_mem_cluster_36_data(proc_1_io_mem_cluster_36_data),
    .io_mem_cluster_37_en(proc_1_io_mem_cluster_37_en),
    .io_mem_cluster_37_addr(proc_1_io_mem_cluster_37_addr),
    .io_mem_cluster_37_data(proc_1_io_mem_cluster_37_data),
    .io_mem_cluster_38_en(proc_1_io_mem_cluster_38_en),
    .io_mem_cluster_38_addr(proc_1_io_mem_cluster_38_addr),
    .io_mem_cluster_38_data(proc_1_io_mem_cluster_38_data),
    .io_mem_cluster_39_en(proc_1_io_mem_cluster_39_en),
    .io_mem_cluster_39_addr(proc_1_io_mem_cluster_39_addr),
    .io_mem_cluster_39_data(proc_1_io_mem_cluster_39_data),
    .io_mem_cluster_40_en(proc_1_io_mem_cluster_40_en),
    .io_mem_cluster_40_addr(proc_1_io_mem_cluster_40_addr),
    .io_mem_cluster_40_data(proc_1_io_mem_cluster_40_data),
    .io_mem_cluster_41_en(proc_1_io_mem_cluster_41_en),
    .io_mem_cluster_41_addr(proc_1_io_mem_cluster_41_addr),
    .io_mem_cluster_41_data(proc_1_io_mem_cluster_41_data),
    .io_mem_cluster_42_en(proc_1_io_mem_cluster_42_en),
    .io_mem_cluster_42_addr(proc_1_io_mem_cluster_42_addr),
    .io_mem_cluster_42_data(proc_1_io_mem_cluster_42_data),
    .io_mem_cluster_43_en(proc_1_io_mem_cluster_43_en),
    .io_mem_cluster_43_addr(proc_1_io_mem_cluster_43_addr),
    .io_mem_cluster_43_data(proc_1_io_mem_cluster_43_data),
    .io_mem_cluster_44_en(proc_1_io_mem_cluster_44_en),
    .io_mem_cluster_44_addr(proc_1_io_mem_cluster_44_addr),
    .io_mem_cluster_44_data(proc_1_io_mem_cluster_44_data),
    .io_mem_cluster_45_en(proc_1_io_mem_cluster_45_en),
    .io_mem_cluster_45_addr(proc_1_io_mem_cluster_45_addr),
    .io_mem_cluster_45_data(proc_1_io_mem_cluster_45_data),
    .io_mem_cluster_46_en(proc_1_io_mem_cluster_46_en),
    .io_mem_cluster_46_addr(proc_1_io_mem_cluster_46_addr),
    .io_mem_cluster_46_data(proc_1_io_mem_cluster_46_data),
    .io_mem_cluster_47_en(proc_1_io_mem_cluster_47_en),
    .io_mem_cluster_47_addr(proc_1_io_mem_cluster_47_addr),
    .io_mem_cluster_47_data(proc_1_io_mem_cluster_47_data),
    .io_mem_cluster_48_en(proc_1_io_mem_cluster_48_en),
    .io_mem_cluster_48_addr(proc_1_io_mem_cluster_48_addr),
    .io_mem_cluster_48_data(proc_1_io_mem_cluster_48_data),
    .io_mem_cluster_49_en(proc_1_io_mem_cluster_49_en),
    .io_mem_cluster_49_addr(proc_1_io_mem_cluster_49_addr),
    .io_mem_cluster_49_data(proc_1_io_mem_cluster_49_data),
    .io_mem_cluster_50_en(proc_1_io_mem_cluster_50_en),
    .io_mem_cluster_50_addr(proc_1_io_mem_cluster_50_addr),
    .io_mem_cluster_50_data(proc_1_io_mem_cluster_50_data),
    .io_mem_cluster_51_en(proc_1_io_mem_cluster_51_en),
    .io_mem_cluster_51_addr(proc_1_io_mem_cluster_51_addr),
    .io_mem_cluster_51_data(proc_1_io_mem_cluster_51_data),
    .io_mem_cluster_52_en(proc_1_io_mem_cluster_52_en),
    .io_mem_cluster_52_addr(proc_1_io_mem_cluster_52_addr),
    .io_mem_cluster_52_data(proc_1_io_mem_cluster_52_data),
    .io_mem_cluster_53_en(proc_1_io_mem_cluster_53_en),
    .io_mem_cluster_53_addr(proc_1_io_mem_cluster_53_addr),
    .io_mem_cluster_53_data(proc_1_io_mem_cluster_53_data),
    .io_mem_cluster_54_en(proc_1_io_mem_cluster_54_en),
    .io_mem_cluster_54_addr(proc_1_io_mem_cluster_54_addr),
    .io_mem_cluster_54_data(proc_1_io_mem_cluster_54_data),
    .io_mem_cluster_55_en(proc_1_io_mem_cluster_55_en),
    .io_mem_cluster_55_addr(proc_1_io_mem_cluster_55_addr),
    .io_mem_cluster_55_data(proc_1_io_mem_cluster_55_data),
    .io_mem_cluster_56_en(proc_1_io_mem_cluster_56_en),
    .io_mem_cluster_56_addr(proc_1_io_mem_cluster_56_addr),
    .io_mem_cluster_56_data(proc_1_io_mem_cluster_56_data),
    .io_mem_cluster_57_en(proc_1_io_mem_cluster_57_en),
    .io_mem_cluster_57_addr(proc_1_io_mem_cluster_57_addr),
    .io_mem_cluster_57_data(proc_1_io_mem_cluster_57_data),
    .io_mem_cluster_58_en(proc_1_io_mem_cluster_58_en),
    .io_mem_cluster_58_addr(proc_1_io_mem_cluster_58_addr),
    .io_mem_cluster_58_data(proc_1_io_mem_cluster_58_data),
    .io_mem_cluster_59_en(proc_1_io_mem_cluster_59_en),
    .io_mem_cluster_59_addr(proc_1_io_mem_cluster_59_addr),
    .io_mem_cluster_59_data(proc_1_io_mem_cluster_59_data),
    .io_mem_cluster_60_en(proc_1_io_mem_cluster_60_en),
    .io_mem_cluster_60_addr(proc_1_io_mem_cluster_60_addr),
    .io_mem_cluster_60_data(proc_1_io_mem_cluster_60_data),
    .io_mem_cluster_61_en(proc_1_io_mem_cluster_61_en),
    .io_mem_cluster_61_addr(proc_1_io_mem_cluster_61_addr),
    .io_mem_cluster_61_data(proc_1_io_mem_cluster_61_data),
    .io_mem_cluster_62_en(proc_1_io_mem_cluster_62_en),
    .io_mem_cluster_62_addr(proc_1_io_mem_cluster_62_addr),
    .io_mem_cluster_62_data(proc_1_io_mem_cluster_62_data),
    .io_mem_cluster_63_en(proc_1_io_mem_cluster_63_en),
    .io_mem_cluster_63_addr(proc_1_io_mem_cluster_63_addr),
    .io_mem_cluster_63_data(proc_1_io_mem_cluster_63_data)
  );
  Processor proc_2 ( // @[ipsa.scala 62:25]
    .clock(proc_2_clock),
    .io_pipe_phv_in_data_0(proc_2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(proc_2_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(proc_2_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(proc_2_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(proc_2_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(proc_2_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(proc_2_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(proc_2_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(proc_2_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(proc_2_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(proc_2_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(proc_2_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(proc_2_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(proc_2_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(proc_2_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(proc_2_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(proc_2_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(proc_2_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(proc_2_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(proc_2_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(proc_2_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(proc_2_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(proc_2_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(proc_2_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(proc_2_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(proc_2_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(proc_2_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(proc_2_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(proc_2_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(proc_2_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(proc_2_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(proc_2_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(proc_2_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(proc_2_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(proc_2_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(proc_2_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(proc_2_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(proc_2_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(proc_2_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(proc_2_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(proc_2_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(proc_2_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(proc_2_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(proc_2_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(proc_2_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(proc_2_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(proc_2_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(proc_2_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(proc_2_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(proc_2_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(proc_2_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(proc_2_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(proc_2_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(proc_2_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(proc_2_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(proc_2_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(proc_2_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(proc_2_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(proc_2_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(proc_2_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(proc_2_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(proc_2_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(proc_2_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(proc_2_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(proc_2_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(proc_2_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(proc_2_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(proc_2_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(proc_2_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(proc_2_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(proc_2_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(proc_2_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(proc_2_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(proc_2_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(proc_2_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(proc_2_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(proc_2_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(proc_2_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(proc_2_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(proc_2_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(proc_2_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(proc_2_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(proc_2_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(proc_2_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(proc_2_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(proc_2_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(proc_2_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(proc_2_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(proc_2_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(proc_2_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(proc_2_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(proc_2_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(proc_2_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(proc_2_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(proc_2_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(proc_2_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(proc_2_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(proc_2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(proc_2_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(proc_2_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(proc_2_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(proc_2_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(proc_2_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(proc_2_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(proc_2_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(proc_2_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(proc_2_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(proc_2_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(proc_2_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(proc_2_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(proc_2_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(proc_2_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(proc_2_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(proc_2_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(proc_2_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(proc_2_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(proc_2_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(proc_2_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(proc_2_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(proc_2_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(proc_2_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(proc_2_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(proc_2_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(proc_2_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(proc_2_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(proc_2_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(proc_2_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(proc_2_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(proc_2_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(proc_2_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(proc_2_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(proc_2_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(proc_2_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(proc_2_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(proc_2_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(proc_2_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(proc_2_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(proc_2_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(proc_2_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(proc_2_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(proc_2_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(proc_2_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(proc_2_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(proc_2_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(proc_2_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(proc_2_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(proc_2_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(proc_2_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(proc_2_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(proc_2_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(proc_2_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(proc_2_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(proc_2_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(proc_2_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(proc_2_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(proc_2_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(proc_2_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(proc_2_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(proc_2_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(proc_2_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(proc_2_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(proc_2_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(proc_2_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(proc_2_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(proc_2_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(proc_2_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(proc_2_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(proc_2_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(proc_2_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(proc_2_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(proc_2_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(proc_2_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(proc_2_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(proc_2_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(proc_2_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(proc_2_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(proc_2_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(proc_2_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(proc_2_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(proc_2_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(proc_2_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(proc_2_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(proc_2_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(proc_2_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(proc_2_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(proc_2_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(proc_2_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(proc_2_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(proc_2_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(proc_2_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(proc_2_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(proc_2_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(proc_2_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(proc_2_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(proc_2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_2_io_pipe_phv_out_next_config_id),
    .io_mod_par_mod_en(proc_2_io_mod_par_mod_en),
    .io_mod_par_mod_last_mau_id_mod(proc_2_io_mod_par_mod_last_mau_id_mod),
    .io_mod_par_mod_last_mau_id(proc_2_io_mod_par_mod_last_mau_id),
    .io_mod_par_mod_cs(proc_2_io_mod_par_mod_cs),
    .io_mod_par_mod_module_mod_state_id_mod(proc_2_io_mod_par_mod_module_mod_state_id_mod),
    .io_mod_par_mod_module_mod_state_id(proc_2_io_mod_par_mod_module_mod_state_id),
    .io_mod_par_mod_module_mod_sram_w_cs(proc_2_io_mod_par_mod_module_mod_sram_w_cs),
    .io_mod_par_mod_module_mod_sram_w_en(proc_2_io_mod_par_mod_module_mod_sram_w_en),
    .io_mod_par_mod_module_mod_sram_w_addr(proc_2_io_mod_par_mod_module_mod_sram_w_addr),
    .io_mod_par_mod_module_mod_sram_w_data(proc_2_io_mod_par_mod_module_mod_sram_w_data),
    .io_mod_mat_mod_en(proc_2_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_2_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_header_id(proc_2_io_mod_mat_mod_key_mod_header_id),
    .io_mod_mat_mod_key_mod_internal_offset(proc_2_io_mod_mat_mod_key_mod_internal_offset),
    .io_mod_mat_mod_key_mod_key_length(proc_2_io_mod_mat_mod_key_mod_key_length),
    .io_mod_mat_mod_table_mod_sram_id_table_0(proc_2_io_mod_mat_mod_table_mod_sram_id_table_0),
    .io_mod_mat_mod_table_mod_sram_id_table_1(proc_2_io_mod_mat_mod_table_mod_sram_id_table_1),
    .io_mod_mat_mod_table_mod_sram_id_table_2(proc_2_io_mod_mat_mod_table_mod_sram_id_table_2),
    .io_mod_mat_mod_table_mod_sram_id_table_3(proc_2_io_mod_mat_mod_table_mod_sram_id_table_3),
    .io_mod_mat_mod_table_mod_sram_id_table_4(proc_2_io_mod_mat_mod_table_mod_sram_id_table_4),
    .io_mod_mat_mod_table_mod_sram_id_table_5(proc_2_io_mod_mat_mod_table_mod_sram_id_table_5),
    .io_mod_mat_mod_table_mod_sram_id_table_6(proc_2_io_mod_mat_mod_table_mod_sram_id_table_6),
    .io_mod_mat_mod_table_mod_sram_id_table_7(proc_2_io_mod_mat_mod_table_mod_sram_id_table_7),
    .io_mod_mat_mod_table_mod_sram_id_table_8(proc_2_io_mod_mat_mod_table_mod_sram_id_table_8),
    .io_mod_mat_mod_table_mod_sram_id_table_9(proc_2_io_mod_mat_mod_table_mod_sram_id_table_9),
    .io_mod_mat_mod_table_mod_sram_id_table_10(proc_2_io_mod_mat_mod_table_mod_sram_id_table_10),
    .io_mod_mat_mod_table_mod_sram_id_table_11(proc_2_io_mod_mat_mod_table_mod_sram_id_table_11),
    .io_mod_mat_mod_table_mod_sram_id_table_12(proc_2_io_mod_mat_mod_table_mod_sram_id_table_12),
    .io_mod_mat_mod_table_mod_sram_id_table_13(proc_2_io_mod_mat_mod_table_mod_sram_id_table_13),
    .io_mod_mat_mod_table_mod_sram_id_table_14(proc_2_io_mod_mat_mod_table_mod_sram_id_table_14),
    .io_mod_mat_mod_table_mod_sram_id_table_15(proc_2_io_mod_mat_mod_table_mod_sram_id_table_15),
    .io_mod_mat_mod_table_mod_sram_id_table_16(proc_2_io_mod_mat_mod_table_mod_sram_id_table_16),
    .io_mod_mat_mod_table_mod_sram_id_table_17(proc_2_io_mod_mat_mod_table_mod_sram_id_table_17),
    .io_mod_mat_mod_table_mod_sram_id_table_18(proc_2_io_mod_mat_mod_table_mod_sram_id_table_18),
    .io_mod_mat_mod_table_mod_sram_id_table_19(proc_2_io_mod_mat_mod_table_mod_sram_id_table_19),
    .io_mod_mat_mod_table_mod_sram_id_table_20(proc_2_io_mod_mat_mod_table_mod_sram_id_table_20),
    .io_mod_mat_mod_table_mod_sram_id_table_21(proc_2_io_mod_mat_mod_table_mod_sram_id_table_21),
    .io_mod_mat_mod_table_mod_sram_id_table_22(proc_2_io_mod_mat_mod_table_mod_sram_id_table_22),
    .io_mod_mat_mod_table_mod_sram_id_table_23(proc_2_io_mod_mat_mod_table_mod_sram_id_table_23),
    .io_mod_mat_mod_table_mod_sram_id_table_24(proc_2_io_mod_mat_mod_table_mod_sram_id_table_24),
    .io_mod_mat_mod_table_mod_sram_id_table_25(proc_2_io_mod_mat_mod_table_mod_sram_id_table_25),
    .io_mod_mat_mod_table_mod_sram_id_table_26(proc_2_io_mod_mat_mod_table_mod_sram_id_table_26),
    .io_mod_mat_mod_table_mod_sram_id_table_27(proc_2_io_mod_mat_mod_table_mod_sram_id_table_27),
    .io_mod_mat_mod_table_mod_sram_id_table_28(proc_2_io_mod_mat_mod_table_mod_sram_id_table_28),
    .io_mod_mat_mod_table_mod_sram_id_table_29(proc_2_io_mod_mat_mod_table_mod_sram_id_table_29),
    .io_mod_mat_mod_table_mod_sram_id_table_30(proc_2_io_mod_mat_mod_table_mod_sram_id_table_30),
    .io_mod_mat_mod_table_mod_sram_id_table_31(proc_2_io_mod_mat_mod_table_mod_sram_id_table_31),
    .io_mod_mat_mod_table_mod_sram_id_table_32(proc_2_io_mod_mat_mod_table_mod_sram_id_table_32),
    .io_mod_mat_mod_table_mod_sram_id_table_33(proc_2_io_mod_mat_mod_table_mod_sram_id_table_33),
    .io_mod_mat_mod_table_mod_sram_id_table_34(proc_2_io_mod_mat_mod_table_mod_sram_id_table_34),
    .io_mod_mat_mod_table_mod_sram_id_table_35(proc_2_io_mod_mat_mod_table_mod_sram_id_table_35),
    .io_mod_mat_mod_table_mod_sram_id_table_36(proc_2_io_mod_mat_mod_table_mod_sram_id_table_36),
    .io_mod_mat_mod_table_mod_sram_id_table_37(proc_2_io_mod_mat_mod_table_mod_sram_id_table_37),
    .io_mod_mat_mod_table_mod_sram_id_table_38(proc_2_io_mod_mat_mod_table_mod_sram_id_table_38),
    .io_mod_mat_mod_table_mod_sram_id_table_39(proc_2_io_mod_mat_mod_table_mod_sram_id_table_39),
    .io_mod_mat_mod_table_mod_sram_id_table_40(proc_2_io_mod_mat_mod_table_mod_sram_id_table_40),
    .io_mod_mat_mod_table_mod_sram_id_table_41(proc_2_io_mod_mat_mod_table_mod_sram_id_table_41),
    .io_mod_mat_mod_table_mod_sram_id_table_42(proc_2_io_mod_mat_mod_table_mod_sram_id_table_42),
    .io_mod_mat_mod_table_mod_sram_id_table_43(proc_2_io_mod_mat_mod_table_mod_sram_id_table_43),
    .io_mod_mat_mod_table_mod_sram_id_table_44(proc_2_io_mod_mat_mod_table_mod_sram_id_table_44),
    .io_mod_mat_mod_table_mod_sram_id_table_45(proc_2_io_mod_mat_mod_table_mod_sram_id_table_45),
    .io_mod_mat_mod_table_mod_sram_id_table_46(proc_2_io_mod_mat_mod_table_mod_sram_id_table_46),
    .io_mod_mat_mod_table_mod_sram_id_table_47(proc_2_io_mod_mat_mod_table_mod_sram_id_table_47),
    .io_mod_mat_mod_table_mod_sram_id_table_48(proc_2_io_mod_mat_mod_table_mod_sram_id_table_48),
    .io_mod_mat_mod_table_mod_sram_id_table_49(proc_2_io_mod_mat_mod_table_mod_sram_id_table_49),
    .io_mod_mat_mod_table_mod_sram_id_table_50(proc_2_io_mod_mat_mod_table_mod_sram_id_table_50),
    .io_mod_mat_mod_table_mod_sram_id_table_51(proc_2_io_mod_mat_mod_table_mod_sram_id_table_51),
    .io_mod_mat_mod_table_mod_sram_id_table_52(proc_2_io_mod_mat_mod_table_mod_sram_id_table_52),
    .io_mod_mat_mod_table_mod_sram_id_table_53(proc_2_io_mod_mat_mod_table_mod_sram_id_table_53),
    .io_mod_mat_mod_table_mod_sram_id_table_54(proc_2_io_mod_mat_mod_table_mod_sram_id_table_54),
    .io_mod_mat_mod_table_mod_sram_id_table_55(proc_2_io_mod_mat_mod_table_mod_sram_id_table_55),
    .io_mod_mat_mod_table_mod_sram_id_table_56(proc_2_io_mod_mat_mod_table_mod_sram_id_table_56),
    .io_mod_mat_mod_table_mod_sram_id_table_57(proc_2_io_mod_mat_mod_table_mod_sram_id_table_57),
    .io_mod_mat_mod_table_mod_sram_id_table_58(proc_2_io_mod_mat_mod_table_mod_sram_id_table_58),
    .io_mod_mat_mod_table_mod_sram_id_table_59(proc_2_io_mod_mat_mod_table_mod_sram_id_table_59),
    .io_mod_mat_mod_table_mod_sram_id_table_60(proc_2_io_mod_mat_mod_table_mod_sram_id_table_60),
    .io_mod_mat_mod_table_mod_sram_id_table_61(proc_2_io_mod_mat_mod_table_mod_sram_id_table_61),
    .io_mod_mat_mod_table_mod_sram_id_table_62(proc_2_io_mod_mat_mod_table_mod_sram_id_table_62),
    .io_mod_mat_mod_table_mod_sram_id_table_63(proc_2_io_mod_mat_mod_table_mod_sram_id_table_63),
    .io_mod_mat_mod_table_mod_table_width(proc_2_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_table_mod_table_depth(proc_2_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_act_mod_en_0(proc_2_io_mod_act_mod_en_0),
    .io_mod_act_mod_en_1(proc_2_io_mod_act_mod_en_1),
    .io_mod_act_mod_addr(proc_2_io_mod_act_mod_addr),
    .io_mod_act_mod_data_0(proc_2_io_mod_act_mod_data_0),
    .io_mod_act_mod_data_1(proc_2_io_mod_act_mod_data_1),
    .io_mem_cluster_0_en(proc_2_io_mem_cluster_0_en),
    .io_mem_cluster_0_addr(proc_2_io_mem_cluster_0_addr),
    .io_mem_cluster_0_data(proc_2_io_mem_cluster_0_data),
    .io_mem_cluster_1_en(proc_2_io_mem_cluster_1_en),
    .io_mem_cluster_1_addr(proc_2_io_mem_cluster_1_addr),
    .io_mem_cluster_1_data(proc_2_io_mem_cluster_1_data),
    .io_mem_cluster_2_en(proc_2_io_mem_cluster_2_en),
    .io_mem_cluster_2_addr(proc_2_io_mem_cluster_2_addr),
    .io_mem_cluster_2_data(proc_2_io_mem_cluster_2_data),
    .io_mem_cluster_3_en(proc_2_io_mem_cluster_3_en),
    .io_mem_cluster_3_addr(proc_2_io_mem_cluster_3_addr),
    .io_mem_cluster_3_data(proc_2_io_mem_cluster_3_data),
    .io_mem_cluster_4_en(proc_2_io_mem_cluster_4_en),
    .io_mem_cluster_4_addr(proc_2_io_mem_cluster_4_addr),
    .io_mem_cluster_4_data(proc_2_io_mem_cluster_4_data),
    .io_mem_cluster_5_en(proc_2_io_mem_cluster_5_en),
    .io_mem_cluster_5_addr(proc_2_io_mem_cluster_5_addr),
    .io_mem_cluster_5_data(proc_2_io_mem_cluster_5_data),
    .io_mem_cluster_6_en(proc_2_io_mem_cluster_6_en),
    .io_mem_cluster_6_addr(proc_2_io_mem_cluster_6_addr),
    .io_mem_cluster_6_data(proc_2_io_mem_cluster_6_data),
    .io_mem_cluster_7_en(proc_2_io_mem_cluster_7_en),
    .io_mem_cluster_7_addr(proc_2_io_mem_cluster_7_addr),
    .io_mem_cluster_7_data(proc_2_io_mem_cluster_7_data),
    .io_mem_cluster_8_en(proc_2_io_mem_cluster_8_en),
    .io_mem_cluster_8_addr(proc_2_io_mem_cluster_8_addr),
    .io_mem_cluster_8_data(proc_2_io_mem_cluster_8_data),
    .io_mem_cluster_9_en(proc_2_io_mem_cluster_9_en),
    .io_mem_cluster_9_addr(proc_2_io_mem_cluster_9_addr),
    .io_mem_cluster_9_data(proc_2_io_mem_cluster_9_data),
    .io_mem_cluster_10_en(proc_2_io_mem_cluster_10_en),
    .io_mem_cluster_10_addr(proc_2_io_mem_cluster_10_addr),
    .io_mem_cluster_10_data(proc_2_io_mem_cluster_10_data),
    .io_mem_cluster_11_en(proc_2_io_mem_cluster_11_en),
    .io_mem_cluster_11_addr(proc_2_io_mem_cluster_11_addr),
    .io_mem_cluster_11_data(proc_2_io_mem_cluster_11_data),
    .io_mem_cluster_12_en(proc_2_io_mem_cluster_12_en),
    .io_mem_cluster_12_addr(proc_2_io_mem_cluster_12_addr),
    .io_mem_cluster_12_data(proc_2_io_mem_cluster_12_data),
    .io_mem_cluster_13_en(proc_2_io_mem_cluster_13_en),
    .io_mem_cluster_13_addr(proc_2_io_mem_cluster_13_addr),
    .io_mem_cluster_13_data(proc_2_io_mem_cluster_13_data),
    .io_mem_cluster_14_en(proc_2_io_mem_cluster_14_en),
    .io_mem_cluster_14_addr(proc_2_io_mem_cluster_14_addr),
    .io_mem_cluster_14_data(proc_2_io_mem_cluster_14_data),
    .io_mem_cluster_15_en(proc_2_io_mem_cluster_15_en),
    .io_mem_cluster_15_addr(proc_2_io_mem_cluster_15_addr),
    .io_mem_cluster_15_data(proc_2_io_mem_cluster_15_data),
    .io_mem_cluster_16_en(proc_2_io_mem_cluster_16_en),
    .io_mem_cluster_16_addr(proc_2_io_mem_cluster_16_addr),
    .io_mem_cluster_16_data(proc_2_io_mem_cluster_16_data),
    .io_mem_cluster_17_en(proc_2_io_mem_cluster_17_en),
    .io_mem_cluster_17_addr(proc_2_io_mem_cluster_17_addr),
    .io_mem_cluster_17_data(proc_2_io_mem_cluster_17_data),
    .io_mem_cluster_18_en(proc_2_io_mem_cluster_18_en),
    .io_mem_cluster_18_addr(proc_2_io_mem_cluster_18_addr),
    .io_mem_cluster_18_data(proc_2_io_mem_cluster_18_data),
    .io_mem_cluster_19_en(proc_2_io_mem_cluster_19_en),
    .io_mem_cluster_19_addr(proc_2_io_mem_cluster_19_addr),
    .io_mem_cluster_19_data(proc_2_io_mem_cluster_19_data),
    .io_mem_cluster_20_en(proc_2_io_mem_cluster_20_en),
    .io_mem_cluster_20_addr(proc_2_io_mem_cluster_20_addr),
    .io_mem_cluster_20_data(proc_2_io_mem_cluster_20_data),
    .io_mem_cluster_21_en(proc_2_io_mem_cluster_21_en),
    .io_mem_cluster_21_addr(proc_2_io_mem_cluster_21_addr),
    .io_mem_cluster_21_data(proc_2_io_mem_cluster_21_data),
    .io_mem_cluster_22_en(proc_2_io_mem_cluster_22_en),
    .io_mem_cluster_22_addr(proc_2_io_mem_cluster_22_addr),
    .io_mem_cluster_22_data(proc_2_io_mem_cluster_22_data),
    .io_mem_cluster_23_en(proc_2_io_mem_cluster_23_en),
    .io_mem_cluster_23_addr(proc_2_io_mem_cluster_23_addr),
    .io_mem_cluster_23_data(proc_2_io_mem_cluster_23_data),
    .io_mem_cluster_24_en(proc_2_io_mem_cluster_24_en),
    .io_mem_cluster_24_addr(proc_2_io_mem_cluster_24_addr),
    .io_mem_cluster_24_data(proc_2_io_mem_cluster_24_data),
    .io_mem_cluster_25_en(proc_2_io_mem_cluster_25_en),
    .io_mem_cluster_25_addr(proc_2_io_mem_cluster_25_addr),
    .io_mem_cluster_25_data(proc_2_io_mem_cluster_25_data),
    .io_mem_cluster_26_en(proc_2_io_mem_cluster_26_en),
    .io_mem_cluster_26_addr(proc_2_io_mem_cluster_26_addr),
    .io_mem_cluster_26_data(proc_2_io_mem_cluster_26_data),
    .io_mem_cluster_27_en(proc_2_io_mem_cluster_27_en),
    .io_mem_cluster_27_addr(proc_2_io_mem_cluster_27_addr),
    .io_mem_cluster_27_data(proc_2_io_mem_cluster_27_data),
    .io_mem_cluster_28_en(proc_2_io_mem_cluster_28_en),
    .io_mem_cluster_28_addr(proc_2_io_mem_cluster_28_addr),
    .io_mem_cluster_28_data(proc_2_io_mem_cluster_28_data),
    .io_mem_cluster_29_en(proc_2_io_mem_cluster_29_en),
    .io_mem_cluster_29_addr(proc_2_io_mem_cluster_29_addr),
    .io_mem_cluster_29_data(proc_2_io_mem_cluster_29_data),
    .io_mem_cluster_30_en(proc_2_io_mem_cluster_30_en),
    .io_mem_cluster_30_addr(proc_2_io_mem_cluster_30_addr),
    .io_mem_cluster_30_data(proc_2_io_mem_cluster_30_data),
    .io_mem_cluster_31_en(proc_2_io_mem_cluster_31_en),
    .io_mem_cluster_31_addr(proc_2_io_mem_cluster_31_addr),
    .io_mem_cluster_31_data(proc_2_io_mem_cluster_31_data),
    .io_mem_cluster_32_en(proc_2_io_mem_cluster_32_en),
    .io_mem_cluster_32_addr(proc_2_io_mem_cluster_32_addr),
    .io_mem_cluster_32_data(proc_2_io_mem_cluster_32_data),
    .io_mem_cluster_33_en(proc_2_io_mem_cluster_33_en),
    .io_mem_cluster_33_addr(proc_2_io_mem_cluster_33_addr),
    .io_mem_cluster_33_data(proc_2_io_mem_cluster_33_data),
    .io_mem_cluster_34_en(proc_2_io_mem_cluster_34_en),
    .io_mem_cluster_34_addr(proc_2_io_mem_cluster_34_addr),
    .io_mem_cluster_34_data(proc_2_io_mem_cluster_34_data),
    .io_mem_cluster_35_en(proc_2_io_mem_cluster_35_en),
    .io_mem_cluster_35_addr(proc_2_io_mem_cluster_35_addr),
    .io_mem_cluster_35_data(proc_2_io_mem_cluster_35_data),
    .io_mem_cluster_36_en(proc_2_io_mem_cluster_36_en),
    .io_mem_cluster_36_addr(proc_2_io_mem_cluster_36_addr),
    .io_mem_cluster_36_data(proc_2_io_mem_cluster_36_data),
    .io_mem_cluster_37_en(proc_2_io_mem_cluster_37_en),
    .io_mem_cluster_37_addr(proc_2_io_mem_cluster_37_addr),
    .io_mem_cluster_37_data(proc_2_io_mem_cluster_37_data),
    .io_mem_cluster_38_en(proc_2_io_mem_cluster_38_en),
    .io_mem_cluster_38_addr(proc_2_io_mem_cluster_38_addr),
    .io_mem_cluster_38_data(proc_2_io_mem_cluster_38_data),
    .io_mem_cluster_39_en(proc_2_io_mem_cluster_39_en),
    .io_mem_cluster_39_addr(proc_2_io_mem_cluster_39_addr),
    .io_mem_cluster_39_data(proc_2_io_mem_cluster_39_data),
    .io_mem_cluster_40_en(proc_2_io_mem_cluster_40_en),
    .io_mem_cluster_40_addr(proc_2_io_mem_cluster_40_addr),
    .io_mem_cluster_40_data(proc_2_io_mem_cluster_40_data),
    .io_mem_cluster_41_en(proc_2_io_mem_cluster_41_en),
    .io_mem_cluster_41_addr(proc_2_io_mem_cluster_41_addr),
    .io_mem_cluster_41_data(proc_2_io_mem_cluster_41_data),
    .io_mem_cluster_42_en(proc_2_io_mem_cluster_42_en),
    .io_mem_cluster_42_addr(proc_2_io_mem_cluster_42_addr),
    .io_mem_cluster_42_data(proc_2_io_mem_cluster_42_data),
    .io_mem_cluster_43_en(proc_2_io_mem_cluster_43_en),
    .io_mem_cluster_43_addr(proc_2_io_mem_cluster_43_addr),
    .io_mem_cluster_43_data(proc_2_io_mem_cluster_43_data),
    .io_mem_cluster_44_en(proc_2_io_mem_cluster_44_en),
    .io_mem_cluster_44_addr(proc_2_io_mem_cluster_44_addr),
    .io_mem_cluster_44_data(proc_2_io_mem_cluster_44_data),
    .io_mem_cluster_45_en(proc_2_io_mem_cluster_45_en),
    .io_mem_cluster_45_addr(proc_2_io_mem_cluster_45_addr),
    .io_mem_cluster_45_data(proc_2_io_mem_cluster_45_data),
    .io_mem_cluster_46_en(proc_2_io_mem_cluster_46_en),
    .io_mem_cluster_46_addr(proc_2_io_mem_cluster_46_addr),
    .io_mem_cluster_46_data(proc_2_io_mem_cluster_46_data),
    .io_mem_cluster_47_en(proc_2_io_mem_cluster_47_en),
    .io_mem_cluster_47_addr(proc_2_io_mem_cluster_47_addr),
    .io_mem_cluster_47_data(proc_2_io_mem_cluster_47_data),
    .io_mem_cluster_48_en(proc_2_io_mem_cluster_48_en),
    .io_mem_cluster_48_addr(proc_2_io_mem_cluster_48_addr),
    .io_mem_cluster_48_data(proc_2_io_mem_cluster_48_data),
    .io_mem_cluster_49_en(proc_2_io_mem_cluster_49_en),
    .io_mem_cluster_49_addr(proc_2_io_mem_cluster_49_addr),
    .io_mem_cluster_49_data(proc_2_io_mem_cluster_49_data),
    .io_mem_cluster_50_en(proc_2_io_mem_cluster_50_en),
    .io_mem_cluster_50_addr(proc_2_io_mem_cluster_50_addr),
    .io_mem_cluster_50_data(proc_2_io_mem_cluster_50_data),
    .io_mem_cluster_51_en(proc_2_io_mem_cluster_51_en),
    .io_mem_cluster_51_addr(proc_2_io_mem_cluster_51_addr),
    .io_mem_cluster_51_data(proc_2_io_mem_cluster_51_data),
    .io_mem_cluster_52_en(proc_2_io_mem_cluster_52_en),
    .io_mem_cluster_52_addr(proc_2_io_mem_cluster_52_addr),
    .io_mem_cluster_52_data(proc_2_io_mem_cluster_52_data),
    .io_mem_cluster_53_en(proc_2_io_mem_cluster_53_en),
    .io_mem_cluster_53_addr(proc_2_io_mem_cluster_53_addr),
    .io_mem_cluster_53_data(proc_2_io_mem_cluster_53_data),
    .io_mem_cluster_54_en(proc_2_io_mem_cluster_54_en),
    .io_mem_cluster_54_addr(proc_2_io_mem_cluster_54_addr),
    .io_mem_cluster_54_data(proc_2_io_mem_cluster_54_data),
    .io_mem_cluster_55_en(proc_2_io_mem_cluster_55_en),
    .io_mem_cluster_55_addr(proc_2_io_mem_cluster_55_addr),
    .io_mem_cluster_55_data(proc_2_io_mem_cluster_55_data),
    .io_mem_cluster_56_en(proc_2_io_mem_cluster_56_en),
    .io_mem_cluster_56_addr(proc_2_io_mem_cluster_56_addr),
    .io_mem_cluster_56_data(proc_2_io_mem_cluster_56_data),
    .io_mem_cluster_57_en(proc_2_io_mem_cluster_57_en),
    .io_mem_cluster_57_addr(proc_2_io_mem_cluster_57_addr),
    .io_mem_cluster_57_data(proc_2_io_mem_cluster_57_data),
    .io_mem_cluster_58_en(proc_2_io_mem_cluster_58_en),
    .io_mem_cluster_58_addr(proc_2_io_mem_cluster_58_addr),
    .io_mem_cluster_58_data(proc_2_io_mem_cluster_58_data),
    .io_mem_cluster_59_en(proc_2_io_mem_cluster_59_en),
    .io_mem_cluster_59_addr(proc_2_io_mem_cluster_59_addr),
    .io_mem_cluster_59_data(proc_2_io_mem_cluster_59_data),
    .io_mem_cluster_60_en(proc_2_io_mem_cluster_60_en),
    .io_mem_cluster_60_addr(proc_2_io_mem_cluster_60_addr),
    .io_mem_cluster_60_data(proc_2_io_mem_cluster_60_data),
    .io_mem_cluster_61_en(proc_2_io_mem_cluster_61_en),
    .io_mem_cluster_61_addr(proc_2_io_mem_cluster_61_addr),
    .io_mem_cluster_61_data(proc_2_io_mem_cluster_61_data),
    .io_mem_cluster_62_en(proc_2_io_mem_cluster_62_en),
    .io_mem_cluster_62_addr(proc_2_io_mem_cluster_62_addr),
    .io_mem_cluster_62_data(proc_2_io_mem_cluster_62_data),
    .io_mem_cluster_63_en(proc_2_io_mem_cluster_63_en),
    .io_mem_cluster_63_addr(proc_2_io_mem_cluster_63_addr),
    .io_mem_cluster_63_data(proc_2_io_mem_cluster_63_data)
  );
  Processor proc_3 ( // @[ipsa.scala 62:25]
    .clock(proc_3_clock),
    .io_pipe_phv_in_data_0(proc_3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_3_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_3_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_3_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_3_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_3_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_3_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_3_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_3_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_3_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_3_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_3_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_3_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_3_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_3_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_3_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_3_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_3_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_3_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_3_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_3_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_3_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_3_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_3_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_3_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_3_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_3_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_3_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_3_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_3_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_3_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_3_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_3_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_3_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_3_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_3_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_3_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_3_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_3_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_3_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_3_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_3_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_3_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_3_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_3_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_3_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_3_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_3_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_3_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_3_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_3_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_3_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_3_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_3_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_3_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_3_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_3_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_3_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_3_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_3_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_3_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_3_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_3_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_3_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_3_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(proc_3_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(proc_3_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(proc_3_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(proc_3_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(proc_3_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(proc_3_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(proc_3_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(proc_3_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(proc_3_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(proc_3_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(proc_3_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(proc_3_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(proc_3_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(proc_3_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(proc_3_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(proc_3_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(proc_3_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(proc_3_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(proc_3_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(proc_3_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(proc_3_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(proc_3_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(proc_3_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(proc_3_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(proc_3_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(proc_3_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(proc_3_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(proc_3_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(proc_3_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(proc_3_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(proc_3_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(proc_3_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(proc_3_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(proc_3_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(proc_3_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(proc_3_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(proc_3_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(proc_3_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(proc_3_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(proc_3_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(proc_3_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(proc_3_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(proc_3_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(proc_3_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(proc_3_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(proc_3_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(proc_3_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(proc_3_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(proc_3_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(proc_3_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(proc_3_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(proc_3_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(proc_3_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(proc_3_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(proc_3_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(proc_3_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(proc_3_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(proc_3_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(proc_3_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(proc_3_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(proc_3_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(proc_3_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(proc_3_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(proc_3_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(proc_3_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(proc_3_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(proc_3_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(proc_3_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(proc_3_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(proc_3_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(proc_3_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(proc_3_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(proc_3_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(proc_3_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(proc_3_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(proc_3_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(proc_3_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(proc_3_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(proc_3_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(proc_3_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(proc_3_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(proc_3_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(proc_3_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(proc_3_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(proc_3_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(proc_3_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(proc_3_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(proc_3_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(proc_3_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(proc_3_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(proc_3_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(proc_3_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(proc_3_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(proc_3_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(proc_3_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(proc_3_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(proc_3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(proc_3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(proc_3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(proc_3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(proc_3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(proc_3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(proc_3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(proc_3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(proc_3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(proc_3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(proc_3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(proc_3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(proc_3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(proc_3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(proc_3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(proc_3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(proc_3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(proc_3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(proc_3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(proc_3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(proc_3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_3_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_3_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_3_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_3_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_3_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_3_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_3_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_3_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_3_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_3_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_3_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_3_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_3_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_3_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_3_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_3_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_3_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_3_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_3_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_3_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_3_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_3_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_3_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_3_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_3_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_3_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_3_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_3_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_3_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_3_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_3_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_3_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_3_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_3_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_3_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_3_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_3_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_3_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_3_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_3_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_3_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_3_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_3_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_3_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_3_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_3_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_3_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_3_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_3_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_3_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_3_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_3_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_3_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_3_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_3_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_3_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_3_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_3_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_3_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_3_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_3_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_3_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_3_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_3_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(proc_3_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(proc_3_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(proc_3_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(proc_3_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(proc_3_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(proc_3_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(proc_3_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(proc_3_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(proc_3_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(proc_3_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(proc_3_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(proc_3_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(proc_3_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(proc_3_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(proc_3_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(proc_3_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(proc_3_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(proc_3_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(proc_3_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(proc_3_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(proc_3_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(proc_3_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(proc_3_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(proc_3_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(proc_3_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(proc_3_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(proc_3_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(proc_3_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(proc_3_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(proc_3_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(proc_3_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(proc_3_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(proc_3_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(proc_3_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(proc_3_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(proc_3_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(proc_3_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(proc_3_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(proc_3_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(proc_3_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(proc_3_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(proc_3_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(proc_3_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(proc_3_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(proc_3_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(proc_3_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(proc_3_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(proc_3_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(proc_3_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(proc_3_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(proc_3_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(proc_3_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(proc_3_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(proc_3_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(proc_3_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(proc_3_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(proc_3_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(proc_3_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(proc_3_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(proc_3_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(proc_3_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(proc_3_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(proc_3_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(proc_3_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(proc_3_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(proc_3_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(proc_3_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(proc_3_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(proc_3_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(proc_3_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(proc_3_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(proc_3_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(proc_3_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(proc_3_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(proc_3_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(proc_3_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(proc_3_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(proc_3_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(proc_3_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(proc_3_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(proc_3_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(proc_3_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(proc_3_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(proc_3_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(proc_3_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(proc_3_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(proc_3_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(proc_3_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(proc_3_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(proc_3_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(proc_3_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(proc_3_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(proc_3_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(proc_3_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(proc_3_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(proc_3_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(proc_3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(proc_3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(proc_3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(proc_3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(proc_3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(proc_3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(proc_3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(proc_3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(proc_3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(proc_3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(proc_3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(proc_3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(proc_3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(proc_3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(proc_3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(proc_3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(proc_3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(proc_3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(proc_3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(proc_3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_3_io_pipe_phv_out_next_config_id),
    .io_mod_par_mod_en(proc_3_io_mod_par_mod_en),
    .io_mod_par_mod_last_mau_id_mod(proc_3_io_mod_par_mod_last_mau_id_mod),
    .io_mod_par_mod_last_mau_id(proc_3_io_mod_par_mod_last_mau_id),
    .io_mod_par_mod_cs(proc_3_io_mod_par_mod_cs),
    .io_mod_par_mod_module_mod_state_id_mod(proc_3_io_mod_par_mod_module_mod_state_id_mod),
    .io_mod_par_mod_module_mod_state_id(proc_3_io_mod_par_mod_module_mod_state_id),
    .io_mod_par_mod_module_mod_sram_w_cs(proc_3_io_mod_par_mod_module_mod_sram_w_cs),
    .io_mod_par_mod_module_mod_sram_w_en(proc_3_io_mod_par_mod_module_mod_sram_w_en),
    .io_mod_par_mod_module_mod_sram_w_addr(proc_3_io_mod_par_mod_module_mod_sram_w_addr),
    .io_mod_par_mod_module_mod_sram_w_data(proc_3_io_mod_par_mod_module_mod_sram_w_data),
    .io_mod_mat_mod_en(proc_3_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_3_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_header_id(proc_3_io_mod_mat_mod_key_mod_header_id),
    .io_mod_mat_mod_key_mod_internal_offset(proc_3_io_mod_mat_mod_key_mod_internal_offset),
    .io_mod_mat_mod_key_mod_key_length(proc_3_io_mod_mat_mod_key_mod_key_length),
    .io_mod_mat_mod_table_mod_sram_id_table_0(proc_3_io_mod_mat_mod_table_mod_sram_id_table_0),
    .io_mod_mat_mod_table_mod_sram_id_table_1(proc_3_io_mod_mat_mod_table_mod_sram_id_table_1),
    .io_mod_mat_mod_table_mod_sram_id_table_2(proc_3_io_mod_mat_mod_table_mod_sram_id_table_2),
    .io_mod_mat_mod_table_mod_sram_id_table_3(proc_3_io_mod_mat_mod_table_mod_sram_id_table_3),
    .io_mod_mat_mod_table_mod_sram_id_table_4(proc_3_io_mod_mat_mod_table_mod_sram_id_table_4),
    .io_mod_mat_mod_table_mod_sram_id_table_5(proc_3_io_mod_mat_mod_table_mod_sram_id_table_5),
    .io_mod_mat_mod_table_mod_sram_id_table_6(proc_3_io_mod_mat_mod_table_mod_sram_id_table_6),
    .io_mod_mat_mod_table_mod_sram_id_table_7(proc_3_io_mod_mat_mod_table_mod_sram_id_table_7),
    .io_mod_mat_mod_table_mod_sram_id_table_8(proc_3_io_mod_mat_mod_table_mod_sram_id_table_8),
    .io_mod_mat_mod_table_mod_sram_id_table_9(proc_3_io_mod_mat_mod_table_mod_sram_id_table_9),
    .io_mod_mat_mod_table_mod_sram_id_table_10(proc_3_io_mod_mat_mod_table_mod_sram_id_table_10),
    .io_mod_mat_mod_table_mod_sram_id_table_11(proc_3_io_mod_mat_mod_table_mod_sram_id_table_11),
    .io_mod_mat_mod_table_mod_sram_id_table_12(proc_3_io_mod_mat_mod_table_mod_sram_id_table_12),
    .io_mod_mat_mod_table_mod_sram_id_table_13(proc_3_io_mod_mat_mod_table_mod_sram_id_table_13),
    .io_mod_mat_mod_table_mod_sram_id_table_14(proc_3_io_mod_mat_mod_table_mod_sram_id_table_14),
    .io_mod_mat_mod_table_mod_sram_id_table_15(proc_3_io_mod_mat_mod_table_mod_sram_id_table_15),
    .io_mod_mat_mod_table_mod_sram_id_table_16(proc_3_io_mod_mat_mod_table_mod_sram_id_table_16),
    .io_mod_mat_mod_table_mod_sram_id_table_17(proc_3_io_mod_mat_mod_table_mod_sram_id_table_17),
    .io_mod_mat_mod_table_mod_sram_id_table_18(proc_3_io_mod_mat_mod_table_mod_sram_id_table_18),
    .io_mod_mat_mod_table_mod_sram_id_table_19(proc_3_io_mod_mat_mod_table_mod_sram_id_table_19),
    .io_mod_mat_mod_table_mod_sram_id_table_20(proc_3_io_mod_mat_mod_table_mod_sram_id_table_20),
    .io_mod_mat_mod_table_mod_sram_id_table_21(proc_3_io_mod_mat_mod_table_mod_sram_id_table_21),
    .io_mod_mat_mod_table_mod_sram_id_table_22(proc_3_io_mod_mat_mod_table_mod_sram_id_table_22),
    .io_mod_mat_mod_table_mod_sram_id_table_23(proc_3_io_mod_mat_mod_table_mod_sram_id_table_23),
    .io_mod_mat_mod_table_mod_sram_id_table_24(proc_3_io_mod_mat_mod_table_mod_sram_id_table_24),
    .io_mod_mat_mod_table_mod_sram_id_table_25(proc_3_io_mod_mat_mod_table_mod_sram_id_table_25),
    .io_mod_mat_mod_table_mod_sram_id_table_26(proc_3_io_mod_mat_mod_table_mod_sram_id_table_26),
    .io_mod_mat_mod_table_mod_sram_id_table_27(proc_3_io_mod_mat_mod_table_mod_sram_id_table_27),
    .io_mod_mat_mod_table_mod_sram_id_table_28(proc_3_io_mod_mat_mod_table_mod_sram_id_table_28),
    .io_mod_mat_mod_table_mod_sram_id_table_29(proc_3_io_mod_mat_mod_table_mod_sram_id_table_29),
    .io_mod_mat_mod_table_mod_sram_id_table_30(proc_3_io_mod_mat_mod_table_mod_sram_id_table_30),
    .io_mod_mat_mod_table_mod_sram_id_table_31(proc_3_io_mod_mat_mod_table_mod_sram_id_table_31),
    .io_mod_mat_mod_table_mod_sram_id_table_32(proc_3_io_mod_mat_mod_table_mod_sram_id_table_32),
    .io_mod_mat_mod_table_mod_sram_id_table_33(proc_3_io_mod_mat_mod_table_mod_sram_id_table_33),
    .io_mod_mat_mod_table_mod_sram_id_table_34(proc_3_io_mod_mat_mod_table_mod_sram_id_table_34),
    .io_mod_mat_mod_table_mod_sram_id_table_35(proc_3_io_mod_mat_mod_table_mod_sram_id_table_35),
    .io_mod_mat_mod_table_mod_sram_id_table_36(proc_3_io_mod_mat_mod_table_mod_sram_id_table_36),
    .io_mod_mat_mod_table_mod_sram_id_table_37(proc_3_io_mod_mat_mod_table_mod_sram_id_table_37),
    .io_mod_mat_mod_table_mod_sram_id_table_38(proc_3_io_mod_mat_mod_table_mod_sram_id_table_38),
    .io_mod_mat_mod_table_mod_sram_id_table_39(proc_3_io_mod_mat_mod_table_mod_sram_id_table_39),
    .io_mod_mat_mod_table_mod_sram_id_table_40(proc_3_io_mod_mat_mod_table_mod_sram_id_table_40),
    .io_mod_mat_mod_table_mod_sram_id_table_41(proc_3_io_mod_mat_mod_table_mod_sram_id_table_41),
    .io_mod_mat_mod_table_mod_sram_id_table_42(proc_3_io_mod_mat_mod_table_mod_sram_id_table_42),
    .io_mod_mat_mod_table_mod_sram_id_table_43(proc_3_io_mod_mat_mod_table_mod_sram_id_table_43),
    .io_mod_mat_mod_table_mod_sram_id_table_44(proc_3_io_mod_mat_mod_table_mod_sram_id_table_44),
    .io_mod_mat_mod_table_mod_sram_id_table_45(proc_3_io_mod_mat_mod_table_mod_sram_id_table_45),
    .io_mod_mat_mod_table_mod_sram_id_table_46(proc_3_io_mod_mat_mod_table_mod_sram_id_table_46),
    .io_mod_mat_mod_table_mod_sram_id_table_47(proc_3_io_mod_mat_mod_table_mod_sram_id_table_47),
    .io_mod_mat_mod_table_mod_sram_id_table_48(proc_3_io_mod_mat_mod_table_mod_sram_id_table_48),
    .io_mod_mat_mod_table_mod_sram_id_table_49(proc_3_io_mod_mat_mod_table_mod_sram_id_table_49),
    .io_mod_mat_mod_table_mod_sram_id_table_50(proc_3_io_mod_mat_mod_table_mod_sram_id_table_50),
    .io_mod_mat_mod_table_mod_sram_id_table_51(proc_3_io_mod_mat_mod_table_mod_sram_id_table_51),
    .io_mod_mat_mod_table_mod_sram_id_table_52(proc_3_io_mod_mat_mod_table_mod_sram_id_table_52),
    .io_mod_mat_mod_table_mod_sram_id_table_53(proc_3_io_mod_mat_mod_table_mod_sram_id_table_53),
    .io_mod_mat_mod_table_mod_sram_id_table_54(proc_3_io_mod_mat_mod_table_mod_sram_id_table_54),
    .io_mod_mat_mod_table_mod_sram_id_table_55(proc_3_io_mod_mat_mod_table_mod_sram_id_table_55),
    .io_mod_mat_mod_table_mod_sram_id_table_56(proc_3_io_mod_mat_mod_table_mod_sram_id_table_56),
    .io_mod_mat_mod_table_mod_sram_id_table_57(proc_3_io_mod_mat_mod_table_mod_sram_id_table_57),
    .io_mod_mat_mod_table_mod_sram_id_table_58(proc_3_io_mod_mat_mod_table_mod_sram_id_table_58),
    .io_mod_mat_mod_table_mod_sram_id_table_59(proc_3_io_mod_mat_mod_table_mod_sram_id_table_59),
    .io_mod_mat_mod_table_mod_sram_id_table_60(proc_3_io_mod_mat_mod_table_mod_sram_id_table_60),
    .io_mod_mat_mod_table_mod_sram_id_table_61(proc_3_io_mod_mat_mod_table_mod_sram_id_table_61),
    .io_mod_mat_mod_table_mod_sram_id_table_62(proc_3_io_mod_mat_mod_table_mod_sram_id_table_62),
    .io_mod_mat_mod_table_mod_sram_id_table_63(proc_3_io_mod_mat_mod_table_mod_sram_id_table_63),
    .io_mod_mat_mod_table_mod_table_width(proc_3_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_table_mod_table_depth(proc_3_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_act_mod_en_0(proc_3_io_mod_act_mod_en_0),
    .io_mod_act_mod_en_1(proc_3_io_mod_act_mod_en_1),
    .io_mod_act_mod_addr(proc_3_io_mod_act_mod_addr),
    .io_mod_act_mod_data_0(proc_3_io_mod_act_mod_data_0),
    .io_mod_act_mod_data_1(proc_3_io_mod_act_mod_data_1),
    .io_mem_cluster_0_en(proc_3_io_mem_cluster_0_en),
    .io_mem_cluster_0_addr(proc_3_io_mem_cluster_0_addr),
    .io_mem_cluster_0_data(proc_3_io_mem_cluster_0_data),
    .io_mem_cluster_1_en(proc_3_io_mem_cluster_1_en),
    .io_mem_cluster_1_addr(proc_3_io_mem_cluster_1_addr),
    .io_mem_cluster_1_data(proc_3_io_mem_cluster_1_data),
    .io_mem_cluster_2_en(proc_3_io_mem_cluster_2_en),
    .io_mem_cluster_2_addr(proc_3_io_mem_cluster_2_addr),
    .io_mem_cluster_2_data(proc_3_io_mem_cluster_2_data),
    .io_mem_cluster_3_en(proc_3_io_mem_cluster_3_en),
    .io_mem_cluster_3_addr(proc_3_io_mem_cluster_3_addr),
    .io_mem_cluster_3_data(proc_3_io_mem_cluster_3_data),
    .io_mem_cluster_4_en(proc_3_io_mem_cluster_4_en),
    .io_mem_cluster_4_addr(proc_3_io_mem_cluster_4_addr),
    .io_mem_cluster_4_data(proc_3_io_mem_cluster_4_data),
    .io_mem_cluster_5_en(proc_3_io_mem_cluster_5_en),
    .io_mem_cluster_5_addr(proc_3_io_mem_cluster_5_addr),
    .io_mem_cluster_5_data(proc_3_io_mem_cluster_5_data),
    .io_mem_cluster_6_en(proc_3_io_mem_cluster_6_en),
    .io_mem_cluster_6_addr(proc_3_io_mem_cluster_6_addr),
    .io_mem_cluster_6_data(proc_3_io_mem_cluster_6_data),
    .io_mem_cluster_7_en(proc_3_io_mem_cluster_7_en),
    .io_mem_cluster_7_addr(proc_3_io_mem_cluster_7_addr),
    .io_mem_cluster_7_data(proc_3_io_mem_cluster_7_data),
    .io_mem_cluster_8_en(proc_3_io_mem_cluster_8_en),
    .io_mem_cluster_8_addr(proc_3_io_mem_cluster_8_addr),
    .io_mem_cluster_8_data(proc_3_io_mem_cluster_8_data),
    .io_mem_cluster_9_en(proc_3_io_mem_cluster_9_en),
    .io_mem_cluster_9_addr(proc_3_io_mem_cluster_9_addr),
    .io_mem_cluster_9_data(proc_3_io_mem_cluster_9_data),
    .io_mem_cluster_10_en(proc_3_io_mem_cluster_10_en),
    .io_mem_cluster_10_addr(proc_3_io_mem_cluster_10_addr),
    .io_mem_cluster_10_data(proc_3_io_mem_cluster_10_data),
    .io_mem_cluster_11_en(proc_3_io_mem_cluster_11_en),
    .io_mem_cluster_11_addr(proc_3_io_mem_cluster_11_addr),
    .io_mem_cluster_11_data(proc_3_io_mem_cluster_11_data),
    .io_mem_cluster_12_en(proc_3_io_mem_cluster_12_en),
    .io_mem_cluster_12_addr(proc_3_io_mem_cluster_12_addr),
    .io_mem_cluster_12_data(proc_3_io_mem_cluster_12_data),
    .io_mem_cluster_13_en(proc_3_io_mem_cluster_13_en),
    .io_mem_cluster_13_addr(proc_3_io_mem_cluster_13_addr),
    .io_mem_cluster_13_data(proc_3_io_mem_cluster_13_data),
    .io_mem_cluster_14_en(proc_3_io_mem_cluster_14_en),
    .io_mem_cluster_14_addr(proc_3_io_mem_cluster_14_addr),
    .io_mem_cluster_14_data(proc_3_io_mem_cluster_14_data),
    .io_mem_cluster_15_en(proc_3_io_mem_cluster_15_en),
    .io_mem_cluster_15_addr(proc_3_io_mem_cluster_15_addr),
    .io_mem_cluster_15_data(proc_3_io_mem_cluster_15_data),
    .io_mem_cluster_16_en(proc_3_io_mem_cluster_16_en),
    .io_mem_cluster_16_addr(proc_3_io_mem_cluster_16_addr),
    .io_mem_cluster_16_data(proc_3_io_mem_cluster_16_data),
    .io_mem_cluster_17_en(proc_3_io_mem_cluster_17_en),
    .io_mem_cluster_17_addr(proc_3_io_mem_cluster_17_addr),
    .io_mem_cluster_17_data(proc_3_io_mem_cluster_17_data),
    .io_mem_cluster_18_en(proc_3_io_mem_cluster_18_en),
    .io_mem_cluster_18_addr(proc_3_io_mem_cluster_18_addr),
    .io_mem_cluster_18_data(proc_3_io_mem_cluster_18_data),
    .io_mem_cluster_19_en(proc_3_io_mem_cluster_19_en),
    .io_mem_cluster_19_addr(proc_3_io_mem_cluster_19_addr),
    .io_mem_cluster_19_data(proc_3_io_mem_cluster_19_data),
    .io_mem_cluster_20_en(proc_3_io_mem_cluster_20_en),
    .io_mem_cluster_20_addr(proc_3_io_mem_cluster_20_addr),
    .io_mem_cluster_20_data(proc_3_io_mem_cluster_20_data),
    .io_mem_cluster_21_en(proc_3_io_mem_cluster_21_en),
    .io_mem_cluster_21_addr(proc_3_io_mem_cluster_21_addr),
    .io_mem_cluster_21_data(proc_3_io_mem_cluster_21_data),
    .io_mem_cluster_22_en(proc_3_io_mem_cluster_22_en),
    .io_mem_cluster_22_addr(proc_3_io_mem_cluster_22_addr),
    .io_mem_cluster_22_data(proc_3_io_mem_cluster_22_data),
    .io_mem_cluster_23_en(proc_3_io_mem_cluster_23_en),
    .io_mem_cluster_23_addr(proc_3_io_mem_cluster_23_addr),
    .io_mem_cluster_23_data(proc_3_io_mem_cluster_23_data),
    .io_mem_cluster_24_en(proc_3_io_mem_cluster_24_en),
    .io_mem_cluster_24_addr(proc_3_io_mem_cluster_24_addr),
    .io_mem_cluster_24_data(proc_3_io_mem_cluster_24_data),
    .io_mem_cluster_25_en(proc_3_io_mem_cluster_25_en),
    .io_mem_cluster_25_addr(proc_3_io_mem_cluster_25_addr),
    .io_mem_cluster_25_data(proc_3_io_mem_cluster_25_data),
    .io_mem_cluster_26_en(proc_3_io_mem_cluster_26_en),
    .io_mem_cluster_26_addr(proc_3_io_mem_cluster_26_addr),
    .io_mem_cluster_26_data(proc_3_io_mem_cluster_26_data),
    .io_mem_cluster_27_en(proc_3_io_mem_cluster_27_en),
    .io_mem_cluster_27_addr(proc_3_io_mem_cluster_27_addr),
    .io_mem_cluster_27_data(proc_3_io_mem_cluster_27_data),
    .io_mem_cluster_28_en(proc_3_io_mem_cluster_28_en),
    .io_mem_cluster_28_addr(proc_3_io_mem_cluster_28_addr),
    .io_mem_cluster_28_data(proc_3_io_mem_cluster_28_data),
    .io_mem_cluster_29_en(proc_3_io_mem_cluster_29_en),
    .io_mem_cluster_29_addr(proc_3_io_mem_cluster_29_addr),
    .io_mem_cluster_29_data(proc_3_io_mem_cluster_29_data),
    .io_mem_cluster_30_en(proc_3_io_mem_cluster_30_en),
    .io_mem_cluster_30_addr(proc_3_io_mem_cluster_30_addr),
    .io_mem_cluster_30_data(proc_3_io_mem_cluster_30_data),
    .io_mem_cluster_31_en(proc_3_io_mem_cluster_31_en),
    .io_mem_cluster_31_addr(proc_3_io_mem_cluster_31_addr),
    .io_mem_cluster_31_data(proc_3_io_mem_cluster_31_data),
    .io_mem_cluster_32_en(proc_3_io_mem_cluster_32_en),
    .io_mem_cluster_32_addr(proc_3_io_mem_cluster_32_addr),
    .io_mem_cluster_32_data(proc_3_io_mem_cluster_32_data),
    .io_mem_cluster_33_en(proc_3_io_mem_cluster_33_en),
    .io_mem_cluster_33_addr(proc_3_io_mem_cluster_33_addr),
    .io_mem_cluster_33_data(proc_3_io_mem_cluster_33_data),
    .io_mem_cluster_34_en(proc_3_io_mem_cluster_34_en),
    .io_mem_cluster_34_addr(proc_3_io_mem_cluster_34_addr),
    .io_mem_cluster_34_data(proc_3_io_mem_cluster_34_data),
    .io_mem_cluster_35_en(proc_3_io_mem_cluster_35_en),
    .io_mem_cluster_35_addr(proc_3_io_mem_cluster_35_addr),
    .io_mem_cluster_35_data(proc_3_io_mem_cluster_35_data),
    .io_mem_cluster_36_en(proc_3_io_mem_cluster_36_en),
    .io_mem_cluster_36_addr(proc_3_io_mem_cluster_36_addr),
    .io_mem_cluster_36_data(proc_3_io_mem_cluster_36_data),
    .io_mem_cluster_37_en(proc_3_io_mem_cluster_37_en),
    .io_mem_cluster_37_addr(proc_3_io_mem_cluster_37_addr),
    .io_mem_cluster_37_data(proc_3_io_mem_cluster_37_data),
    .io_mem_cluster_38_en(proc_3_io_mem_cluster_38_en),
    .io_mem_cluster_38_addr(proc_3_io_mem_cluster_38_addr),
    .io_mem_cluster_38_data(proc_3_io_mem_cluster_38_data),
    .io_mem_cluster_39_en(proc_3_io_mem_cluster_39_en),
    .io_mem_cluster_39_addr(proc_3_io_mem_cluster_39_addr),
    .io_mem_cluster_39_data(proc_3_io_mem_cluster_39_data),
    .io_mem_cluster_40_en(proc_3_io_mem_cluster_40_en),
    .io_mem_cluster_40_addr(proc_3_io_mem_cluster_40_addr),
    .io_mem_cluster_40_data(proc_3_io_mem_cluster_40_data),
    .io_mem_cluster_41_en(proc_3_io_mem_cluster_41_en),
    .io_mem_cluster_41_addr(proc_3_io_mem_cluster_41_addr),
    .io_mem_cluster_41_data(proc_3_io_mem_cluster_41_data),
    .io_mem_cluster_42_en(proc_3_io_mem_cluster_42_en),
    .io_mem_cluster_42_addr(proc_3_io_mem_cluster_42_addr),
    .io_mem_cluster_42_data(proc_3_io_mem_cluster_42_data),
    .io_mem_cluster_43_en(proc_3_io_mem_cluster_43_en),
    .io_mem_cluster_43_addr(proc_3_io_mem_cluster_43_addr),
    .io_mem_cluster_43_data(proc_3_io_mem_cluster_43_data),
    .io_mem_cluster_44_en(proc_3_io_mem_cluster_44_en),
    .io_mem_cluster_44_addr(proc_3_io_mem_cluster_44_addr),
    .io_mem_cluster_44_data(proc_3_io_mem_cluster_44_data),
    .io_mem_cluster_45_en(proc_3_io_mem_cluster_45_en),
    .io_mem_cluster_45_addr(proc_3_io_mem_cluster_45_addr),
    .io_mem_cluster_45_data(proc_3_io_mem_cluster_45_data),
    .io_mem_cluster_46_en(proc_3_io_mem_cluster_46_en),
    .io_mem_cluster_46_addr(proc_3_io_mem_cluster_46_addr),
    .io_mem_cluster_46_data(proc_3_io_mem_cluster_46_data),
    .io_mem_cluster_47_en(proc_3_io_mem_cluster_47_en),
    .io_mem_cluster_47_addr(proc_3_io_mem_cluster_47_addr),
    .io_mem_cluster_47_data(proc_3_io_mem_cluster_47_data),
    .io_mem_cluster_48_en(proc_3_io_mem_cluster_48_en),
    .io_mem_cluster_48_addr(proc_3_io_mem_cluster_48_addr),
    .io_mem_cluster_48_data(proc_3_io_mem_cluster_48_data),
    .io_mem_cluster_49_en(proc_3_io_mem_cluster_49_en),
    .io_mem_cluster_49_addr(proc_3_io_mem_cluster_49_addr),
    .io_mem_cluster_49_data(proc_3_io_mem_cluster_49_data),
    .io_mem_cluster_50_en(proc_3_io_mem_cluster_50_en),
    .io_mem_cluster_50_addr(proc_3_io_mem_cluster_50_addr),
    .io_mem_cluster_50_data(proc_3_io_mem_cluster_50_data),
    .io_mem_cluster_51_en(proc_3_io_mem_cluster_51_en),
    .io_mem_cluster_51_addr(proc_3_io_mem_cluster_51_addr),
    .io_mem_cluster_51_data(proc_3_io_mem_cluster_51_data),
    .io_mem_cluster_52_en(proc_3_io_mem_cluster_52_en),
    .io_mem_cluster_52_addr(proc_3_io_mem_cluster_52_addr),
    .io_mem_cluster_52_data(proc_3_io_mem_cluster_52_data),
    .io_mem_cluster_53_en(proc_3_io_mem_cluster_53_en),
    .io_mem_cluster_53_addr(proc_3_io_mem_cluster_53_addr),
    .io_mem_cluster_53_data(proc_3_io_mem_cluster_53_data),
    .io_mem_cluster_54_en(proc_3_io_mem_cluster_54_en),
    .io_mem_cluster_54_addr(proc_3_io_mem_cluster_54_addr),
    .io_mem_cluster_54_data(proc_3_io_mem_cluster_54_data),
    .io_mem_cluster_55_en(proc_3_io_mem_cluster_55_en),
    .io_mem_cluster_55_addr(proc_3_io_mem_cluster_55_addr),
    .io_mem_cluster_55_data(proc_3_io_mem_cluster_55_data),
    .io_mem_cluster_56_en(proc_3_io_mem_cluster_56_en),
    .io_mem_cluster_56_addr(proc_3_io_mem_cluster_56_addr),
    .io_mem_cluster_56_data(proc_3_io_mem_cluster_56_data),
    .io_mem_cluster_57_en(proc_3_io_mem_cluster_57_en),
    .io_mem_cluster_57_addr(proc_3_io_mem_cluster_57_addr),
    .io_mem_cluster_57_data(proc_3_io_mem_cluster_57_data),
    .io_mem_cluster_58_en(proc_3_io_mem_cluster_58_en),
    .io_mem_cluster_58_addr(proc_3_io_mem_cluster_58_addr),
    .io_mem_cluster_58_data(proc_3_io_mem_cluster_58_data),
    .io_mem_cluster_59_en(proc_3_io_mem_cluster_59_en),
    .io_mem_cluster_59_addr(proc_3_io_mem_cluster_59_addr),
    .io_mem_cluster_59_data(proc_3_io_mem_cluster_59_data),
    .io_mem_cluster_60_en(proc_3_io_mem_cluster_60_en),
    .io_mem_cluster_60_addr(proc_3_io_mem_cluster_60_addr),
    .io_mem_cluster_60_data(proc_3_io_mem_cluster_60_data),
    .io_mem_cluster_61_en(proc_3_io_mem_cluster_61_en),
    .io_mem_cluster_61_addr(proc_3_io_mem_cluster_61_addr),
    .io_mem_cluster_61_data(proc_3_io_mem_cluster_61_data),
    .io_mem_cluster_62_en(proc_3_io_mem_cluster_62_en),
    .io_mem_cluster_62_addr(proc_3_io_mem_cluster_62_addr),
    .io_mem_cluster_62_data(proc_3_io_mem_cluster_62_data),
    .io_mem_cluster_63_en(proc_3_io_mem_cluster_63_en),
    .io_mem_cluster_63_addr(proc_3_io_mem_cluster_63_addr),
    .io_mem_cluster_63_data(proc_3_io_mem_cluster_63_data)
  );
  SRAMCluster sram_cluster_0 ( // @[ipsa.scala 68:25]
    .clock(sram_cluster_0_clock),
    .io_w_wcs(sram_cluster_0_io_w_wcs),
    .io_w_w_en(sram_cluster_0_io_w_w_en),
    .io_w_w_addr(sram_cluster_0_io_w_w_addr),
    .io_w_w_data(sram_cluster_0_io_w_w_data),
    .io_r_0_cluster_0_en(sram_cluster_0_io_r_0_cluster_0_en),
    .io_r_0_cluster_0_addr(sram_cluster_0_io_r_0_cluster_0_addr),
    .io_r_0_cluster_0_data(sram_cluster_0_io_r_0_cluster_0_data),
    .io_r_0_cluster_1_en(sram_cluster_0_io_r_0_cluster_1_en),
    .io_r_0_cluster_1_addr(sram_cluster_0_io_r_0_cluster_1_addr),
    .io_r_0_cluster_1_data(sram_cluster_0_io_r_0_cluster_1_data),
    .io_r_0_cluster_2_en(sram_cluster_0_io_r_0_cluster_2_en),
    .io_r_0_cluster_2_addr(sram_cluster_0_io_r_0_cluster_2_addr),
    .io_r_0_cluster_2_data(sram_cluster_0_io_r_0_cluster_2_data),
    .io_r_0_cluster_3_en(sram_cluster_0_io_r_0_cluster_3_en),
    .io_r_0_cluster_3_addr(sram_cluster_0_io_r_0_cluster_3_addr),
    .io_r_0_cluster_3_data(sram_cluster_0_io_r_0_cluster_3_data),
    .io_r_0_cluster_4_en(sram_cluster_0_io_r_0_cluster_4_en),
    .io_r_0_cluster_4_addr(sram_cluster_0_io_r_0_cluster_4_addr),
    .io_r_0_cluster_4_data(sram_cluster_0_io_r_0_cluster_4_data),
    .io_r_0_cluster_5_en(sram_cluster_0_io_r_0_cluster_5_en),
    .io_r_0_cluster_5_addr(sram_cluster_0_io_r_0_cluster_5_addr),
    .io_r_0_cluster_5_data(sram_cluster_0_io_r_0_cluster_5_data),
    .io_r_0_cluster_6_en(sram_cluster_0_io_r_0_cluster_6_en),
    .io_r_0_cluster_6_addr(sram_cluster_0_io_r_0_cluster_6_addr),
    .io_r_0_cluster_6_data(sram_cluster_0_io_r_0_cluster_6_data),
    .io_r_0_cluster_7_en(sram_cluster_0_io_r_0_cluster_7_en),
    .io_r_0_cluster_7_addr(sram_cluster_0_io_r_0_cluster_7_addr),
    .io_r_0_cluster_7_data(sram_cluster_0_io_r_0_cluster_7_data),
    .io_r_0_cluster_8_en(sram_cluster_0_io_r_0_cluster_8_en),
    .io_r_0_cluster_8_addr(sram_cluster_0_io_r_0_cluster_8_addr),
    .io_r_0_cluster_8_data(sram_cluster_0_io_r_0_cluster_8_data),
    .io_r_0_cluster_9_en(sram_cluster_0_io_r_0_cluster_9_en),
    .io_r_0_cluster_9_addr(sram_cluster_0_io_r_0_cluster_9_addr),
    .io_r_0_cluster_9_data(sram_cluster_0_io_r_0_cluster_9_data),
    .io_r_0_cluster_10_en(sram_cluster_0_io_r_0_cluster_10_en),
    .io_r_0_cluster_10_addr(sram_cluster_0_io_r_0_cluster_10_addr),
    .io_r_0_cluster_10_data(sram_cluster_0_io_r_0_cluster_10_data),
    .io_r_0_cluster_11_en(sram_cluster_0_io_r_0_cluster_11_en),
    .io_r_0_cluster_11_addr(sram_cluster_0_io_r_0_cluster_11_addr),
    .io_r_0_cluster_11_data(sram_cluster_0_io_r_0_cluster_11_data),
    .io_r_0_cluster_12_en(sram_cluster_0_io_r_0_cluster_12_en),
    .io_r_0_cluster_12_addr(sram_cluster_0_io_r_0_cluster_12_addr),
    .io_r_0_cluster_12_data(sram_cluster_0_io_r_0_cluster_12_data),
    .io_r_0_cluster_13_en(sram_cluster_0_io_r_0_cluster_13_en),
    .io_r_0_cluster_13_addr(sram_cluster_0_io_r_0_cluster_13_addr),
    .io_r_0_cluster_13_data(sram_cluster_0_io_r_0_cluster_13_data),
    .io_r_0_cluster_14_en(sram_cluster_0_io_r_0_cluster_14_en),
    .io_r_0_cluster_14_addr(sram_cluster_0_io_r_0_cluster_14_addr),
    .io_r_0_cluster_14_data(sram_cluster_0_io_r_0_cluster_14_data),
    .io_r_0_cluster_15_en(sram_cluster_0_io_r_0_cluster_15_en),
    .io_r_0_cluster_15_addr(sram_cluster_0_io_r_0_cluster_15_addr),
    .io_r_0_cluster_15_data(sram_cluster_0_io_r_0_cluster_15_data),
    .io_r_0_cluster_16_en(sram_cluster_0_io_r_0_cluster_16_en),
    .io_r_0_cluster_16_addr(sram_cluster_0_io_r_0_cluster_16_addr),
    .io_r_0_cluster_16_data(sram_cluster_0_io_r_0_cluster_16_data),
    .io_r_0_cluster_17_en(sram_cluster_0_io_r_0_cluster_17_en),
    .io_r_0_cluster_17_addr(sram_cluster_0_io_r_0_cluster_17_addr),
    .io_r_0_cluster_17_data(sram_cluster_0_io_r_0_cluster_17_data),
    .io_r_0_cluster_18_en(sram_cluster_0_io_r_0_cluster_18_en),
    .io_r_0_cluster_18_addr(sram_cluster_0_io_r_0_cluster_18_addr),
    .io_r_0_cluster_18_data(sram_cluster_0_io_r_0_cluster_18_data),
    .io_r_0_cluster_19_en(sram_cluster_0_io_r_0_cluster_19_en),
    .io_r_0_cluster_19_addr(sram_cluster_0_io_r_0_cluster_19_addr),
    .io_r_0_cluster_19_data(sram_cluster_0_io_r_0_cluster_19_data),
    .io_r_0_cluster_20_en(sram_cluster_0_io_r_0_cluster_20_en),
    .io_r_0_cluster_20_addr(sram_cluster_0_io_r_0_cluster_20_addr),
    .io_r_0_cluster_20_data(sram_cluster_0_io_r_0_cluster_20_data),
    .io_r_0_cluster_21_en(sram_cluster_0_io_r_0_cluster_21_en),
    .io_r_0_cluster_21_addr(sram_cluster_0_io_r_0_cluster_21_addr),
    .io_r_0_cluster_21_data(sram_cluster_0_io_r_0_cluster_21_data),
    .io_r_0_cluster_22_en(sram_cluster_0_io_r_0_cluster_22_en),
    .io_r_0_cluster_22_addr(sram_cluster_0_io_r_0_cluster_22_addr),
    .io_r_0_cluster_22_data(sram_cluster_0_io_r_0_cluster_22_data),
    .io_r_0_cluster_23_en(sram_cluster_0_io_r_0_cluster_23_en),
    .io_r_0_cluster_23_addr(sram_cluster_0_io_r_0_cluster_23_addr),
    .io_r_0_cluster_23_data(sram_cluster_0_io_r_0_cluster_23_data),
    .io_r_0_cluster_24_en(sram_cluster_0_io_r_0_cluster_24_en),
    .io_r_0_cluster_24_addr(sram_cluster_0_io_r_0_cluster_24_addr),
    .io_r_0_cluster_24_data(sram_cluster_0_io_r_0_cluster_24_data),
    .io_r_0_cluster_25_en(sram_cluster_0_io_r_0_cluster_25_en),
    .io_r_0_cluster_25_addr(sram_cluster_0_io_r_0_cluster_25_addr),
    .io_r_0_cluster_25_data(sram_cluster_0_io_r_0_cluster_25_data),
    .io_r_0_cluster_26_en(sram_cluster_0_io_r_0_cluster_26_en),
    .io_r_0_cluster_26_addr(sram_cluster_0_io_r_0_cluster_26_addr),
    .io_r_0_cluster_26_data(sram_cluster_0_io_r_0_cluster_26_data),
    .io_r_0_cluster_27_en(sram_cluster_0_io_r_0_cluster_27_en),
    .io_r_0_cluster_27_addr(sram_cluster_0_io_r_0_cluster_27_addr),
    .io_r_0_cluster_27_data(sram_cluster_0_io_r_0_cluster_27_data),
    .io_r_0_cluster_28_en(sram_cluster_0_io_r_0_cluster_28_en),
    .io_r_0_cluster_28_addr(sram_cluster_0_io_r_0_cluster_28_addr),
    .io_r_0_cluster_28_data(sram_cluster_0_io_r_0_cluster_28_data),
    .io_r_0_cluster_29_en(sram_cluster_0_io_r_0_cluster_29_en),
    .io_r_0_cluster_29_addr(sram_cluster_0_io_r_0_cluster_29_addr),
    .io_r_0_cluster_29_data(sram_cluster_0_io_r_0_cluster_29_data),
    .io_r_0_cluster_30_en(sram_cluster_0_io_r_0_cluster_30_en),
    .io_r_0_cluster_30_addr(sram_cluster_0_io_r_0_cluster_30_addr),
    .io_r_0_cluster_30_data(sram_cluster_0_io_r_0_cluster_30_data),
    .io_r_0_cluster_31_en(sram_cluster_0_io_r_0_cluster_31_en),
    .io_r_0_cluster_31_addr(sram_cluster_0_io_r_0_cluster_31_addr),
    .io_r_0_cluster_31_data(sram_cluster_0_io_r_0_cluster_31_data),
    .io_r_0_cluster_32_en(sram_cluster_0_io_r_0_cluster_32_en),
    .io_r_0_cluster_32_addr(sram_cluster_0_io_r_0_cluster_32_addr),
    .io_r_0_cluster_32_data(sram_cluster_0_io_r_0_cluster_32_data),
    .io_r_0_cluster_33_en(sram_cluster_0_io_r_0_cluster_33_en),
    .io_r_0_cluster_33_addr(sram_cluster_0_io_r_0_cluster_33_addr),
    .io_r_0_cluster_33_data(sram_cluster_0_io_r_0_cluster_33_data),
    .io_r_0_cluster_34_en(sram_cluster_0_io_r_0_cluster_34_en),
    .io_r_0_cluster_34_addr(sram_cluster_0_io_r_0_cluster_34_addr),
    .io_r_0_cluster_34_data(sram_cluster_0_io_r_0_cluster_34_data),
    .io_r_0_cluster_35_en(sram_cluster_0_io_r_0_cluster_35_en),
    .io_r_0_cluster_35_addr(sram_cluster_0_io_r_0_cluster_35_addr),
    .io_r_0_cluster_35_data(sram_cluster_0_io_r_0_cluster_35_data),
    .io_r_0_cluster_36_en(sram_cluster_0_io_r_0_cluster_36_en),
    .io_r_0_cluster_36_addr(sram_cluster_0_io_r_0_cluster_36_addr),
    .io_r_0_cluster_36_data(sram_cluster_0_io_r_0_cluster_36_data),
    .io_r_0_cluster_37_en(sram_cluster_0_io_r_0_cluster_37_en),
    .io_r_0_cluster_37_addr(sram_cluster_0_io_r_0_cluster_37_addr),
    .io_r_0_cluster_37_data(sram_cluster_0_io_r_0_cluster_37_data),
    .io_r_0_cluster_38_en(sram_cluster_0_io_r_0_cluster_38_en),
    .io_r_0_cluster_38_addr(sram_cluster_0_io_r_0_cluster_38_addr),
    .io_r_0_cluster_38_data(sram_cluster_0_io_r_0_cluster_38_data),
    .io_r_0_cluster_39_en(sram_cluster_0_io_r_0_cluster_39_en),
    .io_r_0_cluster_39_addr(sram_cluster_0_io_r_0_cluster_39_addr),
    .io_r_0_cluster_39_data(sram_cluster_0_io_r_0_cluster_39_data),
    .io_r_0_cluster_40_en(sram_cluster_0_io_r_0_cluster_40_en),
    .io_r_0_cluster_40_addr(sram_cluster_0_io_r_0_cluster_40_addr),
    .io_r_0_cluster_40_data(sram_cluster_0_io_r_0_cluster_40_data),
    .io_r_0_cluster_41_en(sram_cluster_0_io_r_0_cluster_41_en),
    .io_r_0_cluster_41_addr(sram_cluster_0_io_r_0_cluster_41_addr),
    .io_r_0_cluster_41_data(sram_cluster_0_io_r_0_cluster_41_data),
    .io_r_0_cluster_42_en(sram_cluster_0_io_r_0_cluster_42_en),
    .io_r_0_cluster_42_addr(sram_cluster_0_io_r_0_cluster_42_addr),
    .io_r_0_cluster_42_data(sram_cluster_0_io_r_0_cluster_42_data),
    .io_r_0_cluster_43_en(sram_cluster_0_io_r_0_cluster_43_en),
    .io_r_0_cluster_43_addr(sram_cluster_0_io_r_0_cluster_43_addr),
    .io_r_0_cluster_43_data(sram_cluster_0_io_r_0_cluster_43_data),
    .io_r_0_cluster_44_en(sram_cluster_0_io_r_0_cluster_44_en),
    .io_r_0_cluster_44_addr(sram_cluster_0_io_r_0_cluster_44_addr),
    .io_r_0_cluster_44_data(sram_cluster_0_io_r_0_cluster_44_data),
    .io_r_0_cluster_45_en(sram_cluster_0_io_r_0_cluster_45_en),
    .io_r_0_cluster_45_addr(sram_cluster_0_io_r_0_cluster_45_addr),
    .io_r_0_cluster_45_data(sram_cluster_0_io_r_0_cluster_45_data),
    .io_r_0_cluster_46_en(sram_cluster_0_io_r_0_cluster_46_en),
    .io_r_0_cluster_46_addr(sram_cluster_0_io_r_0_cluster_46_addr),
    .io_r_0_cluster_46_data(sram_cluster_0_io_r_0_cluster_46_data),
    .io_r_0_cluster_47_en(sram_cluster_0_io_r_0_cluster_47_en),
    .io_r_0_cluster_47_addr(sram_cluster_0_io_r_0_cluster_47_addr),
    .io_r_0_cluster_47_data(sram_cluster_0_io_r_0_cluster_47_data),
    .io_r_0_cluster_48_en(sram_cluster_0_io_r_0_cluster_48_en),
    .io_r_0_cluster_48_addr(sram_cluster_0_io_r_0_cluster_48_addr),
    .io_r_0_cluster_48_data(sram_cluster_0_io_r_0_cluster_48_data),
    .io_r_0_cluster_49_en(sram_cluster_0_io_r_0_cluster_49_en),
    .io_r_0_cluster_49_addr(sram_cluster_0_io_r_0_cluster_49_addr),
    .io_r_0_cluster_49_data(sram_cluster_0_io_r_0_cluster_49_data),
    .io_r_0_cluster_50_en(sram_cluster_0_io_r_0_cluster_50_en),
    .io_r_0_cluster_50_addr(sram_cluster_0_io_r_0_cluster_50_addr),
    .io_r_0_cluster_50_data(sram_cluster_0_io_r_0_cluster_50_data),
    .io_r_0_cluster_51_en(sram_cluster_0_io_r_0_cluster_51_en),
    .io_r_0_cluster_51_addr(sram_cluster_0_io_r_0_cluster_51_addr),
    .io_r_0_cluster_51_data(sram_cluster_0_io_r_0_cluster_51_data),
    .io_r_0_cluster_52_en(sram_cluster_0_io_r_0_cluster_52_en),
    .io_r_0_cluster_52_addr(sram_cluster_0_io_r_0_cluster_52_addr),
    .io_r_0_cluster_52_data(sram_cluster_0_io_r_0_cluster_52_data),
    .io_r_0_cluster_53_en(sram_cluster_0_io_r_0_cluster_53_en),
    .io_r_0_cluster_53_addr(sram_cluster_0_io_r_0_cluster_53_addr),
    .io_r_0_cluster_53_data(sram_cluster_0_io_r_0_cluster_53_data),
    .io_r_0_cluster_54_en(sram_cluster_0_io_r_0_cluster_54_en),
    .io_r_0_cluster_54_addr(sram_cluster_0_io_r_0_cluster_54_addr),
    .io_r_0_cluster_54_data(sram_cluster_0_io_r_0_cluster_54_data),
    .io_r_0_cluster_55_en(sram_cluster_0_io_r_0_cluster_55_en),
    .io_r_0_cluster_55_addr(sram_cluster_0_io_r_0_cluster_55_addr),
    .io_r_0_cluster_55_data(sram_cluster_0_io_r_0_cluster_55_data),
    .io_r_0_cluster_56_en(sram_cluster_0_io_r_0_cluster_56_en),
    .io_r_0_cluster_56_addr(sram_cluster_0_io_r_0_cluster_56_addr),
    .io_r_0_cluster_56_data(sram_cluster_0_io_r_0_cluster_56_data),
    .io_r_0_cluster_57_en(sram_cluster_0_io_r_0_cluster_57_en),
    .io_r_0_cluster_57_addr(sram_cluster_0_io_r_0_cluster_57_addr),
    .io_r_0_cluster_57_data(sram_cluster_0_io_r_0_cluster_57_data),
    .io_r_0_cluster_58_en(sram_cluster_0_io_r_0_cluster_58_en),
    .io_r_0_cluster_58_addr(sram_cluster_0_io_r_0_cluster_58_addr),
    .io_r_0_cluster_58_data(sram_cluster_0_io_r_0_cluster_58_data),
    .io_r_0_cluster_59_en(sram_cluster_0_io_r_0_cluster_59_en),
    .io_r_0_cluster_59_addr(sram_cluster_0_io_r_0_cluster_59_addr),
    .io_r_0_cluster_59_data(sram_cluster_0_io_r_0_cluster_59_data),
    .io_r_0_cluster_60_en(sram_cluster_0_io_r_0_cluster_60_en),
    .io_r_0_cluster_60_addr(sram_cluster_0_io_r_0_cluster_60_addr),
    .io_r_0_cluster_60_data(sram_cluster_0_io_r_0_cluster_60_data),
    .io_r_0_cluster_61_en(sram_cluster_0_io_r_0_cluster_61_en),
    .io_r_0_cluster_61_addr(sram_cluster_0_io_r_0_cluster_61_addr),
    .io_r_0_cluster_61_data(sram_cluster_0_io_r_0_cluster_61_data),
    .io_r_0_cluster_62_en(sram_cluster_0_io_r_0_cluster_62_en),
    .io_r_0_cluster_62_addr(sram_cluster_0_io_r_0_cluster_62_addr),
    .io_r_0_cluster_62_data(sram_cluster_0_io_r_0_cluster_62_data),
    .io_r_0_cluster_63_en(sram_cluster_0_io_r_0_cluster_63_en),
    .io_r_0_cluster_63_addr(sram_cluster_0_io_r_0_cluster_63_addr),
    .io_r_0_cluster_63_data(sram_cluster_0_io_r_0_cluster_63_data),
    .io_r_1_cluster_0_en(sram_cluster_0_io_r_1_cluster_0_en),
    .io_r_1_cluster_0_addr(sram_cluster_0_io_r_1_cluster_0_addr),
    .io_r_1_cluster_0_data(sram_cluster_0_io_r_1_cluster_0_data),
    .io_r_1_cluster_1_en(sram_cluster_0_io_r_1_cluster_1_en),
    .io_r_1_cluster_1_addr(sram_cluster_0_io_r_1_cluster_1_addr),
    .io_r_1_cluster_1_data(sram_cluster_0_io_r_1_cluster_1_data),
    .io_r_1_cluster_2_en(sram_cluster_0_io_r_1_cluster_2_en),
    .io_r_1_cluster_2_addr(sram_cluster_0_io_r_1_cluster_2_addr),
    .io_r_1_cluster_2_data(sram_cluster_0_io_r_1_cluster_2_data),
    .io_r_1_cluster_3_en(sram_cluster_0_io_r_1_cluster_3_en),
    .io_r_1_cluster_3_addr(sram_cluster_0_io_r_1_cluster_3_addr),
    .io_r_1_cluster_3_data(sram_cluster_0_io_r_1_cluster_3_data),
    .io_r_1_cluster_4_en(sram_cluster_0_io_r_1_cluster_4_en),
    .io_r_1_cluster_4_addr(sram_cluster_0_io_r_1_cluster_4_addr),
    .io_r_1_cluster_4_data(sram_cluster_0_io_r_1_cluster_4_data),
    .io_r_1_cluster_5_en(sram_cluster_0_io_r_1_cluster_5_en),
    .io_r_1_cluster_5_addr(sram_cluster_0_io_r_1_cluster_5_addr),
    .io_r_1_cluster_5_data(sram_cluster_0_io_r_1_cluster_5_data),
    .io_r_1_cluster_6_en(sram_cluster_0_io_r_1_cluster_6_en),
    .io_r_1_cluster_6_addr(sram_cluster_0_io_r_1_cluster_6_addr),
    .io_r_1_cluster_6_data(sram_cluster_0_io_r_1_cluster_6_data),
    .io_r_1_cluster_7_en(sram_cluster_0_io_r_1_cluster_7_en),
    .io_r_1_cluster_7_addr(sram_cluster_0_io_r_1_cluster_7_addr),
    .io_r_1_cluster_7_data(sram_cluster_0_io_r_1_cluster_7_data),
    .io_r_1_cluster_8_en(sram_cluster_0_io_r_1_cluster_8_en),
    .io_r_1_cluster_8_addr(sram_cluster_0_io_r_1_cluster_8_addr),
    .io_r_1_cluster_8_data(sram_cluster_0_io_r_1_cluster_8_data),
    .io_r_1_cluster_9_en(sram_cluster_0_io_r_1_cluster_9_en),
    .io_r_1_cluster_9_addr(sram_cluster_0_io_r_1_cluster_9_addr),
    .io_r_1_cluster_9_data(sram_cluster_0_io_r_1_cluster_9_data),
    .io_r_1_cluster_10_en(sram_cluster_0_io_r_1_cluster_10_en),
    .io_r_1_cluster_10_addr(sram_cluster_0_io_r_1_cluster_10_addr),
    .io_r_1_cluster_10_data(sram_cluster_0_io_r_1_cluster_10_data),
    .io_r_1_cluster_11_en(sram_cluster_0_io_r_1_cluster_11_en),
    .io_r_1_cluster_11_addr(sram_cluster_0_io_r_1_cluster_11_addr),
    .io_r_1_cluster_11_data(sram_cluster_0_io_r_1_cluster_11_data),
    .io_r_1_cluster_12_en(sram_cluster_0_io_r_1_cluster_12_en),
    .io_r_1_cluster_12_addr(sram_cluster_0_io_r_1_cluster_12_addr),
    .io_r_1_cluster_12_data(sram_cluster_0_io_r_1_cluster_12_data),
    .io_r_1_cluster_13_en(sram_cluster_0_io_r_1_cluster_13_en),
    .io_r_1_cluster_13_addr(sram_cluster_0_io_r_1_cluster_13_addr),
    .io_r_1_cluster_13_data(sram_cluster_0_io_r_1_cluster_13_data),
    .io_r_1_cluster_14_en(sram_cluster_0_io_r_1_cluster_14_en),
    .io_r_1_cluster_14_addr(sram_cluster_0_io_r_1_cluster_14_addr),
    .io_r_1_cluster_14_data(sram_cluster_0_io_r_1_cluster_14_data),
    .io_r_1_cluster_15_en(sram_cluster_0_io_r_1_cluster_15_en),
    .io_r_1_cluster_15_addr(sram_cluster_0_io_r_1_cluster_15_addr),
    .io_r_1_cluster_15_data(sram_cluster_0_io_r_1_cluster_15_data),
    .io_r_1_cluster_16_en(sram_cluster_0_io_r_1_cluster_16_en),
    .io_r_1_cluster_16_addr(sram_cluster_0_io_r_1_cluster_16_addr),
    .io_r_1_cluster_16_data(sram_cluster_0_io_r_1_cluster_16_data),
    .io_r_1_cluster_17_en(sram_cluster_0_io_r_1_cluster_17_en),
    .io_r_1_cluster_17_addr(sram_cluster_0_io_r_1_cluster_17_addr),
    .io_r_1_cluster_17_data(sram_cluster_0_io_r_1_cluster_17_data),
    .io_r_1_cluster_18_en(sram_cluster_0_io_r_1_cluster_18_en),
    .io_r_1_cluster_18_addr(sram_cluster_0_io_r_1_cluster_18_addr),
    .io_r_1_cluster_18_data(sram_cluster_0_io_r_1_cluster_18_data),
    .io_r_1_cluster_19_en(sram_cluster_0_io_r_1_cluster_19_en),
    .io_r_1_cluster_19_addr(sram_cluster_0_io_r_1_cluster_19_addr),
    .io_r_1_cluster_19_data(sram_cluster_0_io_r_1_cluster_19_data),
    .io_r_1_cluster_20_en(sram_cluster_0_io_r_1_cluster_20_en),
    .io_r_1_cluster_20_addr(sram_cluster_0_io_r_1_cluster_20_addr),
    .io_r_1_cluster_20_data(sram_cluster_0_io_r_1_cluster_20_data),
    .io_r_1_cluster_21_en(sram_cluster_0_io_r_1_cluster_21_en),
    .io_r_1_cluster_21_addr(sram_cluster_0_io_r_1_cluster_21_addr),
    .io_r_1_cluster_21_data(sram_cluster_0_io_r_1_cluster_21_data),
    .io_r_1_cluster_22_en(sram_cluster_0_io_r_1_cluster_22_en),
    .io_r_1_cluster_22_addr(sram_cluster_0_io_r_1_cluster_22_addr),
    .io_r_1_cluster_22_data(sram_cluster_0_io_r_1_cluster_22_data),
    .io_r_1_cluster_23_en(sram_cluster_0_io_r_1_cluster_23_en),
    .io_r_1_cluster_23_addr(sram_cluster_0_io_r_1_cluster_23_addr),
    .io_r_1_cluster_23_data(sram_cluster_0_io_r_1_cluster_23_data),
    .io_r_1_cluster_24_en(sram_cluster_0_io_r_1_cluster_24_en),
    .io_r_1_cluster_24_addr(sram_cluster_0_io_r_1_cluster_24_addr),
    .io_r_1_cluster_24_data(sram_cluster_0_io_r_1_cluster_24_data),
    .io_r_1_cluster_25_en(sram_cluster_0_io_r_1_cluster_25_en),
    .io_r_1_cluster_25_addr(sram_cluster_0_io_r_1_cluster_25_addr),
    .io_r_1_cluster_25_data(sram_cluster_0_io_r_1_cluster_25_data),
    .io_r_1_cluster_26_en(sram_cluster_0_io_r_1_cluster_26_en),
    .io_r_1_cluster_26_addr(sram_cluster_0_io_r_1_cluster_26_addr),
    .io_r_1_cluster_26_data(sram_cluster_0_io_r_1_cluster_26_data),
    .io_r_1_cluster_27_en(sram_cluster_0_io_r_1_cluster_27_en),
    .io_r_1_cluster_27_addr(sram_cluster_0_io_r_1_cluster_27_addr),
    .io_r_1_cluster_27_data(sram_cluster_0_io_r_1_cluster_27_data),
    .io_r_1_cluster_28_en(sram_cluster_0_io_r_1_cluster_28_en),
    .io_r_1_cluster_28_addr(sram_cluster_0_io_r_1_cluster_28_addr),
    .io_r_1_cluster_28_data(sram_cluster_0_io_r_1_cluster_28_data),
    .io_r_1_cluster_29_en(sram_cluster_0_io_r_1_cluster_29_en),
    .io_r_1_cluster_29_addr(sram_cluster_0_io_r_1_cluster_29_addr),
    .io_r_1_cluster_29_data(sram_cluster_0_io_r_1_cluster_29_data),
    .io_r_1_cluster_30_en(sram_cluster_0_io_r_1_cluster_30_en),
    .io_r_1_cluster_30_addr(sram_cluster_0_io_r_1_cluster_30_addr),
    .io_r_1_cluster_30_data(sram_cluster_0_io_r_1_cluster_30_data),
    .io_r_1_cluster_31_en(sram_cluster_0_io_r_1_cluster_31_en),
    .io_r_1_cluster_31_addr(sram_cluster_0_io_r_1_cluster_31_addr),
    .io_r_1_cluster_31_data(sram_cluster_0_io_r_1_cluster_31_data),
    .io_r_1_cluster_32_en(sram_cluster_0_io_r_1_cluster_32_en),
    .io_r_1_cluster_32_addr(sram_cluster_0_io_r_1_cluster_32_addr),
    .io_r_1_cluster_32_data(sram_cluster_0_io_r_1_cluster_32_data),
    .io_r_1_cluster_33_en(sram_cluster_0_io_r_1_cluster_33_en),
    .io_r_1_cluster_33_addr(sram_cluster_0_io_r_1_cluster_33_addr),
    .io_r_1_cluster_33_data(sram_cluster_0_io_r_1_cluster_33_data),
    .io_r_1_cluster_34_en(sram_cluster_0_io_r_1_cluster_34_en),
    .io_r_1_cluster_34_addr(sram_cluster_0_io_r_1_cluster_34_addr),
    .io_r_1_cluster_34_data(sram_cluster_0_io_r_1_cluster_34_data),
    .io_r_1_cluster_35_en(sram_cluster_0_io_r_1_cluster_35_en),
    .io_r_1_cluster_35_addr(sram_cluster_0_io_r_1_cluster_35_addr),
    .io_r_1_cluster_35_data(sram_cluster_0_io_r_1_cluster_35_data),
    .io_r_1_cluster_36_en(sram_cluster_0_io_r_1_cluster_36_en),
    .io_r_1_cluster_36_addr(sram_cluster_0_io_r_1_cluster_36_addr),
    .io_r_1_cluster_36_data(sram_cluster_0_io_r_1_cluster_36_data),
    .io_r_1_cluster_37_en(sram_cluster_0_io_r_1_cluster_37_en),
    .io_r_1_cluster_37_addr(sram_cluster_0_io_r_1_cluster_37_addr),
    .io_r_1_cluster_37_data(sram_cluster_0_io_r_1_cluster_37_data),
    .io_r_1_cluster_38_en(sram_cluster_0_io_r_1_cluster_38_en),
    .io_r_1_cluster_38_addr(sram_cluster_0_io_r_1_cluster_38_addr),
    .io_r_1_cluster_38_data(sram_cluster_0_io_r_1_cluster_38_data),
    .io_r_1_cluster_39_en(sram_cluster_0_io_r_1_cluster_39_en),
    .io_r_1_cluster_39_addr(sram_cluster_0_io_r_1_cluster_39_addr),
    .io_r_1_cluster_39_data(sram_cluster_0_io_r_1_cluster_39_data),
    .io_r_1_cluster_40_en(sram_cluster_0_io_r_1_cluster_40_en),
    .io_r_1_cluster_40_addr(sram_cluster_0_io_r_1_cluster_40_addr),
    .io_r_1_cluster_40_data(sram_cluster_0_io_r_1_cluster_40_data),
    .io_r_1_cluster_41_en(sram_cluster_0_io_r_1_cluster_41_en),
    .io_r_1_cluster_41_addr(sram_cluster_0_io_r_1_cluster_41_addr),
    .io_r_1_cluster_41_data(sram_cluster_0_io_r_1_cluster_41_data),
    .io_r_1_cluster_42_en(sram_cluster_0_io_r_1_cluster_42_en),
    .io_r_1_cluster_42_addr(sram_cluster_0_io_r_1_cluster_42_addr),
    .io_r_1_cluster_42_data(sram_cluster_0_io_r_1_cluster_42_data),
    .io_r_1_cluster_43_en(sram_cluster_0_io_r_1_cluster_43_en),
    .io_r_1_cluster_43_addr(sram_cluster_0_io_r_1_cluster_43_addr),
    .io_r_1_cluster_43_data(sram_cluster_0_io_r_1_cluster_43_data),
    .io_r_1_cluster_44_en(sram_cluster_0_io_r_1_cluster_44_en),
    .io_r_1_cluster_44_addr(sram_cluster_0_io_r_1_cluster_44_addr),
    .io_r_1_cluster_44_data(sram_cluster_0_io_r_1_cluster_44_data),
    .io_r_1_cluster_45_en(sram_cluster_0_io_r_1_cluster_45_en),
    .io_r_1_cluster_45_addr(sram_cluster_0_io_r_1_cluster_45_addr),
    .io_r_1_cluster_45_data(sram_cluster_0_io_r_1_cluster_45_data),
    .io_r_1_cluster_46_en(sram_cluster_0_io_r_1_cluster_46_en),
    .io_r_1_cluster_46_addr(sram_cluster_0_io_r_1_cluster_46_addr),
    .io_r_1_cluster_46_data(sram_cluster_0_io_r_1_cluster_46_data),
    .io_r_1_cluster_47_en(sram_cluster_0_io_r_1_cluster_47_en),
    .io_r_1_cluster_47_addr(sram_cluster_0_io_r_1_cluster_47_addr),
    .io_r_1_cluster_47_data(sram_cluster_0_io_r_1_cluster_47_data),
    .io_r_1_cluster_48_en(sram_cluster_0_io_r_1_cluster_48_en),
    .io_r_1_cluster_48_addr(sram_cluster_0_io_r_1_cluster_48_addr),
    .io_r_1_cluster_48_data(sram_cluster_0_io_r_1_cluster_48_data),
    .io_r_1_cluster_49_en(sram_cluster_0_io_r_1_cluster_49_en),
    .io_r_1_cluster_49_addr(sram_cluster_0_io_r_1_cluster_49_addr),
    .io_r_1_cluster_49_data(sram_cluster_0_io_r_1_cluster_49_data),
    .io_r_1_cluster_50_en(sram_cluster_0_io_r_1_cluster_50_en),
    .io_r_1_cluster_50_addr(sram_cluster_0_io_r_1_cluster_50_addr),
    .io_r_1_cluster_50_data(sram_cluster_0_io_r_1_cluster_50_data),
    .io_r_1_cluster_51_en(sram_cluster_0_io_r_1_cluster_51_en),
    .io_r_1_cluster_51_addr(sram_cluster_0_io_r_1_cluster_51_addr),
    .io_r_1_cluster_51_data(sram_cluster_0_io_r_1_cluster_51_data),
    .io_r_1_cluster_52_en(sram_cluster_0_io_r_1_cluster_52_en),
    .io_r_1_cluster_52_addr(sram_cluster_0_io_r_1_cluster_52_addr),
    .io_r_1_cluster_52_data(sram_cluster_0_io_r_1_cluster_52_data),
    .io_r_1_cluster_53_en(sram_cluster_0_io_r_1_cluster_53_en),
    .io_r_1_cluster_53_addr(sram_cluster_0_io_r_1_cluster_53_addr),
    .io_r_1_cluster_53_data(sram_cluster_0_io_r_1_cluster_53_data),
    .io_r_1_cluster_54_en(sram_cluster_0_io_r_1_cluster_54_en),
    .io_r_1_cluster_54_addr(sram_cluster_0_io_r_1_cluster_54_addr),
    .io_r_1_cluster_54_data(sram_cluster_0_io_r_1_cluster_54_data),
    .io_r_1_cluster_55_en(sram_cluster_0_io_r_1_cluster_55_en),
    .io_r_1_cluster_55_addr(sram_cluster_0_io_r_1_cluster_55_addr),
    .io_r_1_cluster_55_data(sram_cluster_0_io_r_1_cluster_55_data),
    .io_r_1_cluster_56_en(sram_cluster_0_io_r_1_cluster_56_en),
    .io_r_1_cluster_56_addr(sram_cluster_0_io_r_1_cluster_56_addr),
    .io_r_1_cluster_56_data(sram_cluster_0_io_r_1_cluster_56_data),
    .io_r_1_cluster_57_en(sram_cluster_0_io_r_1_cluster_57_en),
    .io_r_1_cluster_57_addr(sram_cluster_0_io_r_1_cluster_57_addr),
    .io_r_1_cluster_57_data(sram_cluster_0_io_r_1_cluster_57_data),
    .io_r_1_cluster_58_en(sram_cluster_0_io_r_1_cluster_58_en),
    .io_r_1_cluster_58_addr(sram_cluster_0_io_r_1_cluster_58_addr),
    .io_r_1_cluster_58_data(sram_cluster_0_io_r_1_cluster_58_data),
    .io_r_1_cluster_59_en(sram_cluster_0_io_r_1_cluster_59_en),
    .io_r_1_cluster_59_addr(sram_cluster_0_io_r_1_cluster_59_addr),
    .io_r_1_cluster_59_data(sram_cluster_0_io_r_1_cluster_59_data),
    .io_r_1_cluster_60_en(sram_cluster_0_io_r_1_cluster_60_en),
    .io_r_1_cluster_60_addr(sram_cluster_0_io_r_1_cluster_60_addr),
    .io_r_1_cluster_60_data(sram_cluster_0_io_r_1_cluster_60_data),
    .io_r_1_cluster_61_en(sram_cluster_0_io_r_1_cluster_61_en),
    .io_r_1_cluster_61_addr(sram_cluster_0_io_r_1_cluster_61_addr),
    .io_r_1_cluster_61_data(sram_cluster_0_io_r_1_cluster_61_data),
    .io_r_1_cluster_62_en(sram_cluster_0_io_r_1_cluster_62_en),
    .io_r_1_cluster_62_addr(sram_cluster_0_io_r_1_cluster_62_addr),
    .io_r_1_cluster_62_data(sram_cluster_0_io_r_1_cluster_62_data),
    .io_r_1_cluster_63_en(sram_cluster_0_io_r_1_cluster_63_en),
    .io_r_1_cluster_63_addr(sram_cluster_0_io_r_1_cluster_63_addr),
    .io_r_1_cluster_63_data(sram_cluster_0_io_r_1_cluster_63_data),
    .io_r_2_cluster_0_en(sram_cluster_0_io_r_2_cluster_0_en),
    .io_r_2_cluster_0_addr(sram_cluster_0_io_r_2_cluster_0_addr),
    .io_r_2_cluster_0_data(sram_cluster_0_io_r_2_cluster_0_data),
    .io_r_2_cluster_1_en(sram_cluster_0_io_r_2_cluster_1_en),
    .io_r_2_cluster_1_addr(sram_cluster_0_io_r_2_cluster_1_addr),
    .io_r_2_cluster_1_data(sram_cluster_0_io_r_2_cluster_1_data),
    .io_r_2_cluster_2_en(sram_cluster_0_io_r_2_cluster_2_en),
    .io_r_2_cluster_2_addr(sram_cluster_0_io_r_2_cluster_2_addr),
    .io_r_2_cluster_2_data(sram_cluster_0_io_r_2_cluster_2_data),
    .io_r_2_cluster_3_en(sram_cluster_0_io_r_2_cluster_3_en),
    .io_r_2_cluster_3_addr(sram_cluster_0_io_r_2_cluster_3_addr),
    .io_r_2_cluster_3_data(sram_cluster_0_io_r_2_cluster_3_data),
    .io_r_2_cluster_4_en(sram_cluster_0_io_r_2_cluster_4_en),
    .io_r_2_cluster_4_addr(sram_cluster_0_io_r_2_cluster_4_addr),
    .io_r_2_cluster_4_data(sram_cluster_0_io_r_2_cluster_4_data),
    .io_r_2_cluster_5_en(sram_cluster_0_io_r_2_cluster_5_en),
    .io_r_2_cluster_5_addr(sram_cluster_0_io_r_2_cluster_5_addr),
    .io_r_2_cluster_5_data(sram_cluster_0_io_r_2_cluster_5_data),
    .io_r_2_cluster_6_en(sram_cluster_0_io_r_2_cluster_6_en),
    .io_r_2_cluster_6_addr(sram_cluster_0_io_r_2_cluster_6_addr),
    .io_r_2_cluster_6_data(sram_cluster_0_io_r_2_cluster_6_data),
    .io_r_2_cluster_7_en(sram_cluster_0_io_r_2_cluster_7_en),
    .io_r_2_cluster_7_addr(sram_cluster_0_io_r_2_cluster_7_addr),
    .io_r_2_cluster_7_data(sram_cluster_0_io_r_2_cluster_7_data),
    .io_r_2_cluster_8_en(sram_cluster_0_io_r_2_cluster_8_en),
    .io_r_2_cluster_8_addr(sram_cluster_0_io_r_2_cluster_8_addr),
    .io_r_2_cluster_8_data(sram_cluster_0_io_r_2_cluster_8_data),
    .io_r_2_cluster_9_en(sram_cluster_0_io_r_2_cluster_9_en),
    .io_r_2_cluster_9_addr(sram_cluster_0_io_r_2_cluster_9_addr),
    .io_r_2_cluster_9_data(sram_cluster_0_io_r_2_cluster_9_data),
    .io_r_2_cluster_10_en(sram_cluster_0_io_r_2_cluster_10_en),
    .io_r_2_cluster_10_addr(sram_cluster_0_io_r_2_cluster_10_addr),
    .io_r_2_cluster_10_data(sram_cluster_0_io_r_2_cluster_10_data),
    .io_r_2_cluster_11_en(sram_cluster_0_io_r_2_cluster_11_en),
    .io_r_2_cluster_11_addr(sram_cluster_0_io_r_2_cluster_11_addr),
    .io_r_2_cluster_11_data(sram_cluster_0_io_r_2_cluster_11_data),
    .io_r_2_cluster_12_en(sram_cluster_0_io_r_2_cluster_12_en),
    .io_r_2_cluster_12_addr(sram_cluster_0_io_r_2_cluster_12_addr),
    .io_r_2_cluster_12_data(sram_cluster_0_io_r_2_cluster_12_data),
    .io_r_2_cluster_13_en(sram_cluster_0_io_r_2_cluster_13_en),
    .io_r_2_cluster_13_addr(sram_cluster_0_io_r_2_cluster_13_addr),
    .io_r_2_cluster_13_data(sram_cluster_0_io_r_2_cluster_13_data),
    .io_r_2_cluster_14_en(sram_cluster_0_io_r_2_cluster_14_en),
    .io_r_2_cluster_14_addr(sram_cluster_0_io_r_2_cluster_14_addr),
    .io_r_2_cluster_14_data(sram_cluster_0_io_r_2_cluster_14_data),
    .io_r_2_cluster_15_en(sram_cluster_0_io_r_2_cluster_15_en),
    .io_r_2_cluster_15_addr(sram_cluster_0_io_r_2_cluster_15_addr),
    .io_r_2_cluster_15_data(sram_cluster_0_io_r_2_cluster_15_data),
    .io_r_2_cluster_16_en(sram_cluster_0_io_r_2_cluster_16_en),
    .io_r_2_cluster_16_addr(sram_cluster_0_io_r_2_cluster_16_addr),
    .io_r_2_cluster_16_data(sram_cluster_0_io_r_2_cluster_16_data),
    .io_r_2_cluster_17_en(sram_cluster_0_io_r_2_cluster_17_en),
    .io_r_2_cluster_17_addr(sram_cluster_0_io_r_2_cluster_17_addr),
    .io_r_2_cluster_17_data(sram_cluster_0_io_r_2_cluster_17_data),
    .io_r_2_cluster_18_en(sram_cluster_0_io_r_2_cluster_18_en),
    .io_r_2_cluster_18_addr(sram_cluster_0_io_r_2_cluster_18_addr),
    .io_r_2_cluster_18_data(sram_cluster_0_io_r_2_cluster_18_data),
    .io_r_2_cluster_19_en(sram_cluster_0_io_r_2_cluster_19_en),
    .io_r_2_cluster_19_addr(sram_cluster_0_io_r_2_cluster_19_addr),
    .io_r_2_cluster_19_data(sram_cluster_0_io_r_2_cluster_19_data),
    .io_r_2_cluster_20_en(sram_cluster_0_io_r_2_cluster_20_en),
    .io_r_2_cluster_20_addr(sram_cluster_0_io_r_2_cluster_20_addr),
    .io_r_2_cluster_20_data(sram_cluster_0_io_r_2_cluster_20_data),
    .io_r_2_cluster_21_en(sram_cluster_0_io_r_2_cluster_21_en),
    .io_r_2_cluster_21_addr(sram_cluster_0_io_r_2_cluster_21_addr),
    .io_r_2_cluster_21_data(sram_cluster_0_io_r_2_cluster_21_data),
    .io_r_2_cluster_22_en(sram_cluster_0_io_r_2_cluster_22_en),
    .io_r_2_cluster_22_addr(sram_cluster_0_io_r_2_cluster_22_addr),
    .io_r_2_cluster_22_data(sram_cluster_0_io_r_2_cluster_22_data),
    .io_r_2_cluster_23_en(sram_cluster_0_io_r_2_cluster_23_en),
    .io_r_2_cluster_23_addr(sram_cluster_0_io_r_2_cluster_23_addr),
    .io_r_2_cluster_23_data(sram_cluster_0_io_r_2_cluster_23_data),
    .io_r_2_cluster_24_en(sram_cluster_0_io_r_2_cluster_24_en),
    .io_r_2_cluster_24_addr(sram_cluster_0_io_r_2_cluster_24_addr),
    .io_r_2_cluster_24_data(sram_cluster_0_io_r_2_cluster_24_data),
    .io_r_2_cluster_25_en(sram_cluster_0_io_r_2_cluster_25_en),
    .io_r_2_cluster_25_addr(sram_cluster_0_io_r_2_cluster_25_addr),
    .io_r_2_cluster_25_data(sram_cluster_0_io_r_2_cluster_25_data),
    .io_r_2_cluster_26_en(sram_cluster_0_io_r_2_cluster_26_en),
    .io_r_2_cluster_26_addr(sram_cluster_0_io_r_2_cluster_26_addr),
    .io_r_2_cluster_26_data(sram_cluster_0_io_r_2_cluster_26_data),
    .io_r_2_cluster_27_en(sram_cluster_0_io_r_2_cluster_27_en),
    .io_r_2_cluster_27_addr(sram_cluster_0_io_r_2_cluster_27_addr),
    .io_r_2_cluster_27_data(sram_cluster_0_io_r_2_cluster_27_data),
    .io_r_2_cluster_28_en(sram_cluster_0_io_r_2_cluster_28_en),
    .io_r_2_cluster_28_addr(sram_cluster_0_io_r_2_cluster_28_addr),
    .io_r_2_cluster_28_data(sram_cluster_0_io_r_2_cluster_28_data),
    .io_r_2_cluster_29_en(sram_cluster_0_io_r_2_cluster_29_en),
    .io_r_2_cluster_29_addr(sram_cluster_0_io_r_2_cluster_29_addr),
    .io_r_2_cluster_29_data(sram_cluster_0_io_r_2_cluster_29_data),
    .io_r_2_cluster_30_en(sram_cluster_0_io_r_2_cluster_30_en),
    .io_r_2_cluster_30_addr(sram_cluster_0_io_r_2_cluster_30_addr),
    .io_r_2_cluster_30_data(sram_cluster_0_io_r_2_cluster_30_data),
    .io_r_2_cluster_31_en(sram_cluster_0_io_r_2_cluster_31_en),
    .io_r_2_cluster_31_addr(sram_cluster_0_io_r_2_cluster_31_addr),
    .io_r_2_cluster_31_data(sram_cluster_0_io_r_2_cluster_31_data),
    .io_r_2_cluster_32_en(sram_cluster_0_io_r_2_cluster_32_en),
    .io_r_2_cluster_32_addr(sram_cluster_0_io_r_2_cluster_32_addr),
    .io_r_2_cluster_32_data(sram_cluster_0_io_r_2_cluster_32_data),
    .io_r_2_cluster_33_en(sram_cluster_0_io_r_2_cluster_33_en),
    .io_r_2_cluster_33_addr(sram_cluster_0_io_r_2_cluster_33_addr),
    .io_r_2_cluster_33_data(sram_cluster_0_io_r_2_cluster_33_data),
    .io_r_2_cluster_34_en(sram_cluster_0_io_r_2_cluster_34_en),
    .io_r_2_cluster_34_addr(sram_cluster_0_io_r_2_cluster_34_addr),
    .io_r_2_cluster_34_data(sram_cluster_0_io_r_2_cluster_34_data),
    .io_r_2_cluster_35_en(sram_cluster_0_io_r_2_cluster_35_en),
    .io_r_2_cluster_35_addr(sram_cluster_0_io_r_2_cluster_35_addr),
    .io_r_2_cluster_35_data(sram_cluster_0_io_r_2_cluster_35_data),
    .io_r_2_cluster_36_en(sram_cluster_0_io_r_2_cluster_36_en),
    .io_r_2_cluster_36_addr(sram_cluster_0_io_r_2_cluster_36_addr),
    .io_r_2_cluster_36_data(sram_cluster_0_io_r_2_cluster_36_data),
    .io_r_2_cluster_37_en(sram_cluster_0_io_r_2_cluster_37_en),
    .io_r_2_cluster_37_addr(sram_cluster_0_io_r_2_cluster_37_addr),
    .io_r_2_cluster_37_data(sram_cluster_0_io_r_2_cluster_37_data),
    .io_r_2_cluster_38_en(sram_cluster_0_io_r_2_cluster_38_en),
    .io_r_2_cluster_38_addr(sram_cluster_0_io_r_2_cluster_38_addr),
    .io_r_2_cluster_38_data(sram_cluster_0_io_r_2_cluster_38_data),
    .io_r_2_cluster_39_en(sram_cluster_0_io_r_2_cluster_39_en),
    .io_r_2_cluster_39_addr(sram_cluster_0_io_r_2_cluster_39_addr),
    .io_r_2_cluster_39_data(sram_cluster_0_io_r_2_cluster_39_data),
    .io_r_2_cluster_40_en(sram_cluster_0_io_r_2_cluster_40_en),
    .io_r_2_cluster_40_addr(sram_cluster_0_io_r_2_cluster_40_addr),
    .io_r_2_cluster_40_data(sram_cluster_0_io_r_2_cluster_40_data),
    .io_r_2_cluster_41_en(sram_cluster_0_io_r_2_cluster_41_en),
    .io_r_2_cluster_41_addr(sram_cluster_0_io_r_2_cluster_41_addr),
    .io_r_2_cluster_41_data(sram_cluster_0_io_r_2_cluster_41_data),
    .io_r_2_cluster_42_en(sram_cluster_0_io_r_2_cluster_42_en),
    .io_r_2_cluster_42_addr(sram_cluster_0_io_r_2_cluster_42_addr),
    .io_r_2_cluster_42_data(sram_cluster_0_io_r_2_cluster_42_data),
    .io_r_2_cluster_43_en(sram_cluster_0_io_r_2_cluster_43_en),
    .io_r_2_cluster_43_addr(sram_cluster_0_io_r_2_cluster_43_addr),
    .io_r_2_cluster_43_data(sram_cluster_0_io_r_2_cluster_43_data),
    .io_r_2_cluster_44_en(sram_cluster_0_io_r_2_cluster_44_en),
    .io_r_2_cluster_44_addr(sram_cluster_0_io_r_2_cluster_44_addr),
    .io_r_2_cluster_44_data(sram_cluster_0_io_r_2_cluster_44_data),
    .io_r_2_cluster_45_en(sram_cluster_0_io_r_2_cluster_45_en),
    .io_r_2_cluster_45_addr(sram_cluster_0_io_r_2_cluster_45_addr),
    .io_r_2_cluster_45_data(sram_cluster_0_io_r_2_cluster_45_data),
    .io_r_2_cluster_46_en(sram_cluster_0_io_r_2_cluster_46_en),
    .io_r_2_cluster_46_addr(sram_cluster_0_io_r_2_cluster_46_addr),
    .io_r_2_cluster_46_data(sram_cluster_0_io_r_2_cluster_46_data),
    .io_r_2_cluster_47_en(sram_cluster_0_io_r_2_cluster_47_en),
    .io_r_2_cluster_47_addr(sram_cluster_0_io_r_2_cluster_47_addr),
    .io_r_2_cluster_47_data(sram_cluster_0_io_r_2_cluster_47_data),
    .io_r_2_cluster_48_en(sram_cluster_0_io_r_2_cluster_48_en),
    .io_r_2_cluster_48_addr(sram_cluster_0_io_r_2_cluster_48_addr),
    .io_r_2_cluster_48_data(sram_cluster_0_io_r_2_cluster_48_data),
    .io_r_2_cluster_49_en(sram_cluster_0_io_r_2_cluster_49_en),
    .io_r_2_cluster_49_addr(sram_cluster_0_io_r_2_cluster_49_addr),
    .io_r_2_cluster_49_data(sram_cluster_0_io_r_2_cluster_49_data),
    .io_r_2_cluster_50_en(sram_cluster_0_io_r_2_cluster_50_en),
    .io_r_2_cluster_50_addr(sram_cluster_0_io_r_2_cluster_50_addr),
    .io_r_2_cluster_50_data(sram_cluster_0_io_r_2_cluster_50_data),
    .io_r_2_cluster_51_en(sram_cluster_0_io_r_2_cluster_51_en),
    .io_r_2_cluster_51_addr(sram_cluster_0_io_r_2_cluster_51_addr),
    .io_r_2_cluster_51_data(sram_cluster_0_io_r_2_cluster_51_data),
    .io_r_2_cluster_52_en(sram_cluster_0_io_r_2_cluster_52_en),
    .io_r_2_cluster_52_addr(sram_cluster_0_io_r_2_cluster_52_addr),
    .io_r_2_cluster_52_data(sram_cluster_0_io_r_2_cluster_52_data),
    .io_r_2_cluster_53_en(sram_cluster_0_io_r_2_cluster_53_en),
    .io_r_2_cluster_53_addr(sram_cluster_0_io_r_2_cluster_53_addr),
    .io_r_2_cluster_53_data(sram_cluster_0_io_r_2_cluster_53_data),
    .io_r_2_cluster_54_en(sram_cluster_0_io_r_2_cluster_54_en),
    .io_r_2_cluster_54_addr(sram_cluster_0_io_r_2_cluster_54_addr),
    .io_r_2_cluster_54_data(sram_cluster_0_io_r_2_cluster_54_data),
    .io_r_2_cluster_55_en(sram_cluster_0_io_r_2_cluster_55_en),
    .io_r_2_cluster_55_addr(sram_cluster_0_io_r_2_cluster_55_addr),
    .io_r_2_cluster_55_data(sram_cluster_0_io_r_2_cluster_55_data),
    .io_r_2_cluster_56_en(sram_cluster_0_io_r_2_cluster_56_en),
    .io_r_2_cluster_56_addr(sram_cluster_0_io_r_2_cluster_56_addr),
    .io_r_2_cluster_56_data(sram_cluster_0_io_r_2_cluster_56_data),
    .io_r_2_cluster_57_en(sram_cluster_0_io_r_2_cluster_57_en),
    .io_r_2_cluster_57_addr(sram_cluster_0_io_r_2_cluster_57_addr),
    .io_r_2_cluster_57_data(sram_cluster_0_io_r_2_cluster_57_data),
    .io_r_2_cluster_58_en(sram_cluster_0_io_r_2_cluster_58_en),
    .io_r_2_cluster_58_addr(sram_cluster_0_io_r_2_cluster_58_addr),
    .io_r_2_cluster_58_data(sram_cluster_0_io_r_2_cluster_58_data),
    .io_r_2_cluster_59_en(sram_cluster_0_io_r_2_cluster_59_en),
    .io_r_2_cluster_59_addr(sram_cluster_0_io_r_2_cluster_59_addr),
    .io_r_2_cluster_59_data(sram_cluster_0_io_r_2_cluster_59_data),
    .io_r_2_cluster_60_en(sram_cluster_0_io_r_2_cluster_60_en),
    .io_r_2_cluster_60_addr(sram_cluster_0_io_r_2_cluster_60_addr),
    .io_r_2_cluster_60_data(sram_cluster_0_io_r_2_cluster_60_data),
    .io_r_2_cluster_61_en(sram_cluster_0_io_r_2_cluster_61_en),
    .io_r_2_cluster_61_addr(sram_cluster_0_io_r_2_cluster_61_addr),
    .io_r_2_cluster_61_data(sram_cluster_0_io_r_2_cluster_61_data),
    .io_r_2_cluster_62_en(sram_cluster_0_io_r_2_cluster_62_en),
    .io_r_2_cluster_62_addr(sram_cluster_0_io_r_2_cluster_62_addr),
    .io_r_2_cluster_62_data(sram_cluster_0_io_r_2_cluster_62_data),
    .io_r_2_cluster_63_en(sram_cluster_0_io_r_2_cluster_63_en),
    .io_r_2_cluster_63_addr(sram_cluster_0_io_r_2_cluster_63_addr),
    .io_r_2_cluster_63_data(sram_cluster_0_io_r_2_cluster_63_data),
    .io_r_3_cluster_0_en(sram_cluster_0_io_r_3_cluster_0_en),
    .io_r_3_cluster_0_addr(sram_cluster_0_io_r_3_cluster_0_addr),
    .io_r_3_cluster_0_data(sram_cluster_0_io_r_3_cluster_0_data),
    .io_r_3_cluster_1_en(sram_cluster_0_io_r_3_cluster_1_en),
    .io_r_3_cluster_1_addr(sram_cluster_0_io_r_3_cluster_1_addr),
    .io_r_3_cluster_1_data(sram_cluster_0_io_r_3_cluster_1_data),
    .io_r_3_cluster_2_en(sram_cluster_0_io_r_3_cluster_2_en),
    .io_r_3_cluster_2_addr(sram_cluster_0_io_r_3_cluster_2_addr),
    .io_r_3_cluster_2_data(sram_cluster_0_io_r_3_cluster_2_data),
    .io_r_3_cluster_3_en(sram_cluster_0_io_r_3_cluster_3_en),
    .io_r_3_cluster_3_addr(sram_cluster_0_io_r_3_cluster_3_addr),
    .io_r_3_cluster_3_data(sram_cluster_0_io_r_3_cluster_3_data),
    .io_r_3_cluster_4_en(sram_cluster_0_io_r_3_cluster_4_en),
    .io_r_3_cluster_4_addr(sram_cluster_0_io_r_3_cluster_4_addr),
    .io_r_3_cluster_4_data(sram_cluster_0_io_r_3_cluster_4_data),
    .io_r_3_cluster_5_en(sram_cluster_0_io_r_3_cluster_5_en),
    .io_r_3_cluster_5_addr(sram_cluster_0_io_r_3_cluster_5_addr),
    .io_r_3_cluster_5_data(sram_cluster_0_io_r_3_cluster_5_data),
    .io_r_3_cluster_6_en(sram_cluster_0_io_r_3_cluster_6_en),
    .io_r_3_cluster_6_addr(sram_cluster_0_io_r_3_cluster_6_addr),
    .io_r_3_cluster_6_data(sram_cluster_0_io_r_3_cluster_6_data),
    .io_r_3_cluster_7_en(sram_cluster_0_io_r_3_cluster_7_en),
    .io_r_3_cluster_7_addr(sram_cluster_0_io_r_3_cluster_7_addr),
    .io_r_3_cluster_7_data(sram_cluster_0_io_r_3_cluster_7_data),
    .io_r_3_cluster_8_en(sram_cluster_0_io_r_3_cluster_8_en),
    .io_r_3_cluster_8_addr(sram_cluster_0_io_r_3_cluster_8_addr),
    .io_r_3_cluster_8_data(sram_cluster_0_io_r_3_cluster_8_data),
    .io_r_3_cluster_9_en(sram_cluster_0_io_r_3_cluster_9_en),
    .io_r_3_cluster_9_addr(sram_cluster_0_io_r_3_cluster_9_addr),
    .io_r_3_cluster_9_data(sram_cluster_0_io_r_3_cluster_9_data),
    .io_r_3_cluster_10_en(sram_cluster_0_io_r_3_cluster_10_en),
    .io_r_3_cluster_10_addr(sram_cluster_0_io_r_3_cluster_10_addr),
    .io_r_3_cluster_10_data(sram_cluster_0_io_r_3_cluster_10_data),
    .io_r_3_cluster_11_en(sram_cluster_0_io_r_3_cluster_11_en),
    .io_r_3_cluster_11_addr(sram_cluster_0_io_r_3_cluster_11_addr),
    .io_r_3_cluster_11_data(sram_cluster_0_io_r_3_cluster_11_data),
    .io_r_3_cluster_12_en(sram_cluster_0_io_r_3_cluster_12_en),
    .io_r_3_cluster_12_addr(sram_cluster_0_io_r_3_cluster_12_addr),
    .io_r_3_cluster_12_data(sram_cluster_0_io_r_3_cluster_12_data),
    .io_r_3_cluster_13_en(sram_cluster_0_io_r_3_cluster_13_en),
    .io_r_3_cluster_13_addr(sram_cluster_0_io_r_3_cluster_13_addr),
    .io_r_3_cluster_13_data(sram_cluster_0_io_r_3_cluster_13_data),
    .io_r_3_cluster_14_en(sram_cluster_0_io_r_3_cluster_14_en),
    .io_r_3_cluster_14_addr(sram_cluster_0_io_r_3_cluster_14_addr),
    .io_r_3_cluster_14_data(sram_cluster_0_io_r_3_cluster_14_data),
    .io_r_3_cluster_15_en(sram_cluster_0_io_r_3_cluster_15_en),
    .io_r_3_cluster_15_addr(sram_cluster_0_io_r_3_cluster_15_addr),
    .io_r_3_cluster_15_data(sram_cluster_0_io_r_3_cluster_15_data),
    .io_r_3_cluster_16_en(sram_cluster_0_io_r_3_cluster_16_en),
    .io_r_3_cluster_16_addr(sram_cluster_0_io_r_3_cluster_16_addr),
    .io_r_3_cluster_16_data(sram_cluster_0_io_r_3_cluster_16_data),
    .io_r_3_cluster_17_en(sram_cluster_0_io_r_3_cluster_17_en),
    .io_r_3_cluster_17_addr(sram_cluster_0_io_r_3_cluster_17_addr),
    .io_r_3_cluster_17_data(sram_cluster_0_io_r_3_cluster_17_data),
    .io_r_3_cluster_18_en(sram_cluster_0_io_r_3_cluster_18_en),
    .io_r_3_cluster_18_addr(sram_cluster_0_io_r_3_cluster_18_addr),
    .io_r_3_cluster_18_data(sram_cluster_0_io_r_3_cluster_18_data),
    .io_r_3_cluster_19_en(sram_cluster_0_io_r_3_cluster_19_en),
    .io_r_3_cluster_19_addr(sram_cluster_0_io_r_3_cluster_19_addr),
    .io_r_3_cluster_19_data(sram_cluster_0_io_r_3_cluster_19_data),
    .io_r_3_cluster_20_en(sram_cluster_0_io_r_3_cluster_20_en),
    .io_r_3_cluster_20_addr(sram_cluster_0_io_r_3_cluster_20_addr),
    .io_r_3_cluster_20_data(sram_cluster_0_io_r_3_cluster_20_data),
    .io_r_3_cluster_21_en(sram_cluster_0_io_r_3_cluster_21_en),
    .io_r_3_cluster_21_addr(sram_cluster_0_io_r_3_cluster_21_addr),
    .io_r_3_cluster_21_data(sram_cluster_0_io_r_3_cluster_21_data),
    .io_r_3_cluster_22_en(sram_cluster_0_io_r_3_cluster_22_en),
    .io_r_3_cluster_22_addr(sram_cluster_0_io_r_3_cluster_22_addr),
    .io_r_3_cluster_22_data(sram_cluster_0_io_r_3_cluster_22_data),
    .io_r_3_cluster_23_en(sram_cluster_0_io_r_3_cluster_23_en),
    .io_r_3_cluster_23_addr(sram_cluster_0_io_r_3_cluster_23_addr),
    .io_r_3_cluster_23_data(sram_cluster_0_io_r_3_cluster_23_data),
    .io_r_3_cluster_24_en(sram_cluster_0_io_r_3_cluster_24_en),
    .io_r_3_cluster_24_addr(sram_cluster_0_io_r_3_cluster_24_addr),
    .io_r_3_cluster_24_data(sram_cluster_0_io_r_3_cluster_24_data),
    .io_r_3_cluster_25_en(sram_cluster_0_io_r_3_cluster_25_en),
    .io_r_3_cluster_25_addr(sram_cluster_0_io_r_3_cluster_25_addr),
    .io_r_3_cluster_25_data(sram_cluster_0_io_r_3_cluster_25_data),
    .io_r_3_cluster_26_en(sram_cluster_0_io_r_3_cluster_26_en),
    .io_r_3_cluster_26_addr(sram_cluster_0_io_r_3_cluster_26_addr),
    .io_r_3_cluster_26_data(sram_cluster_0_io_r_3_cluster_26_data),
    .io_r_3_cluster_27_en(sram_cluster_0_io_r_3_cluster_27_en),
    .io_r_3_cluster_27_addr(sram_cluster_0_io_r_3_cluster_27_addr),
    .io_r_3_cluster_27_data(sram_cluster_0_io_r_3_cluster_27_data),
    .io_r_3_cluster_28_en(sram_cluster_0_io_r_3_cluster_28_en),
    .io_r_3_cluster_28_addr(sram_cluster_0_io_r_3_cluster_28_addr),
    .io_r_3_cluster_28_data(sram_cluster_0_io_r_3_cluster_28_data),
    .io_r_3_cluster_29_en(sram_cluster_0_io_r_3_cluster_29_en),
    .io_r_3_cluster_29_addr(sram_cluster_0_io_r_3_cluster_29_addr),
    .io_r_3_cluster_29_data(sram_cluster_0_io_r_3_cluster_29_data),
    .io_r_3_cluster_30_en(sram_cluster_0_io_r_3_cluster_30_en),
    .io_r_3_cluster_30_addr(sram_cluster_0_io_r_3_cluster_30_addr),
    .io_r_3_cluster_30_data(sram_cluster_0_io_r_3_cluster_30_data),
    .io_r_3_cluster_31_en(sram_cluster_0_io_r_3_cluster_31_en),
    .io_r_3_cluster_31_addr(sram_cluster_0_io_r_3_cluster_31_addr),
    .io_r_3_cluster_31_data(sram_cluster_0_io_r_3_cluster_31_data),
    .io_r_3_cluster_32_en(sram_cluster_0_io_r_3_cluster_32_en),
    .io_r_3_cluster_32_addr(sram_cluster_0_io_r_3_cluster_32_addr),
    .io_r_3_cluster_32_data(sram_cluster_0_io_r_3_cluster_32_data),
    .io_r_3_cluster_33_en(sram_cluster_0_io_r_3_cluster_33_en),
    .io_r_3_cluster_33_addr(sram_cluster_0_io_r_3_cluster_33_addr),
    .io_r_3_cluster_33_data(sram_cluster_0_io_r_3_cluster_33_data),
    .io_r_3_cluster_34_en(sram_cluster_0_io_r_3_cluster_34_en),
    .io_r_3_cluster_34_addr(sram_cluster_0_io_r_3_cluster_34_addr),
    .io_r_3_cluster_34_data(sram_cluster_0_io_r_3_cluster_34_data),
    .io_r_3_cluster_35_en(sram_cluster_0_io_r_3_cluster_35_en),
    .io_r_3_cluster_35_addr(sram_cluster_0_io_r_3_cluster_35_addr),
    .io_r_3_cluster_35_data(sram_cluster_0_io_r_3_cluster_35_data),
    .io_r_3_cluster_36_en(sram_cluster_0_io_r_3_cluster_36_en),
    .io_r_3_cluster_36_addr(sram_cluster_0_io_r_3_cluster_36_addr),
    .io_r_3_cluster_36_data(sram_cluster_0_io_r_3_cluster_36_data),
    .io_r_3_cluster_37_en(sram_cluster_0_io_r_3_cluster_37_en),
    .io_r_3_cluster_37_addr(sram_cluster_0_io_r_3_cluster_37_addr),
    .io_r_3_cluster_37_data(sram_cluster_0_io_r_3_cluster_37_data),
    .io_r_3_cluster_38_en(sram_cluster_0_io_r_3_cluster_38_en),
    .io_r_3_cluster_38_addr(sram_cluster_0_io_r_3_cluster_38_addr),
    .io_r_3_cluster_38_data(sram_cluster_0_io_r_3_cluster_38_data),
    .io_r_3_cluster_39_en(sram_cluster_0_io_r_3_cluster_39_en),
    .io_r_3_cluster_39_addr(sram_cluster_0_io_r_3_cluster_39_addr),
    .io_r_3_cluster_39_data(sram_cluster_0_io_r_3_cluster_39_data),
    .io_r_3_cluster_40_en(sram_cluster_0_io_r_3_cluster_40_en),
    .io_r_3_cluster_40_addr(sram_cluster_0_io_r_3_cluster_40_addr),
    .io_r_3_cluster_40_data(sram_cluster_0_io_r_3_cluster_40_data),
    .io_r_3_cluster_41_en(sram_cluster_0_io_r_3_cluster_41_en),
    .io_r_3_cluster_41_addr(sram_cluster_0_io_r_3_cluster_41_addr),
    .io_r_3_cluster_41_data(sram_cluster_0_io_r_3_cluster_41_data),
    .io_r_3_cluster_42_en(sram_cluster_0_io_r_3_cluster_42_en),
    .io_r_3_cluster_42_addr(sram_cluster_0_io_r_3_cluster_42_addr),
    .io_r_3_cluster_42_data(sram_cluster_0_io_r_3_cluster_42_data),
    .io_r_3_cluster_43_en(sram_cluster_0_io_r_3_cluster_43_en),
    .io_r_3_cluster_43_addr(sram_cluster_0_io_r_3_cluster_43_addr),
    .io_r_3_cluster_43_data(sram_cluster_0_io_r_3_cluster_43_data),
    .io_r_3_cluster_44_en(sram_cluster_0_io_r_3_cluster_44_en),
    .io_r_3_cluster_44_addr(sram_cluster_0_io_r_3_cluster_44_addr),
    .io_r_3_cluster_44_data(sram_cluster_0_io_r_3_cluster_44_data),
    .io_r_3_cluster_45_en(sram_cluster_0_io_r_3_cluster_45_en),
    .io_r_3_cluster_45_addr(sram_cluster_0_io_r_3_cluster_45_addr),
    .io_r_3_cluster_45_data(sram_cluster_0_io_r_3_cluster_45_data),
    .io_r_3_cluster_46_en(sram_cluster_0_io_r_3_cluster_46_en),
    .io_r_3_cluster_46_addr(sram_cluster_0_io_r_3_cluster_46_addr),
    .io_r_3_cluster_46_data(sram_cluster_0_io_r_3_cluster_46_data),
    .io_r_3_cluster_47_en(sram_cluster_0_io_r_3_cluster_47_en),
    .io_r_3_cluster_47_addr(sram_cluster_0_io_r_3_cluster_47_addr),
    .io_r_3_cluster_47_data(sram_cluster_0_io_r_3_cluster_47_data),
    .io_r_3_cluster_48_en(sram_cluster_0_io_r_3_cluster_48_en),
    .io_r_3_cluster_48_addr(sram_cluster_0_io_r_3_cluster_48_addr),
    .io_r_3_cluster_48_data(sram_cluster_0_io_r_3_cluster_48_data),
    .io_r_3_cluster_49_en(sram_cluster_0_io_r_3_cluster_49_en),
    .io_r_3_cluster_49_addr(sram_cluster_0_io_r_3_cluster_49_addr),
    .io_r_3_cluster_49_data(sram_cluster_0_io_r_3_cluster_49_data),
    .io_r_3_cluster_50_en(sram_cluster_0_io_r_3_cluster_50_en),
    .io_r_3_cluster_50_addr(sram_cluster_0_io_r_3_cluster_50_addr),
    .io_r_3_cluster_50_data(sram_cluster_0_io_r_3_cluster_50_data),
    .io_r_3_cluster_51_en(sram_cluster_0_io_r_3_cluster_51_en),
    .io_r_3_cluster_51_addr(sram_cluster_0_io_r_3_cluster_51_addr),
    .io_r_3_cluster_51_data(sram_cluster_0_io_r_3_cluster_51_data),
    .io_r_3_cluster_52_en(sram_cluster_0_io_r_3_cluster_52_en),
    .io_r_3_cluster_52_addr(sram_cluster_0_io_r_3_cluster_52_addr),
    .io_r_3_cluster_52_data(sram_cluster_0_io_r_3_cluster_52_data),
    .io_r_3_cluster_53_en(sram_cluster_0_io_r_3_cluster_53_en),
    .io_r_3_cluster_53_addr(sram_cluster_0_io_r_3_cluster_53_addr),
    .io_r_3_cluster_53_data(sram_cluster_0_io_r_3_cluster_53_data),
    .io_r_3_cluster_54_en(sram_cluster_0_io_r_3_cluster_54_en),
    .io_r_3_cluster_54_addr(sram_cluster_0_io_r_3_cluster_54_addr),
    .io_r_3_cluster_54_data(sram_cluster_0_io_r_3_cluster_54_data),
    .io_r_3_cluster_55_en(sram_cluster_0_io_r_3_cluster_55_en),
    .io_r_3_cluster_55_addr(sram_cluster_0_io_r_3_cluster_55_addr),
    .io_r_3_cluster_55_data(sram_cluster_0_io_r_3_cluster_55_data),
    .io_r_3_cluster_56_en(sram_cluster_0_io_r_3_cluster_56_en),
    .io_r_3_cluster_56_addr(sram_cluster_0_io_r_3_cluster_56_addr),
    .io_r_3_cluster_56_data(sram_cluster_0_io_r_3_cluster_56_data),
    .io_r_3_cluster_57_en(sram_cluster_0_io_r_3_cluster_57_en),
    .io_r_3_cluster_57_addr(sram_cluster_0_io_r_3_cluster_57_addr),
    .io_r_3_cluster_57_data(sram_cluster_0_io_r_3_cluster_57_data),
    .io_r_3_cluster_58_en(sram_cluster_0_io_r_3_cluster_58_en),
    .io_r_3_cluster_58_addr(sram_cluster_0_io_r_3_cluster_58_addr),
    .io_r_3_cluster_58_data(sram_cluster_0_io_r_3_cluster_58_data),
    .io_r_3_cluster_59_en(sram_cluster_0_io_r_3_cluster_59_en),
    .io_r_3_cluster_59_addr(sram_cluster_0_io_r_3_cluster_59_addr),
    .io_r_3_cluster_59_data(sram_cluster_0_io_r_3_cluster_59_data),
    .io_r_3_cluster_60_en(sram_cluster_0_io_r_3_cluster_60_en),
    .io_r_3_cluster_60_addr(sram_cluster_0_io_r_3_cluster_60_addr),
    .io_r_3_cluster_60_data(sram_cluster_0_io_r_3_cluster_60_data),
    .io_r_3_cluster_61_en(sram_cluster_0_io_r_3_cluster_61_en),
    .io_r_3_cluster_61_addr(sram_cluster_0_io_r_3_cluster_61_addr),
    .io_r_3_cluster_61_data(sram_cluster_0_io_r_3_cluster_61_data),
    .io_r_3_cluster_62_en(sram_cluster_0_io_r_3_cluster_62_en),
    .io_r_3_cluster_62_addr(sram_cluster_0_io_r_3_cluster_62_addr),
    .io_r_3_cluster_62_data(sram_cluster_0_io_r_3_cluster_62_data),
    .io_r_3_cluster_63_en(sram_cluster_0_io_r_3_cluster_63_en),
    .io_r_3_cluster_63_addr(sram_cluster_0_io_r_3_cluster_63_addr),
    .io_r_3_cluster_63_data(sram_cluster_0_io_r_3_cluster_63_data)
  );
  Initializer init ( // @[ipsa.scala 80:22]
    .clock(init_clock),
    .io_pipe_phv_in_data_0(init_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(init_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(init_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(init_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(init_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(init_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(init_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(init_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(init_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(init_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(init_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(init_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(init_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(init_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(init_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(init_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(init_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(init_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(init_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(init_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(init_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(init_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(init_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(init_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(init_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(init_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(init_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(init_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(init_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(init_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(init_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(init_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(init_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(init_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(init_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(init_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(init_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(init_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(init_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(init_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(init_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(init_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(init_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(init_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(init_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(init_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(init_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(init_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(init_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(init_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(init_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(init_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(init_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(init_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(init_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(init_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(init_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(init_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(init_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(init_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(init_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(init_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(init_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(init_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(init_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(init_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(init_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(init_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(init_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(init_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(init_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(init_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(init_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(init_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(init_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(init_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(init_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(init_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(init_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(init_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(init_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(init_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(init_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(init_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(init_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(init_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(init_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(init_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(init_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(init_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(init_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(init_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(init_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(init_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(init_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(init_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(init_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(init_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(init_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(init_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(init_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(init_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(init_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(init_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(init_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(init_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(init_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(init_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(init_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(init_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(init_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(init_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(init_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(init_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(init_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(init_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(init_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(init_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(init_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(init_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(init_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(init_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(init_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(init_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(init_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(init_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(init_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(init_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(init_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(init_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(init_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(init_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(init_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(init_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(init_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(init_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(init_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(init_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(init_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(init_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(init_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(init_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(init_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(init_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(init_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(init_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(init_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(init_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(init_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(init_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(init_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(init_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(init_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(init_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(init_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(init_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(init_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(init_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(init_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(init_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(init_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(init_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(init_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(init_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(init_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(init_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(init_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(init_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(init_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(init_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(init_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(init_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(init_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(init_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(init_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(init_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(init_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(init_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(init_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(init_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(init_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(init_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(init_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(init_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(init_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(init_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(init_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(init_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(init_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(init_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(init_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(init_io_pipe_phv_in_data_191),
    .io_pipe_phv_out_data_0(init_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(init_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(init_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(init_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(init_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(init_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(init_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(init_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(init_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(init_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(init_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(init_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(init_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(init_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(init_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(init_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(init_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(init_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(init_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(init_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(init_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(init_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(init_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(init_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(init_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(init_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(init_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(init_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(init_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(init_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(init_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(init_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(init_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(init_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(init_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(init_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(init_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(init_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(init_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(init_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(init_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(init_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(init_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(init_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(init_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(init_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(init_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(init_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(init_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(init_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(init_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(init_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(init_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(init_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(init_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(init_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(init_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(init_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(init_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(init_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(init_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(init_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(init_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(init_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(init_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(init_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(init_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(init_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(init_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(init_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(init_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(init_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(init_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(init_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(init_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(init_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(init_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(init_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(init_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(init_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(init_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(init_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(init_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(init_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(init_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(init_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(init_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(init_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(init_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(init_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(init_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(init_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(init_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(init_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(init_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(init_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(init_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(init_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(init_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(init_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(init_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(init_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(init_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(init_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(init_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(init_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(init_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(init_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(init_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(init_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(init_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(init_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(init_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(init_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(init_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(init_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(init_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(init_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(init_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(init_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(init_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(init_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(init_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(init_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(init_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(init_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(init_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(init_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(init_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(init_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(init_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(init_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(init_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(init_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(init_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(init_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(init_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(init_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(init_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(init_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(init_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(init_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(init_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(init_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(init_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(init_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(init_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(init_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(init_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(init_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(init_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(init_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(init_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(init_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(init_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(init_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(init_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(init_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(init_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(init_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(init_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(init_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(init_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(init_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(init_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(init_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(init_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(init_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(init_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(init_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(init_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(init_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(init_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(init_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(init_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(init_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(init_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(init_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(init_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(init_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(init_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(init_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(init_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(init_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(init_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(init_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(init_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(init_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(init_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(init_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(init_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(init_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_next_processor_id(init_io_pipe_phv_out_next_processor_id),
    .io_first_proc_id(init_io_first_proc_id)
  );
  InterProcessorTransfer trans_0 ( // @[ipsa.scala 85:25]
    .clock(trans_0_clock),
    .io_pipe_phv_in_data_0(trans_0_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_0_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_0_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_0_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_0_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_0_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_0_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_0_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_0_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_0_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_0_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_0_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_0_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_0_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_0_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_0_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_0_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_0_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_0_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_0_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_0_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_0_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_0_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_0_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_0_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_0_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_0_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_0_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_0_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_0_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_0_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_0_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_0_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_0_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_0_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_0_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_0_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_0_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_0_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_0_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_0_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_0_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_0_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_0_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_0_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_0_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_0_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_0_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_0_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_0_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_0_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_0_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_0_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_0_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_0_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_0_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_0_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_0_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_0_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_0_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_0_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_0_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_0_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_0_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_0_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_0_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_0_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_0_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_0_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_0_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_0_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_0_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_0_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_0_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_0_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_0_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_0_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_0_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_0_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_0_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_0_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_0_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_0_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_0_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_0_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_0_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_0_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_0_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_0_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_0_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_0_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_0_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_0_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_0_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_0_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_0_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_0_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_0_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_0_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_0_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_0_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_0_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_0_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_0_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_0_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_0_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_0_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_0_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_0_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_0_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_0_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_0_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_0_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_0_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_0_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_0_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_0_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_0_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_0_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_0_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_0_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_0_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_0_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_0_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_0_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_0_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_0_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_0_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_0_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_0_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_0_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_0_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_0_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_0_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_0_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_0_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_0_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_0_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_0_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_0_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_0_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_0_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_0_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_0_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_0_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_0_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_0_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_0_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_0_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_0_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_0_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_0_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_0_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_0_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_0_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_0_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_0_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_0_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_0_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_0_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(trans_0_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(trans_0_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(trans_0_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(trans_0_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(trans_0_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(trans_0_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(trans_0_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(trans_0_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(trans_0_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(trans_0_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(trans_0_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(trans_0_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(trans_0_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(trans_0_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(trans_0_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(trans_0_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(trans_0_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(trans_0_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(trans_0_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(trans_0_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(trans_0_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(trans_0_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(trans_0_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(trans_0_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(trans_0_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(trans_0_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(trans_0_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(trans_0_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(trans_0_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(trans_0_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(trans_0_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(trans_0_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(trans_0_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(trans_0_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(trans_0_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(trans_0_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(trans_0_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(trans_0_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(trans_0_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(trans_0_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(trans_0_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(trans_0_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(trans_0_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(trans_0_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(trans_0_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(trans_0_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(trans_0_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(trans_0_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(trans_0_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(trans_0_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(trans_0_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(trans_0_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(trans_0_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(trans_0_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(trans_0_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(trans_0_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(trans_0_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(trans_0_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(trans_0_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(trans_0_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(trans_0_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(trans_0_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(trans_0_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(trans_0_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(trans_0_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(trans_0_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(trans_0_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(trans_0_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(trans_0_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(trans_0_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(trans_0_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(trans_0_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(trans_0_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(trans_0_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(trans_0_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(trans_0_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(trans_0_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(trans_0_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(trans_0_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(trans_0_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(trans_0_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(trans_0_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(trans_0_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(trans_0_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(trans_0_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(trans_0_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(trans_0_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(trans_0_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(trans_0_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(trans_0_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(trans_0_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(trans_0_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(trans_0_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(trans_0_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(trans_0_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(trans_0_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(trans_0_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_0_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_0_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_0_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_0_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_0_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_0_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_0_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_0_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_0_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_0_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_0_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_0_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_0_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_0_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_0_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_0_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_0_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_0_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_0_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_0_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_out_data_0(trans_0_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_0_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_0_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_0_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_0_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_0_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_0_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_0_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_0_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_0_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_0_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_0_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_0_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_0_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_0_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_0_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_0_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_0_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_0_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_0_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_0_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_0_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_0_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_0_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_0_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_0_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_0_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_0_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_0_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_0_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_0_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_0_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_0_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_0_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_0_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_0_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_0_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_0_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_0_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_0_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_0_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_0_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_0_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_0_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_0_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_0_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_0_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_0_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_0_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_0_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_0_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_0_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_0_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_0_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_0_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_0_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_0_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_0_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_0_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_0_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_0_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_0_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_0_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_0_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_0_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_0_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_0_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_0_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_0_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_0_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_0_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_0_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_0_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_0_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_0_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_0_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_0_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_0_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_0_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_0_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_0_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_0_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_0_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_0_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_0_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_0_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_0_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_0_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_0_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_0_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_0_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_0_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_0_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_0_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_0_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_0_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_0_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_0_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_0_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_0_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_0_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_0_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_0_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_0_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_0_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_0_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_0_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_0_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_0_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_0_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_0_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_0_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_0_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_0_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_0_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_0_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_0_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_0_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_0_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_0_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_0_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_0_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_0_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_0_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_0_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_0_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_0_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_0_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_0_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_0_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_0_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_0_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_0_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_0_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_0_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_0_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_0_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_0_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_0_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_0_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_0_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_0_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_0_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_0_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_0_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_0_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_0_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_0_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_0_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_0_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_0_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_0_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_0_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_0_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_0_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_0_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_0_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_0_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_0_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_0_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(trans_0_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(trans_0_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(trans_0_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(trans_0_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(trans_0_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(trans_0_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(trans_0_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(trans_0_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(trans_0_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(trans_0_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(trans_0_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(trans_0_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(trans_0_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(trans_0_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(trans_0_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(trans_0_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(trans_0_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(trans_0_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(trans_0_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(trans_0_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(trans_0_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(trans_0_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(trans_0_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(trans_0_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(trans_0_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(trans_0_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(trans_0_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(trans_0_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(trans_0_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(trans_0_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(trans_0_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(trans_0_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(trans_0_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(trans_0_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(trans_0_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(trans_0_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(trans_0_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(trans_0_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(trans_0_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(trans_0_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(trans_0_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(trans_0_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(trans_0_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(trans_0_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(trans_0_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(trans_0_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(trans_0_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(trans_0_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(trans_0_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(trans_0_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(trans_0_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(trans_0_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(trans_0_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(trans_0_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(trans_0_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(trans_0_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(trans_0_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(trans_0_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(trans_0_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(trans_0_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(trans_0_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(trans_0_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(trans_0_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(trans_0_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(trans_0_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(trans_0_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(trans_0_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(trans_0_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(trans_0_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(trans_0_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(trans_0_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(trans_0_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(trans_0_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(trans_0_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(trans_0_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(trans_0_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(trans_0_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(trans_0_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(trans_0_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(trans_0_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(trans_0_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(trans_0_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(trans_0_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(trans_0_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(trans_0_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(trans_0_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(trans_0_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(trans_0_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(trans_0_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(trans_0_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(trans_0_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(trans_0_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(trans_0_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(trans_0_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(trans_0_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(trans_0_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(trans_0_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_0_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_0_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_0_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_0_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_0_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_0_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_0_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_0_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_0_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_0_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_0_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_0_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_0_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_0_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_0_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_0_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_0_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_0_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_0_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_0_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_0_io_pipe_phv_out_is_valid_processor),
    .io_next_proc_exist(trans_0_io_next_proc_exist),
    .io_next_proc_id_in(trans_0_io_next_proc_id_in),
    .io_next_proc_id_out(trans_0_io_next_proc_id_out)
  );
  InterProcessorTransfer trans_1 ( // @[ipsa.scala 85:25]
    .clock(trans_1_clock),
    .io_pipe_phv_in_data_0(trans_1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(trans_1_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(trans_1_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(trans_1_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(trans_1_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(trans_1_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(trans_1_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(trans_1_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(trans_1_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(trans_1_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(trans_1_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(trans_1_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(trans_1_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(trans_1_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(trans_1_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(trans_1_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(trans_1_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(trans_1_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(trans_1_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(trans_1_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(trans_1_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(trans_1_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(trans_1_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(trans_1_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(trans_1_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(trans_1_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(trans_1_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(trans_1_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(trans_1_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(trans_1_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(trans_1_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(trans_1_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(trans_1_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(trans_1_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(trans_1_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(trans_1_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(trans_1_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(trans_1_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(trans_1_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(trans_1_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(trans_1_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(trans_1_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(trans_1_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(trans_1_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(trans_1_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(trans_1_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(trans_1_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(trans_1_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(trans_1_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(trans_1_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(trans_1_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(trans_1_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(trans_1_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(trans_1_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(trans_1_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(trans_1_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(trans_1_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(trans_1_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(trans_1_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(trans_1_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(trans_1_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(trans_1_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(trans_1_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(trans_1_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(trans_1_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(trans_1_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(trans_1_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(trans_1_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(trans_1_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(trans_1_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(trans_1_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(trans_1_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(trans_1_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(trans_1_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(trans_1_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(trans_1_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(trans_1_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(trans_1_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(trans_1_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(trans_1_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(trans_1_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(trans_1_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(trans_1_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(trans_1_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(trans_1_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(trans_1_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(trans_1_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(trans_1_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(trans_1_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(trans_1_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(trans_1_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(trans_1_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(trans_1_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(trans_1_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(trans_1_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(trans_1_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(trans_1_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(trans_1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_out_data_0(trans_1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(trans_1_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(trans_1_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(trans_1_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(trans_1_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(trans_1_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(trans_1_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(trans_1_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(trans_1_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(trans_1_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(trans_1_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(trans_1_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(trans_1_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(trans_1_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(trans_1_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(trans_1_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(trans_1_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(trans_1_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(trans_1_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(trans_1_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(trans_1_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(trans_1_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(trans_1_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(trans_1_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(trans_1_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(trans_1_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(trans_1_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(trans_1_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(trans_1_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(trans_1_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(trans_1_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(trans_1_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(trans_1_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(trans_1_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(trans_1_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(trans_1_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(trans_1_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(trans_1_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(trans_1_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(trans_1_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(trans_1_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(trans_1_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(trans_1_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(trans_1_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(trans_1_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(trans_1_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(trans_1_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(trans_1_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(trans_1_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(trans_1_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(trans_1_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(trans_1_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(trans_1_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(trans_1_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(trans_1_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(trans_1_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(trans_1_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(trans_1_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(trans_1_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(trans_1_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(trans_1_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(trans_1_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(trans_1_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(trans_1_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(trans_1_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(trans_1_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(trans_1_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(trans_1_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(trans_1_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(trans_1_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(trans_1_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(trans_1_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(trans_1_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(trans_1_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(trans_1_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(trans_1_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(trans_1_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(trans_1_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(trans_1_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(trans_1_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(trans_1_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(trans_1_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(trans_1_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(trans_1_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(trans_1_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(trans_1_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(trans_1_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(trans_1_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(trans_1_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(trans_1_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(trans_1_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(trans_1_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(trans_1_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(trans_1_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(trans_1_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(trans_1_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(trans_1_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(trans_1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_1_io_pipe_phv_out_is_valid_processor),
    .io_next_proc_exist(trans_1_io_next_proc_exist),
    .io_next_proc_id_in(trans_1_io_next_proc_id_in),
    .io_next_proc_id_out(trans_1_io_next_proc_id_out)
  );
  InterProcessorTransfer trans_2 ( // @[ipsa.scala 85:25]
    .clock(trans_2_clock),
    .io_pipe_phv_in_data_0(trans_2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(trans_2_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(trans_2_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(trans_2_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(trans_2_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(trans_2_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(trans_2_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(trans_2_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(trans_2_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(trans_2_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(trans_2_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(trans_2_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(trans_2_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(trans_2_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(trans_2_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(trans_2_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(trans_2_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(trans_2_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(trans_2_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(trans_2_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(trans_2_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(trans_2_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(trans_2_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(trans_2_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(trans_2_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(trans_2_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(trans_2_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(trans_2_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(trans_2_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(trans_2_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(trans_2_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(trans_2_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(trans_2_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(trans_2_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(trans_2_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(trans_2_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(trans_2_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(trans_2_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(trans_2_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(trans_2_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(trans_2_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(trans_2_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(trans_2_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(trans_2_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(trans_2_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(trans_2_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(trans_2_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(trans_2_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(trans_2_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(trans_2_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(trans_2_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(trans_2_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(trans_2_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(trans_2_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(trans_2_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(trans_2_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(trans_2_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(trans_2_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(trans_2_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(trans_2_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(trans_2_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(trans_2_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(trans_2_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(trans_2_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(trans_2_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(trans_2_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(trans_2_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(trans_2_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(trans_2_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(trans_2_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(trans_2_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(trans_2_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(trans_2_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(trans_2_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(trans_2_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(trans_2_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(trans_2_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(trans_2_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(trans_2_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(trans_2_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(trans_2_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(trans_2_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(trans_2_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(trans_2_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(trans_2_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(trans_2_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(trans_2_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(trans_2_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(trans_2_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(trans_2_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(trans_2_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(trans_2_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(trans_2_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(trans_2_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(trans_2_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(trans_2_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(trans_2_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(trans_2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_out_data_0(trans_2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(trans_2_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(trans_2_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(trans_2_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(trans_2_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(trans_2_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(trans_2_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(trans_2_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(trans_2_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(trans_2_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(trans_2_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(trans_2_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(trans_2_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(trans_2_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(trans_2_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(trans_2_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(trans_2_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(trans_2_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(trans_2_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(trans_2_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(trans_2_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(trans_2_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(trans_2_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(trans_2_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(trans_2_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(trans_2_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(trans_2_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(trans_2_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(trans_2_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(trans_2_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(trans_2_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(trans_2_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(trans_2_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(trans_2_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(trans_2_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(trans_2_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(trans_2_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(trans_2_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(trans_2_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(trans_2_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(trans_2_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(trans_2_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(trans_2_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(trans_2_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(trans_2_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(trans_2_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(trans_2_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(trans_2_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(trans_2_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(trans_2_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(trans_2_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(trans_2_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(trans_2_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(trans_2_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(trans_2_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(trans_2_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(trans_2_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(trans_2_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(trans_2_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(trans_2_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(trans_2_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(trans_2_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(trans_2_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(trans_2_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(trans_2_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(trans_2_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(trans_2_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(trans_2_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(trans_2_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(trans_2_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(trans_2_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(trans_2_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(trans_2_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(trans_2_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(trans_2_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(trans_2_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(trans_2_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(trans_2_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(trans_2_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(trans_2_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(trans_2_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(trans_2_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(trans_2_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(trans_2_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(trans_2_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(trans_2_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(trans_2_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(trans_2_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(trans_2_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(trans_2_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(trans_2_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(trans_2_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(trans_2_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(trans_2_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(trans_2_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(trans_2_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(trans_2_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(trans_2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_2_io_pipe_phv_out_is_valid_processor),
    .io_next_proc_exist(trans_2_io_next_proc_exist),
    .io_next_proc_id_in(trans_2_io_next_proc_id_in),
    .io_next_proc_id_out(trans_2_io_next_proc_id_out)
  );
  InterProcessorTransfer trans_3 ( // @[ipsa.scala 85:25]
    .clock(trans_3_clock),
    .io_pipe_phv_in_data_0(trans_3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(trans_3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(trans_3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(trans_3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(trans_3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(trans_3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(trans_3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(trans_3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(trans_3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(trans_3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(trans_3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(trans_3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(trans_3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(trans_3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(trans_3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(trans_3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(trans_3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(trans_3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(trans_3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(trans_3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(trans_3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(trans_3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(trans_3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(trans_3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(trans_3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(trans_3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(trans_3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(trans_3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(trans_3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(trans_3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(trans_3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(trans_3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(trans_3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(trans_3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(trans_3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(trans_3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(trans_3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(trans_3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(trans_3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(trans_3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(trans_3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(trans_3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(trans_3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(trans_3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(trans_3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(trans_3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(trans_3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(trans_3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(trans_3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(trans_3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(trans_3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(trans_3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(trans_3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(trans_3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(trans_3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(trans_3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(trans_3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(trans_3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(trans_3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(trans_3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(trans_3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(trans_3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(trans_3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(trans_3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(trans_3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(trans_3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(trans_3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(trans_3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(trans_3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(trans_3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(trans_3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(trans_3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(trans_3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(trans_3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(trans_3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(trans_3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(trans_3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(trans_3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(trans_3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(trans_3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(trans_3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(trans_3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(trans_3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(trans_3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(trans_3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(trans_3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(trans_3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(trans_3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(trans_3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(trans_3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(trans_3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(trans_3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(trans_3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(trans_3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(trans_3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(trans_3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(trans_3_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(trans_3_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(trans_3_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(trans_3_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(trans_3_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(trans_3_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(trans_3_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(trans_3_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(trans_3_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(trans_3_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(trans_3_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(trans_3_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(trans_3_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(trans_3_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(trans_3_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(trans_3_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(trans_3_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(trans_3_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(trans_3_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(trans_3_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(trans_3_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(trans_3_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(trans_3_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(trans_3_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(trans_3_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(trans_3_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(trans_3_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(trans_3_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(trans_3_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(trans_3_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(trans_3_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(trans_3_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(trans_3_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(trans_3_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(trans_3_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(trans_3_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(trans_3_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(trans_3_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(trans_3_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(trans_3_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(trans_3_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(trans_3_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(trans_3_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(trans_3_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(trans_3_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(trans_3_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(trans_3_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(trans_3_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(trans_3_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(trans_3_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(trans_3_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(trans_3_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(trans_3_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(trans_3_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(trans_3_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(trans_3_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(trans_3_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(trans_3_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(trans_3_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(trans_3_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(trans_3_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(trans_3_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(trans_3_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(trans_3_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(trans_3_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(trans_3_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(trans_3_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(trans_3_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(trans_3_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(trans_3_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(trans_3_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(trans_3_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(trans_3_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(trans_3_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(trans_3_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(trans_3_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(trans_3_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(trans_3_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(trans_3_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(trans_3_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(trans_3_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(trans_3_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(trans_3_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(trans_3_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(trans_3_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(trans_3_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(trans_3_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(trans_3_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(trans_3_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(trans_3_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(trans_3_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(trans_3_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(trans_3_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(trans_3_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(trans_3_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(trans_3_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(trans_3_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(trans_3_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(trans_3_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(trans_3_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(trans_3_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(trans_3_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(trans_3_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(trans_3_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(trans_3_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(trans_3_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(trans_3_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(trans_3_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(trans_3_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(trans_3_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(trans_3_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(trans_3_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(trans_3_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(trans_3_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(trans_3_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(trans_3_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(trans_3_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(trans_3_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(trans_3_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(trans_3_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(trans_3_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(trans_3_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(trans_3_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(trans_3_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(trans_3_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(trans_3_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(trans_3_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(trans_3_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(trans_3_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(trans_3_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(trans_3_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(trans_3_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(trans_3_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(trans_3_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(trans_3_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(trans_3_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(trans_3_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(trans_3_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(trans_3_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(trans_3_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(trans_3_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(trans_3_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(trans_3_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(trans_3_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(trans_3_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(trans_3_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(trans_3_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(trans_3_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(trans_3_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(trans_3_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(trans_3_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(trans_3_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(trans_3_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(trans_3_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(trans_3_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(trans_3_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(trans_3_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(trans_3_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(trans_3_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(trans_3_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(trans_3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(trans_3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(trans_3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(trans_3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(trans_3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(trans_3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(trans_3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(trans_3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(trans_3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(trans_3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(trans_3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(trans_3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(trans_3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(trans_3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(trans_3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(trans_3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(trans_3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(trans_3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(trans_3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(trans_3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(trans_3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_out_data_0(trans_3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(trans_3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(trans_3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(trans_3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(trans_3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(trans_3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(trans_3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(trans_3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(trans_3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(trans_3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(trans_3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(trans_3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(trans_3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(trans_3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(trans_3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(trans_3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(trans_3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(trans_3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(trans_3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(trans_3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(trans_3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(trans_3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(trans_3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(trans_3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(trans_3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(trans_3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(trans_3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(trans_3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(trans_3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(trans_3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(trans_3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(trans_3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(trans_3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(trans_3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(trans_3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(trans_3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(trans_3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(trans_3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(trans_3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(trans_3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(trans_3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(trans_3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(trans_3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(trans_3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(trans_3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(trans_3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(trans_3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(trans_3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(trans_3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(trans_3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(trans_3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(trans_3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(trans_3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(trans_3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(trans_3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(trans_3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(trans_3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(trans_3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(trans_3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(trans_3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(trans_3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(trans_3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(trans_3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(trans_3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(trans_3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(trans_3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(trans_3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(trans_3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(trans_3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(trans_3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(trans_3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(trans_3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(trans_3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(trans_3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(trans_3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(trans_3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(trans_3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(trans_3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(trans_3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(trans_3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(trans_3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(trans_3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(trans_3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(trans_3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(trans_3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(trans_3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(trans_3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(trans_3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(trans_3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(trans_3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(trans_3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(trans_3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(trans_3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(trans_3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(trans_3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(trans_3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(trans_3_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(trans_3_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(trans_3_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(trans_3_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(trans_3_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(trans_3_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(trans_3_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(trans_3_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(trans_3_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(trans_3_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(trans_3_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(trans_3_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(trans_3_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(trans_3_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(trans_3_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(trans_3_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(trans_3_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(trans_3_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(trans_3_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(trans_3_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(trans_3_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(trans_3_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(trans_3_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(trans_3_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(trans_3_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(trans_3_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(trans_3_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(trans_3_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(trans_3_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(trans_3_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(trans_3_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(trans_3_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(trans_3_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(trans_3_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(trans_3_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(trans_3_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(trans_3_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(trans_3_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(trans_3_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(trans_3_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(trans_3_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(trans_3_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(trans_3_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(trans_3_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(trans_3_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(trans_3_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(trans_3_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(trans_3_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(trans_3_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(trans_3_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(trans_3_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(trans_3_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(trans_3_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(trans_3_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(trans_3_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(trans_3_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(trans_3_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(trans_3_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(trans_3_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(trans_3_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(trans_3_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(trans_3_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(trans_3_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(trans_3_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(trans_3_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(trans_3_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(trans_3_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(trans_3_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(trans_3_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(trans_3_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(trans_3_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(trans_3_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(trans_3_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(trans_3_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(trans_3_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(trans_3_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(trans_3_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(trans_3_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(trans_3_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(trans_3_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(trans_3_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(trans_3_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(trans_3_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(trans_3_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(trans_3_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(trans_3_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(trans_3_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(trans_3_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(trans_3_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(trans_3_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(trans_3_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(trans_3_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(trans_3_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(trans_3_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(trans_3_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(trans_3_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(trans_3_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(trans_3_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(trans_3_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(trans_3_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(trans_3_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(trans_3_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(trans_3_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(trans_3_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(trans_3_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(trans_3_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(trans_3_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(trans_3_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(trans_3_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(trans_3_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(trans_3_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(trans_3_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(trans_3_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(trans_3_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(trans_3_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(trans_3_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(trans_3_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(trans_3_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(trans_3_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(trans_3_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(trans_3_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(trans_3_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(trans_3_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(trans_3_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(trans_3_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(trans_3_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(trans_3_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(trans_3_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(trans_3_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(trans_3_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(trans_3_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(trans_3_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(trans_3_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(trans_3_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(trans_3_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(trans_3_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(trans_3_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(trans_3_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(trans_3_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(trans_3_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(trans_3_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(trans_3_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(trans_3_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(trans_3_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(trans_3_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(trans_3_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(trans_3_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(trans_3_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(trans_3_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(trans_3_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(trans_3_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(trans_3_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(trans_3_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(trans_3_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(trans_3_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(trans_3_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(trans_3_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(trans_3_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(trans_3_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(trans_3_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(trans_3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(trans_3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(trans_3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(trans_3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(trans_3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(trans_3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(trans_3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(trans_3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(trans_3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(trans_3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(trans_3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(trans_3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(trans_3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(trans_3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(trans_3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(trans_3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(trans_3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(trans_3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(trans_3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(trans_3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(trans_3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(trans_3_io_pipe_phv_out_is_valid_processor),
    .io_next_proc_exist(trans_3_io_next_proc_exist),
    .io_next_proc_id_in(trans_3_io_next_proc_id_in),
    .io_next_proc_id_out(trans_3_io_next_proc_id_out)
  );
  assign io_pipe_phv_out_data_0 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_0 : _GEN_584; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_1 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_1 : _GEN_585; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_2 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_2 : _GEN_586; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_3 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_3 : _GEN_587; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_4 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_4 : _GEN_588; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_5 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_5 : _GEN_589; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_6 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_6 : _GEN_590; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_7 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_7 : _GEN_591; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_8 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_8 : _GEN_592; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_9 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_9 : _GEN_593; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_10 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_10 : _GEN_594; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_11 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_11 : _GEN_595; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_12 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_12 : _GEN_596; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_13 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_13 : _GEN_597; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_14 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_14 : _GEN_598; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_15 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_15 : _GEN_599; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_16 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_16 : _GEN_600; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_17 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_17 : _GEN_601; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_18 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_18 : _GEN_602; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_19 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_19 : _GEN_603; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_20 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_20 : _GEN_604; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_21 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_21 : _GEN_605; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_22 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_22 : _GEN_606; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_23 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_23 : _GEN_607; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_24 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_24 : _GEN_608; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_25 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_25 : _GEN_609; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_26 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_26 : _GEN_610; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_27 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_27 : _GEN_611; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_28 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_28 : _GEN_612; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_29 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_29 : _GEN_613; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_30 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_30 : _GEN_614; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_31 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_31 : _GEN_615; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_32 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_32 : _GEN_616; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_33 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_33 : _GEN_617; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_34 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_34 : _GEN_618; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_35 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_35 : _GEN_619; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_36 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_36 : _GEN_620; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_37 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_37 : _GEN_621; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_38 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_38 : _GEN_622; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_39 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_39 : _GEN_623; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_40 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_40 : _GEN_624; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_41 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_41 : _GEN_625; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_42 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_42 : _GEN_626; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_43 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_43 : _GEN_627; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_44 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_44 : _GEN_628; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_45 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_45 : _GEN_629; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_46 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_46 : _GEN_630; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_47 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_47 : _GEN_631; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_48 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_48 : _GEN_632; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_49 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_49 : _GEN_633; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_50 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_50 : _GEN_634; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_51 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_51 : _GEN_635; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_52 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_52 : _GEN_636; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_53 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_53 : _GEN_637; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_54 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_54 : _GEN_638; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_55 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_55 : _GEN_639; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_56 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_56 : _GEN_640; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_57 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_57 : _GEN_641; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_58 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_58 : _GEN_642; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_59 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_59 : _GEN_643; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_60 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_60 : _GEN_644; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_61 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_61 : _GEN_645; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_62 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_62 : _GEN_646; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_63 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_63 : _GEN_647; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_64 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_64 : _GEN_648; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_65 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_65 : _GEN_649; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_66 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_66 : _GEN_650; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_67 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_67 : _GEN_651; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_68 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_68 : _GEN_652; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_69 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_69 : _GEN_653; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_70 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_70 : _GEN_654; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_71 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_71 : _GEN_655; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_72 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_72 : _GEN_656; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_73 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_73 : _GEN_657; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_74 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_74 : _GEN_658; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_75 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_75 : _GEN_659; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_76 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_76 : _GEN_660; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_77 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_77 : _GEN_661; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_78 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_78 : _GEN_662; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_79 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_79 : _GEN_663; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_80 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_80 : _GEN_664; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_81 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_81 : _GEN_665; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_82 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_82 : _GEN_666; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_83 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_83 : _GEN_667; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_84 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_84 : _GEN_668; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_85 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_85 : _GEN_669; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_86 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_86 : _GEN_670; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_87 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_87 : _GEN_671; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_88 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_88 : _GEN_672; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_89 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_89 : _GEN_673; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_90 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_90 : _GEN_674; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_91 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_91 : _GEN_675; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_92 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_92 : _GEN_676; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_93 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_93 : _GEN_677; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_94 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_94 : _GEN_678; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_95 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_95 : _GEN_679; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_96 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_96 : _GEN_680; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_97 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_97 : _GEN_681; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_98 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_98 : _GEN_682; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_99 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_99 : _GEN_683; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_100 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_100 : _GEN_684; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_101 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_101 : _GEN_685; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_102 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_102 : _GEN_686; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_103 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_103 : _GEN_687; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_104 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_104 : _GEN_688; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_105 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_105 : _GEN_689; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_106 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_106 : _GEN_690; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_107 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_107 : _GEN_691; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_108 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_108 : _GEN_692; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_109 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_109 : _GEN_693; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_110 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_110 : _GEN_694; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_111 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_111 : _GEN_695; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_112 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_112 : _GEN_696; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_113 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_113 : _GEN_697; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_114 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_114 : _GEN_698; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_115 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_115 : _GEN_699; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_116 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_116 : _GEN_700; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_117 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_117 : _GEN_701; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_118 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_118 : _GEN_702; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_119 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_119 : _GEN_703; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_120 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_120 : _GEN_704; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_121 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_121 : _GEN_705; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_122 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_122 : _GEN_706; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_123 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_123 : _GEN_707; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_124 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_124 : _GEN_708; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_125 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_125 : _GEN_709; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_126 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_126 : _GEN_710; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_127 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_127 : _GEN_711; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_128 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_128 : _GEN_712; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_129 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_129 : _GEN_713; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_130 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_130 : _GEN_714; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_131 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_131 : _GEN_715; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_132 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_132 : _GEN_716; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_133 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_133 : _GEN_717; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_134 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_134 : _GEN_718; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_135 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_135 : _GEN_719; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_136 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_136 : _GEN_720; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_137 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_137 : _GEN_721; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_138 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_138 : _GEN_722; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_139 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_139 : _GEN_723; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_140 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_140 : _GEN_724; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_141 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_141 : _GEN_725; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_142 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_142 : _GEN_726; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_143 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_143 : _GEN_727; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_144 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_144 : _GEN_728; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_145 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_145 : _GEN_729; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_146 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_146 : _GEN_730; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_147 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_147 : _GEN_731; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_148 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_148 : _GEN_732; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_149 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_149 : _GEN_733; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_150 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_150 : _GEN_734; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_151 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_151 : _GEN_735; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_152 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_152 : _GEN_736; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_153 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_153 : _GEN_737; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_154 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_154 : _GEN_738; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_155 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_155 : _GEN_739; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_156 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_156 : _GEN_740; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_157 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_157 : _GEN_741; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_158 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_158 : _GEN_742; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_159 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_159 : _GEN_743; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_160 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_160 : _GEN_744; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_161 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_161 : _GEN_745; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_162 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_162 : _GEN_746; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_163 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_163 : _GEN_747; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_164 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_164 : _GEN_748; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_165 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_165 : _GEN_749; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_166 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_166 : _GEN_750; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_167 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_167 : _GEN_751; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_168 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_168 : _GEN_752; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_169 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_169 : _GEN_753; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_170 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_170 : _GEN_754; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_171 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_171 : _GEN_755; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_172 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_172 : _GEN_756; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_173 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_173 : _GEN_757; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_174 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_174 : _GEN_758; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_175 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_175 : _GEN_759; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_176 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_176 : _GEN_760; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_177 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_177 : _GEN_761; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_178 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_178 : _GEN_762; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_179 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_179 : _GEN_763; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_180 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_180 : _GEN_764; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_181 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_181 : _GEN_765; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_182 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_182 : _GEN_766; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_183 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_183 : _GEN_767; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_184 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_184 : _GEN_768; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_185 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_185 : _GEN_769; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_186 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_186 : _GEN_770; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_187 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_187 : _GEN_771; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_188 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_188 : _GEN_772; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_189 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_189 : _GEN_773; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_190 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_190 : _GEN_774; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_191 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_191 : _GEN_775; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_192 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_192 : _GEN_776; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_193 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_193 : _GEN_777; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_194 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_194 : _GEN_778; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_195 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_195 : _GEN_779; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_196 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_196 : _GEN_780; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_197 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_197 : _GEN_781; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_198 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_198 : _GEN_782; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_199 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_199 : _GEN_783; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_200 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_200 : _GEN_784; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_201 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_201 : _GEN_785; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_202 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_202 : _GEN_786; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_203 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_203 : _GEN_787; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_204 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_204 : _GEN_788; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_205 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_205 : _GEN_789; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_206 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_206 : _GEN_790; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_207 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_207 : _GEN_791; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_208 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_208 : _GEN_792; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_209 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_209 : _GEN_793; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_210 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_210 : _GEN_794; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_211 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_211 : _GEN_795; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_212 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_212 : _GEN_796; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_213 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_213 : _GEN_797; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_214 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_214 : _GEN_798; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_215 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_215 : _GEN_799; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_216 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_216 : _GEN_800; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_217 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_217 : _GEN_801; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_218 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_218 : _GEN_802; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_219 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_219 : _GEN_803; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_220 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_220 : _GEN_804; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_221 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_221 : _GEN_805; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_222 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_222 : _GEN_806; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_223 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_223 : _GEN_807; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_224 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_224 : _GEN_808; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_225 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_225 : _GEN_809; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_226 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_226 : _GEN_810; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_227 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_227 : _GEN_811; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_228 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_228 : _GEN_812; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_229 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_229 : _GEN_813; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_230 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_230 : _GEN_814; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_231 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_231 : _GEN_815; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_232 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_232 : _GEN_816; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_233 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_233 : _GEN_817; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_234 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_234 : _GEN_818; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_235 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_235 : _GEN_819; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_236 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_236 : _GEN_820; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_237 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_237 : _GEN_821; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_238 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_238 : _GEN_822; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_239 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_239 : _GEN_823; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_240 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_240 : _GEN_824; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_241 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_241 : _GEN_825; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_242 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_242 : _GEN_826; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_243 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_243 : _GEN_827; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_244 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_244 : _GEN_828; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_245 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_245 : _GEN_829; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_246 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_246 : _GEN_830; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_247 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_247 : _GEN_831; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_248 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_248 : _GEN_832; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_249 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_249 : _GEN_833; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_250 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_250 : _GEN_834; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_251 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_251 : _GEN_835; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_252 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_252 : _GEN_836; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_253 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_253 : _GEN_837; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_254 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_254 : _GEN_838; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign io_pipe_phv_out_data_255 = 2'h3 == last_proc_id ? trans_3_io_pipe_phv_out_data_255 : _GEN_839; // @[ipsa.scala 96:65 ipsa.scala 97:29]
  assign proc_0_clock = clock;
  assign proc_0_io_pipe_phv_in_data_0 = recv_0_data_0; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_1 = recv_0_data_1; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_2 = recv_0_data_2; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_3 = recv_0_data_3; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_4 = recv_0_data_4; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_5 = recv_0_data_5; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_6 = recv_0_data_6; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_7 = recv_0_data_7; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_8 = recv_0_data_8; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_9 = recv_0_data_9; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_10 = recv_0_data_10; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_11 = recv_0_data_11; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_12 = recv_0_data_12; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_13 = recv_0_data_13; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_14 = recv_0_data_14; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_15 = recv_0_data_15; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_16 = recv_0_data_16; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_17 = recv_0_data_17; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_18 = recv_0_data_18; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_19 = recv_0_data_19; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_20 = recv_0_data_20; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_21 = recv_0_data_21; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_22 = recv_0_data_22; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_23 = recv_0_data_23; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_24 = recv_0_data_24; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_25 = recv_0_data_25; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_26 = recv_0_data_26; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_27 = recv_0_data_27; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_28 = recv_0_data_28; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_29 = recv_0_data_29; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_30 = recv_0_data_30; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_31 = recv_0_data_31; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_32 = recv_0_data_32; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_33 = recv_0_data_33; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_34 = recv_0_data_34; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_35 = recv_0_data_35; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_36 = recv_0_data_36; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_37 = recv_0_data_37; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_38 = recv_0_data_38; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_39 = recv_0_data_39; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_40 = recv_0_data_40; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_41 = recv_0_data_41; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_42 = recv_0_data_42; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_43 = recv_0_data_43; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_44 = recv_0_data_44; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_45 = recv_0_data_45; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_46 = recv_0_data_46; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_47 = recv_0_data_47; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_48 = recv_0_data_48; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_49 = recv_0_data_49; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_50 = recv_0_data_50; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_51 = recv_0_data_51; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_52 = recv_0_data_52; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_53 = recv_0_data_53; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_54 = recv_0_data_54; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_55 = recv_0_data_55; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_56 = recv_0_data_56; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_57 = recv_0_data_57; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_58 = recv_0_data_58; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_59 = recv_0_data_59; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_60 = recv_0_data_60; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_61 = recv_0_data_61; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_62 = recv_0_data_62; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_63 = recv_0_data_63; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_64 = recv_0_data_64; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_65 = recv_0_data_65; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_66 = recv_0_data_66; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_67 = recv_0_data_67; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_68 = recv_0_data_68; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_69 = recv_0_data_69; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_70 = recv_0_data_70; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_71 = recv_0_data_71; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_72 = recv_0_data_72; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_73 = recv_0_data_73; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_74 = recv_0_data_74; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_75 = recv_0_data_75; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_76 = recv_0_data_76; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_77 = recv_0_data_77; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_78 = recv_0_data_78; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_79 = recv_0_data_79; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_80 = recv_0_data_80; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_81 = recv_0_data_81; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_82 = recv_0_data_82; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_83 = recv_0_data_83; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_84 = recv_0_data_84; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_85 = recv_0_data_85; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_86 = recv_0_data_86; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_87 = recv_0_data_87; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_88 = recv_0_data_88; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_89 = recv_0_data_89; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_90 = recv_0_data_90; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_91 = recv_0_data_91; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_92 = recv_0_data_92; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_93 = recv_0_data_93; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_94 = recv_0_data_94; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_95 = recv_0_data_95; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_96 = recv_0_data_96; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_97 = recv_0_data_97; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_98 = recv_0_data_98; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_99 = recv_0_data_99; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_100 = recv_0_data_100; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_101 = recv_0_data_101; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_102 = recv_0_data_102; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_103 = recv_0_data_103; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_104 = recv_0_data_104; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_105 = recv_0_data_105; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_106 = recv_0_data_106; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_107 = recv_0_data_107; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_108 = recv_0_data_108; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_109 = recv_0_data_109; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_110 = recv_0_data_110; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_111 = recv_0_data_111; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_112 = recv_0_data_112; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_113 = recv_0_data_113; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_114 = recv_0_data_114; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_115 = recv_0_data_115; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_116 = recv_0_data_116; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_117 = recv_0_data_117; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_118 = recv_0_data_118; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_119 = recv_0_data_119; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_120 = recv_0_data_120; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_121 = recv_0_data_121; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_122 = recv_0_data_122; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_123 = recv_0_data_123; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_124 = recv_0_data_124; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_125 = recv_0_data_125; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_126 = recv_0_data_126; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_127 = recv_0_data_127; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_128 = recv_0_data_128; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_129 = recv_0_data_129; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_130 = recv_0_data_130; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_131 = recv_0_data_131; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_132 = recv_0_data_132; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_133 = recv_0_data_133; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_134 = recv_0_data_134; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_135 = recv_0_data_135; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_136 = recv_0_data_136; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_137 = recv_0_data_137; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_138 = recv_0_data_138; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_139 = recv_0_data_139; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_140 = recv_0_data_140; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_141 = recv_0_data_141; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_142 = recv_0_data_142; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_143 = recv_0_data_143; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_144 = recv_0_data_144; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_145 = recv_0_data_145; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_146 = recv_0_data_146; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_147 = recv_0_data_147; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_148 = recv_0_data_148; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_149 = recv_0_data_149; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_150 = recv_0_data_150; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_151 = recv_0_data_151; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_152 = recv_0_data_152; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_153 = recv_0_data_153; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_154 = recv_0_data_154; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_155 = recv_0_data_155; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_156 = recv_0_data_156; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_157 = recv_0_data_157; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_158 = recv_0_data_158; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_159 = recv_0_data_159; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_160 = recv_0_data_160; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_161 = recv_0_data_161; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_162 = recv_0_data_162; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_163 = recv_0_data_163; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_164 = recv_0_data_164; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_165 = recv_0_data_165; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_166 = recv_0_data_166; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_167 = recv_0_data_167; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_168 = recv_0_data_168; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_169 = recv_0_data_169; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_170 = recv_0_data_170; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_171 = recv_0_data_171; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_172 = recv_0_data_172; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_173 = recv_0_data_173; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_174 = recv_0_data_174; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_175 = recv_0_data_175; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_176 = recv_0_data_176; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_177 = recv_0_data_177; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_178 = recv_0_data_178; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_179 = recv_0_data_179; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_180 = recv_0_data_180; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_181 = recv_0_data_181; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_182 = recv_0_data_182; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_183 = recv_0_data_183; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_184 = recv_0_data_184; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_185 = recv_0_data_185; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_186 = recv_0_data_186; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_187 = recv_0_data_187; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_188 = recv_0_data_188; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_189 = recv_0_data_189; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_190 = recv_0_data_190; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_191 = recv_0_data_191; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_192 = recv_0_data_192; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_193 = recv_0_data_193; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_194 = recv_0_data_194; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_195 = recv_0_data_195; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_196 = recv_0_data_196; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_197 = recv_0_data_197; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_198 = recv_0_data_198; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_199 = recv_0_data_199; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_200 = recv_0_data_200; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_201 = recv_0_data_201; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_202 = recv_0_data_202; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_203 = recv_0_data_203; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_204 = recv_0_data_204; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_205 = recv_0_data_205; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_206 = recv_0_data_206; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_207 = recv_0_data_207; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_208 = recv_0_data_208; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_209 = recv_0_data_209; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_210 = recv_0_data_210; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_211 = recv_0_data_211; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_212 = recv_0_data_212; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_213 = recv_0_data_213; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_214 = recv_0_data_214; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_215 = recv_0_data_215; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_216 = recv_0_data_216; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_217 = recv_0_data_217; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_218 = recv_0_data_218; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_219 = recv_0_data_219; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_220 = recv_0_data_220; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_221 = recv_0_data_221; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_222 = recv_0_data_222; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_223 = recv_0_data_223; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_224 = recv_0_data_224; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_225 = recv_0_data_225; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_226 = recv_0_data_226; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_227 = recv_0_data_227; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_228 = recv_0_data_228; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_229 = recv_0_data_229; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_230 = recv_0_data_230; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_231 = recv_0_data_231; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_232 = recv_0_data_232; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_233 = recv_0_data_233; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_234 = recv_0_data_234; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_235 = recv_0_data_235; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_236 = recv_0_data_236; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_237 = recv_0_data_237; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_238 = recv_0_data_238; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_239 = recv_0_data_239; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_240 = recv_0_data_240; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_241 = recv_0_data_241; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_242 = recv_0_data_242; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_243 = recv_0_data_243; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_244 = recv_0_data_244; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_245 = recv_0_data_245; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_246 = recv_0_data_246; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_247 = recv_0_data_247; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_248 = recv_0_data_248; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_249 = recv_0_data_249; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_250 = recv_0_data_250; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_251 = recv_0_data_251; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_252 = recv_0_data_252; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_253 = recv_0_data_253; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_254 = recv_0_data_254; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_data_255 = recv_0_data_255; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_header_0 = recv_0_header_0; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_header_1 = recv_0_header_1; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_header_2 = recv_0_header_2; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_header_3 = recv_0_header_3; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_header_4 = recv_0_header_4; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_header_5 = recv_0_header_5; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_header_6 = recv_0_header_6; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_header_7 = recv_0_header_7; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_header_8 = recv_0_header_8; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_header_9 = recv_0_header_9; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_header_10 = recv_0_header_10; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_header_11 = recv_0_header_11; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_header_12 = recv_0_header_12; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_header_13 = recv_0_header_13; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_header_14 = recv_0_header_14; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_header_15 = recv_0_header_15; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_parse_current_state = recv_0_parse_current_state; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_parse_current_offset = recv_0_parse_current_offset; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_parse_transition_field = recv_0_parse_transition_field; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_next_processor_id = recv_0_next_processor_id; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_next_config_id = recv_0_next_config_id; // @[ipsa.scala 161:32]
  assign proc_0_io_pipe_phv_in_is_valid_processor = recv_0_is_valid_processor; // @[ipsa.scala 161:32]
  assign proc_0_io_mod_par_mod_en = io_mod_proc_mod_0_par_mod_en; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_par_mod_last_mau_id_mod = io_mod_proc_mod_0_par_mod_last_mau_id_mod; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_par_mod_last_mau_id = io_mod_proc_mod_0_par_mod_last_mau_id; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_par_mod_cs = io_mod_proc_mod_0_par_mod_cs; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_par_mod_module_mod_state_id_mod = io_mod_proc_mod_0_par_mod_module_mod_state_id_mod; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_par_mod_module_mod_state_id = io_mod_proc_mod_0_par_mod_module_mod_state_id; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_par_mod_module_mod_sram_w_cs = io_mod_proc_mod_0_par_mod_module_mod_sram_w_cs; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_par_mod_module_mod_sram_w_en = io_mod_proc_mod_0_par_mod_module_mod_sram_w_en; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_par_mod_module_mod_sram_w_addr = io_mod_proc_mod_0_par_mod_module_mod_sram_w_addr; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_par_mod_module_mod_sram_w_data = io_mod_proc_mod_0_par_mod_module_mod_sram_w_data; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_en = io_mod_proc_mod_0_mat_mod_en; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_config_id = io_mod_proc_mod_0_mat_mod_config_id; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_key_mod_header_id = io_mod_proc_mod_0_mat_mod_key_mod_header_id; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_key_mod_internal_offset = io_mod_proc_mod_0_mat_mod_key_mod_internal_offset; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_key_mod_key_length = io_mod_proc_mod_0_mat_mod_key_mod_key_length; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_0 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_0; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_1 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_1; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_2 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_2; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_3 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_3; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_4 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_4; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_5 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_5; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_6 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_6; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_7 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_7; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_8 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_8; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_9 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_9; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_10 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_10; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_11 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_11; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_12 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_12; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_13 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_13; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_14 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_14; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_15 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_15; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_16 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_16; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_17 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_17; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_18 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_18; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_19 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_19; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_20 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_20; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_21 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_21; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_22 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_22; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_23 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_23; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_24 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_24; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_25 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_25; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_26 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_26; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_27 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_27; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_28 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_28; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_29 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_29; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_30 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_30; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_31 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_31; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_32 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_32; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_33 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_33; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_34 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_34; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_35 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_35; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_36 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_36; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_37 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_37; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_38 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_38; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_39 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_39; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_40 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_40; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_41 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_41; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_42 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_42; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_43 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_43; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_44 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_44; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_45 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_45; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_46 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_46; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_47 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_47; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_48 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_48; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_49 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_49; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_50 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_50; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_51 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_51; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_52 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_52; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_53 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_53; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_54 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_54; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_55 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_55; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_56 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_56; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_57 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_57; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_58 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_58; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_59 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_59; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_60 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_60; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_61 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_61; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_62 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_62; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_sram_id_table_63 = io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_63; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_0_mat_mod_table_mod_table_width; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_0_mat_mod_table_mod_table_depth; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_act_mod_en_0 = io_mod_proc_mod_0_act_mod_en_0; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_act_mod_en_1 = io_mod_proc_mod_0_act_mod_en_1; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_act_mod_addr = io_mod_proc_mod_0_act_mod_addr; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_act_mod_data_0 = io_mod_proc_mod_0_act_mod_data_0; // @[ipsa.scala 63:20]
  assign proc_0_io_mod_act_mod_data_1 = io_mod_proc_mod_0_act_mod_data_1; // @[ipsa.scala 63:20]
  assign proc_0_io_mem_cluster_0_data = sram_cluster_0_io_r_0_cluster_0_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_1_data = sram_cluster_0_io_r_0_cluster_1_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_2_data = sram_cluster_0_io_r_0_cluster_2_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_3_data = sram_cluster_0_io_r_0_cluster_3_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_4_data = sram_cluster_0_io_r_0_cluster_4_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_5_data = sram_cluster_0_io_r_0_cluster_5_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_6_data = sram_cluster_0_io_r_0_cluster_6_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_7_data = sram_cluster_0_io_r_0_cluster_7_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_8_data = sram_cluster_0_io_r_0_cluster_8_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_9_data = sram_cluster_0_io_r_0_cluster_9_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_10_data = sram_cluster_0_io_r_0_cluster_10_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_11_data = sram_cluster_0_io_r_0_cluster_11_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_12_data = sram_cluster_0_io_r_0_cluster_12_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_13_data = sram_cluster_0_io_r_0_cluster_13_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_14_data = sram_cluster_0_io_r_0_cluster_14_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_15_data = sram_cluster_0_io_r_0_cluster_15_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_16_data = sram_cluster_0_io_r_0_cluster_16_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_17_data = sram_cluster_0_io_r_0_cluster_17_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_18_data = sram_cluster_0_io_r_0_cluster_18_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_19_data = sram_cluster_0_io_r_0_cluster_19_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_20_data = sram_cluster_0_io_r_0_cluster_20_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_21_data = sram_cluster_0_io_r_0_cluster_21_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_22_data = sram_cluster_0_io_r_0_cluster_22_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_23_data = sram_cluster_0_io_r_0_cluster_23_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_24_data = sram_cluster_0_io_r_0_cluster_24_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_25_data = sram_cluster_0_io_r_0_cluster_25_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_26_data = sram_cluster_0_io_r_0_cluster_26_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_27_data = sram_cluster_0_io_r_0_cluster_27_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_28_data = sram_cluster_0_io_r_0_cluster_28_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_29_data = sram_cluster_0_io_r_0_cluster_29_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_30_data = sram_cluster_0_io_r_0_cluster_30_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_31_data = sram_cluster_0_io_r_0_cluster_31_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_32_data = sram_cluster_0_io_r_0_cluster_32_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_33_data = sram_cluster_0_io_r_0_cluster_33_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_34_data = sram_cluster_0_io_r_0_cluster_34_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_35_data = sram_cluster_0_io_r_0_cluster_35_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_36_data = sram_cluster_0_io_r_0_cluster_36_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_37_data = sram_cluster_0_io_r_0_cluster_37_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_38_data = sram_cluster_0_io_r_0_cluster_38_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_39_data = sram_cluster_0_io_r_0_cluster_39_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_40_data = sram_cluster_0_io_r_0_cluster_40_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_41_data = sram_cluster_0_io_r_0_cluster_41_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_42_data = sram_cluster_0_io_r_0_cluster_42_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_43_data = sram_cluster_0_io_r_0_cluster_43_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_44_data = sram_cluster_0_io_r_0_cluster_44_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_45_data = sram_cluster_0_io_r_0_cluster_45_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_46_data = sram_cluster_0_io_r_0_cluster_46_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_47_data = sram_cluster_0_io_r_0_cluster_47_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_48_data = sram_cluster_0_io_r_0_cluster_48_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_49_data = sram_cluster_0_io_r_0_cluster_49_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_50_data = sram_cluster_0_io_r_0_cluster_50_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_51_data = sram_cluster_0_io_r_0_cluster_51_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_52_data = sram_cluster_0_io_r_0_cluster_52_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_53_data = sram_cluster_0_io_r_0_cluster_53_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_54_data = sram_cluster_0_io_r_0_cluster_54_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_55_data = sram_cluster_0_io_r_0_cluster_55_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_56_data = sram_cluster_0_io_r_0_cluster_56_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_57_data = sram_cluster_0_io_r_0_cluster_57_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_58_data = sram_cluster_0_io_r_0_cluster_58_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_59_data = sram_cluster_0_io_r_0_cluster_59_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_60_data = sram_cluster_0_io_r_0_cluster_60_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_61_data = sram_cluster_0_io_r_0_cluster_61_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_62_data = sram_cluster_0_io_r_0_cluster_62_data; // @[ipsa.scala 76:37]
  assign proc_0_io_mem_cluster_63_data = sram_cluster_0_io_r_0_cluster_63_data; // @[ipsa.scala 76:37]
  assign proc_1_clock = clock;
  assign proc_1_io_pipe_phv_in_data_0 = recv_1_data_0; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_1 = recv_1_data_1; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_2 = recv_1_data_2; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_3 = recv_1_data_3; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_4 = recv_1_data_4; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_5 = recv_1_data_5; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_6 = recv_1_data_6; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_7 = recv_1_data_7; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_8 = recv_1_data_8; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_9 = recv_1_data_9; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_10 = recv_1_data_10; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_11 = recv_1_data_11; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_12 = recv_1_data_12; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_13 = recv_1_data_13; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_14 = recv_1_data_14; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_15 = recv_1_data_15; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_16 = recv_1_data_16; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_17 = recv_1_data_17; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_18 = recv_1_data_18; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_19 = recv_1_data_19; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_20 = recv_1_data_20; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_21 = recv_1_data_21; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_22 = recv_1_data_22; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_23 = recv_1_data_23; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_24 = recv_1_data_24; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_25 = recv_1_data_25; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_26 = recv_1_data_26; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_27 = recv_1_data_27; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_28 = recv_1_data_28; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_29 = recv_1_data_29; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_30 = recv_1_data_30; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_31 = recv_1_data_31; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_32 = recv_1_data_32; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_33 = recv_1_data_33; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_34 = recv_1_data_34; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_35 = recv_1_data_35; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_36 = recv_1_data_36; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_37 = recv_1_data_37; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_38 = recv_1_data_38; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_39 = recv_1_data_39; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_40 = recv_1_data_40; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_41 = recv_1_data_41; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_42 = recv_1_data_42; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_43 = recv_1_data_43; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_44 = recv_1_data_44; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_45 = recv_1_data_45; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_46 = recv_1_data_46; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_47 = recv_1_data_47; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_48 = recv_1_data_48; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_49 = recv_1_data_49; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_50 = recv_1_data_50; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_51 = recv_1_data_51; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_52 = recv_1_data_52; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_53 = recv_1_data_53; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_54 = recv_1_data_54; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_55 = recv_1_data_55; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_56 = recv_1_data_56; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_57 = recv_1_data_57; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_58 = recv_1_data_58; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_59 = recv_1_data_59; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_60 = recv_1_data_60; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_61 = recv_1_data_61; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_62 = recv_1_data_62; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_63 = recv_1_data_63; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_64 = recv_1_data_64; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_65 = recv_1_data_65; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_66 = recv_1_data_66; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_67 = recv_1_data_67; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_68 = recv_1_data_68; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_69 = recv_1_data_69; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_70 = recv_1_data_70; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_71 = recv_1_data_71; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_72 = recv_1_data_72; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_73 = recv_1_data_73; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_74 = recv_1_data_74; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_75 = recv_1_data_75; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_76 = recv_1_data_76; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_77 = recv_1_data_77; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_78 = recv_1_data_78; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_79 = recv_1_data_79; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_80 = recv_1_data_80; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_81 = recv_1_data_81; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_82 = recv_1_data_82; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_83 = recv_1_data_83; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_84 = recv_1_data_84; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_85 = recv_1_data_85; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_86 = recv_1_data_86; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_87 = recv_1_data_87; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_88 = recv_1_data_88; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_89 = recv_1_data_89; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_90 = recv_1_data_90; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_91 = recv_1_data_91; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_92 = recv_1_data_92; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_93 = recv_1_data_93; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_94 = recv_1_data_94; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_95 = recv_1_data_95; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_96 = recv_1_data_96; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_97 = recv_1_data_97; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_98 = recv_1_data_98; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_99 = recv_1_data_99; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_100 = recv_1_data_100; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_101 = recv_1_data_101; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_102 = recv_1_data_102; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_103 = recv_1_data_103; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_104 = recv_1_data_104; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_105 = recv_1_data_105; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_106 = recv_1_data_106; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_107 = recv_1_data_107; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_108 = recv_1_data_108; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_109 = recv_1_data_109; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_110 = recv_1_data_110; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_111 = recv_1_data_111; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_112 = recv_1_data_112; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_113 = recv_1_data_113; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_114 = recv_1_data_114; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_115 = recv_1_data_115; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_116 = recv_1_data_116; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_117 = recv_1_data_117; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_118 = recv_1_data_118; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_119 = recv_1_data_119; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_120 = recv_1_data_120; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_121 = recv_1_data_121; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_122 = recv_1_data_122; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_123 = recv_1_data_123; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_124 = recv_1_data_124; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_125 = recv_1_data_125; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_126 = recv_1_data_126; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_127 = recv_1_data_127; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_128 = recv_1_data_128; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_129 = recv_1_data_129; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_130 = recv_1_data_130; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_131 = recv_1_data_131; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_132 = recv_1_data_132; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_133 = recv_1_data_133; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_134 = recv_1_data_134; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_135 = recv_1_data_135; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_136 = recv_1_data_136; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_137 = recv_1_data_137; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_138 = recv_1_data_138; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_139 = recv_1_data_139; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_140 = recv_1_data_140; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_141 = recv_1_data_141; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_142 = recv_1_data_142; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_143 = recv_1_data_143; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_144 = recv_1_data_144; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_145 = recv_1_data_145; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_146 = recv_1_data_146; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_147 = recv_1_data_147; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_148 = recv_1_data_148; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_149 = recv_1_data_149; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_150 = recv_1_data_150; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_151 = recv_1_data_151; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_152 = recv_1_data_152; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_153 = recv_1_data_153; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_154 = recv_1_data_154; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_155 = recv_1_data_155; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_156 = recv_1_data_156; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_157 = recv_1_data_157; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_158 = recv_1_data_158; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_159 = recv_1_data_159; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_160 = recv_1_data_160; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_161 = recv_1_data_161; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_162 = recv_1_data_162; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_163 = recv_1_data_163; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_164 = recv_1_data_164; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_165 = recv_1_data_165; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_166 = recv_1_data_166; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_167 = recv_1_data_167; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_168 = recv_1_data_168; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_169 = recv_1_data_169; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_170 = recv_1_data_170; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_171 = recv_1_data_171; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_172 = recv_1_data_172; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_173 = recv_1_data_173; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_174 = recv_1_data_174; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_175 = recv_1_data_175; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_176 = recv_1_data_176; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_177 = recv_1_data_177; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_178 = recv_1_data_178; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_179 = recv_1_data_179; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_180 = recv_1_data_180; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_181 = recv_1_data_181; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_182 = recv_1_data_182; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_183 = recv_1_data_183; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_184 = recv_1_data_184; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_185 = recv_1_data_185; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_186 = recv_1_data_186; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_187 = recv_1_data_187; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_188 = recv_1_data_188; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_189 = recv_1_data_189; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_190 = recv_1_data_190; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_191 = recv_1_data_191; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_192 = recv_1_data_192; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_193 = recv_1_data_193; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_194 = recv_1_data_194; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_195 = recv_1_data_195; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_196 = recv_1_data_196; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_197 = recv_1_data_197; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_198 = recv_1_data_198; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_199 = recv_1_data_199; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_200 = recv_1_data_200; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_201 = recv_1_data_201; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_202 = recv_1_data_202; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_203 = recv_1_data_203; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_204 = recv_1_data_204; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_205 = recv_1_data_205; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_206 = recv_1_data_206; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_207 = recv_1_data_207; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_208 = recv_1_data_208; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_209 = recv_1_data_209; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_210 = recv_1_data_210; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_211 = recv_1_data_211; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_212 = recv_1_data_212; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_213 = recv_1_data_213; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_214 = recv_1_data_214; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_215 = recv_1_data_215; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_216 = recv_1_data_216; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_217 = recv_1_data_217; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_218 = recv_1_data_218; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_219 = recv_1_data_219; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_220 = recv_1_data_220; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_221 = recv_1_data_221; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_222 = recv_1_data_222; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_223 = recv_1_data_223; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_224 = recv_1_data_224; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_225 = recv_1_data_225; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_226 = recv_1_data_226; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_227 = recv_1_data_227; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_228 = recv_1_data_228; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_229 = recv_1_data_229; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_230 = recv_1_data_230; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_231 = recv_1_data_231; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_232 = recv_1_data_232; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_233 = recv_1_data_233; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_234 = recv_1_data_234; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_235 = recv_1_data_235; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_236 = recv_1_data_236; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_237 = recv_1_data_237; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_238 = recv_1_data_238; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_239 = recv_1_data_239; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_240 = recv_1_data_240; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_241 = recv_1_data_241; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_242 = recv_1_data_242; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_243 = recv_1_data_243; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_244 = recv_1_data_244; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_245 = recv_1_data_245; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_246 = recv_1_data_246; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_247 = recv_1_data_247; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_248 = recv_1_data_248; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_249 = recv_1_data_249; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_250 = recv_1_data_250; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_251 = recv_1_data_251; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_252 = recv_1_data_252; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_253 = recv_1_data_253; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_254 = recv_1_data_254; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_data_255 = recv_1_data_255; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_header_0 = recv_1_header_0; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_header_1 = recv_1_header_1; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_header_2 = recv_1_header_2; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_header_3 = recv_1_header_3; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_header_4 = recv_1_header_4; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_header_5 = recv_1_header_5; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_header_6 = recv_1_header_6; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_header_7 = recv_1_header_7; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_header_8 = recv_1_header_8; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_header_9 = recv_1_header_9; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_header_10 = recv_1_header_10; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_header_11 = recv_1_header_11; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_header_12 = recv_1_header_12; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_header_13 = recv_1_header_13; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_header_14 = recv_1_header_14; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_header_15 = recv_1_header_15; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_parse_current_state = recv_1_parse_current_state; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_parse_current_offset = recv_1_parse_current_offset; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_parse_transition_field = recv_1_parse_transition_field; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_next_processor_id = recv_1_next_processor_id; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_next_config_id = recv_1_next_config_id; // @[ipsa.scala 161:32]
  assign proc_1_io_pipe_phv_in_is_valid_processor = recv_1_is_valid_processor; // @[ipsa.scala 161:32]
  assign proc_1_io_mod_par_mod_en = io_mod_proc_mod_1_par_mod_en; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_par_mod_last_mau_id_mod = io_mod_proc_mod_1_par_mod_last_mau_id_mod; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_par_mod_last_mau_id = io_mod_proc_mod_1_par_mod_last_mau_id; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_par_mod_cs = io_mod_proc_mod_1_par_mod_cs; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_par_mod_module_mod_state_id_mod = io_mod_proc_mod_1_par_mod_module_mod_state_id_mod; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_par_mod_module_mod_state_id = io_mod_proc_mod_1_par_mod_module_mod_state_id; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_par_mod_module_mod_sram_w_cs = io_mod_proc_mod_1_par_mod_module_mod_sram_w_cs; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_par_mod_module_mod_sram_w_en = io_mod_proc_mod_1_par_mod_module_mod_sram_w_en; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_par_mod_module_mod_sram_w_addr = io_mod_proc_mod_1_par_mod_module_mod_sram_w_addr; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_par_mod_module_mod_sram_w_data = io_mod_proc_mod_1_par_mod_module_mod_sram_w_data; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_en = io_mod_proc_mod_1_mat_mod_en; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_config_id = io_mod_proc_mod_1_mat_mod_config_id; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_key_mod_header_id = io_mod_proc_mod_1_mat_mod_key_mod_header_id; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_key_mod_internal_offset = io_mod_proc_mod_1_mat_mod_key_mod_internal_offset; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_key_mod_key_length = io_mod_proc_mod_1_mat_mod_key_mod_key_length; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_0 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_0; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_1 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_1; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_2 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_2; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_3 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_3; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_4 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_4; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_5 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_5; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_6 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_6; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_7 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_7; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_8 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_8; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_9 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_9; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_10 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_10; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_11 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_11; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_12 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_12; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_13 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_13; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_14 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_14; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_15 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_15; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_16 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_16; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_17 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_17; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_18 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_18; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_19 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_19; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_20 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_20; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_21 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_21; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_22 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_22; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_23 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_23; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_24 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_24; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_25 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_25; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_26 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_26; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_27 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_27; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_28 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_28; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_29 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_29; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_30 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_30; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_31 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_31; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_32 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_32; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_33 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_33; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_34 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_34; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_35 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_35; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_36 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_36; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_37 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_37; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_38 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_38; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_39 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_39; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_40 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_40; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_41 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_41; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_42 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_42; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_43 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_43; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_44 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_44; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_45 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_45; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_46 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_46; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_47 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_47; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_48 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_48; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_49 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_49; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_50 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_50; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_51 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_51; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_52 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_52; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_53 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_53; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_54 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_54; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_55 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_55; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_56 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_56; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_57 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_57; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_58 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_58; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_59 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_59; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_60 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_60; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_61 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_61; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_62 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_62; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_sram_id_table_63 = io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_63; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_1_mat_mod_table_mod_table_width; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_1_mat_mod_table_mod_table_depth; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_act_mod_en_0 = io_mod_proc_mod_1_act_mod_en_0; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_act_mod_en_1 = io_mod_proc_mod_1_act_mod_en_1; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_act_mod_addr = io_mod_proc_mod_1_act_mod_addr; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_act_mod_data_0 = io_mod_proc_mod_1_act_mod_data_0; // @[ipsa.scala 63:20]
  assign proc_1_io_mod_act_mod_data_1 = io_mod_proc_mod_1_act_mod_data_1; // @[ipsa.scala 63:20]
  assign proc_1_io_mem_cluster_0_data = sram_cluster_0_io_r_1_cluster_0_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_1_data = sram_cluster_0_io_r_1_cluster_1_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_2_data = sram_cluster_0_io_r_1_cluster_2_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_3_data = sram_cluster_0_io_r_1_cluster_3_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_4_data = sram_cluster_0_io_r_1_cluster_4_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_5_data = sram_cluster_0_io_r_1_cluster_5_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_6_data = sram_cluster_0_io_r_1_cluster_6_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_7_data = sram_cluster_0_io_r_1_cluster_7_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_8_data = sram_cluster_0_io_r_1_cluster_8_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_9_data = sram_cluster_0_io_r_1_cluster_9_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_10_data = sram_cluster_0_io_r_1_cluster_10_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_11_data = sram_cluster_0_io_r_1_cluster_11_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_12_data = sram_cluster_0_io_r_1_cluster_12_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_13_data = sram_cluster_0_io_r_1_cluster_13_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_14_data = sram_cluster_0_io_r_1_cluster_14_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_15_data = sram_cluster_0_io_r_1_cluster_15_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_16_data = sram_cluster_0_io_r_1_cluster_16_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_17_data = sram_cluster_0_io_r_1_cluster_17_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_18_data = sram_cluster_0_io_r_1_cluster_18_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_19_data = sram_cluster_0_io_r_1_cluster_19_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_20_data = sram_cluster_0_io_r_1_cluster_20_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_21_data = sram_cluster_0_io_r_1_cluster_21_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_22_data = sram_cluster_0_io_r_1_cluster_22_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_23_data = sram_cluster_0_io_r_1_cluster_23_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_24_data = sram_cluster_0_io_r_1_cluster_24_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_25_data = sram_cluster_0_io_r_1_cluster_25_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_26_data = sram_cluster_0_io_r_1_cluster_26_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_27_data = sram_cluster_0_io_r_1_cluster_27_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_28_data = sram_cluster_0_io_r_1_cluster_28_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_29_data = sram_cluster_0_io_r_1_cluster_29_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_30_data = sram_cluster_0_io_r_1_cluster_30_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_31_data = sram_cluster_0_io_r_1_cluster_31_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_32_data = sram_cluster_0_io_r_1_cluster_32_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_33_data = sram_cluster_0_io_r_1_cluster_33_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_34_data = sram_cluster_0_io_r_1_cluster_34_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_35_data = sram_cluster_0_io_r_1_cluster_35_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_36_data = sram_cluster_0_io_r_1_cluster_36_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_37_data = sram_cluster_0_io_r_1_cluster_37_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_38_data = sram_cluster_0_io_r_1_cluster_38_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_39_data = sram_cluster_0_io_r_1_cluster_39_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_40_data = sram_cluster_0_io_r_1_cluster_40_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_41_data = sram_cluster_0_io_r_1_cluster_41_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_42_data = sram_cluster_0_io_r_1_cluster_42_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_43_data = sram_cluster_0_io_r_1_cluster_43_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_44_data = sram_cluster_0_io_r_1_cluster_44_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_45_data = sram_cluster_0_io_r_1_cluster_45_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_46_data = sram_cluster_0_io_r_1_cluster_46_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_47_data = sram_cluster_0_io_r_1_cluster_47_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_48_data = sram_cluster_0_io_r_1_cluster_48_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_49_data = sram_cluster_0_io_r_1_cluster_49_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_50_data = sram_cluster_0_io_r_1_cluster_50_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_51_data = sram_cluster_0_io_r_1_cluster_51_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_52_data = sram_cluster_0_io_r_1_cluster_52_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_53_data = sram_cluster_0_io_r_1_cluster_53_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_54_data = sram_cluster_0_io_r_1_cluster_54_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_55_data = sram_cluster_0_io_r_1_cluster_55_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_56_data = sram_cluster_0_io_r_1_cluster_56_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_57_data = sram_cluster_0_io_r_1_cluster_57_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_58_data = sram_cluster_0_io_r_1_cluster_58_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_59_data = sram_cluster_0_io_r_1_cluster_59_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_60_data = sram_cluster_0_io_r_1_cluster_60_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_61_data = sram_cluster_0_io_r_1_cluster_61_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_62_data = sram_cluster_0_io_r_1_cluster_62_data; // @[ipsa.scala 76:37]
  assign proc_1_io_mem_cluster_63_data = sram_cluster_0_io_r_1_cluster_63_data; // @[ipsa.scala 76:37]
  assign proc_2_clock = clock;
  assign proc_2_io_pipe_phv_in_data_0 = recv_2_data_0; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_1 = recv_2_data_1; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_2 = recv_2_data_2; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_3 = recv_2_data_3; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_4 = recv_2_data_4; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_5 = recv_2_data_5; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_6 = recv_2_data_6; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_7 = recv_2_data_7; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_8 = recv_2_data_8; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_9 = recv_2_data_9; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_10 = recv_2_data_10; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_11 = recv_2_data_11; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_12 = recv_2_data_12; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_13 = recv_2_data_13; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_14 = recv_2_data_14; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_15 = recv_2_data_15; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_16 = recv_2_data_16; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_17 = recv_2_data_17; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_18 = recv_2_data_18; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_19 = recv_2_data_19; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_20 = recv_2_data_20; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_21 = recv_2_data_21; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_22 = recv_2_data_22; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_23 = recv_2_data_23; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_24 = recv_2_data_24; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_25 = recv_2_data_25; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_26 = recv_2_data_26; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_27 = recv_2_data_27; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_28 = recv_2_data_28; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_29 = recv_2_data_29; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_30 = recv_2_data_30; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_31 = recv_2_data_31; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_32 = recv_2_data_32; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_33 = recv_2_data_33; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_34 = recv_2_data_34; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_35 = recv_2_data_35; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_36 = recv_2_data_36; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_37 = recv_2_data_37; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_38 = recv_2_data_38; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_39 = recv_2_data_39; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_40 = recv_2_data_40; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_41 = recv_2_data_41; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_42 = recv_2_data_42; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_43 = recv_2_data_43; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_44 = recv_2_data_44; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_45 = recv_2_data_45; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_46 = recv_2_data_46; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_47 = recv_2_data_47; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_48 = recv_2_data_48; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_49 = recv_2_data_49; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_50 = recv_2_data_50; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_51 = recv_2_data_51; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_52 = recv_2_data_52; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_53 = recv_2_data_53; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_54 = recv_2_data_54; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_55 = recv_2_data_55; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_56 = recv_2_data_56; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_57 = recv_2_data_57; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_58 = recv_2_data_58; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_59 = recv_2_data_59; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_60 = recv_2_data_60; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_61 = recv_2_data_61; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_62 = recv_2_data_62; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_63 = recv_2_data_63; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_64 = recv_2_data_64; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_65 = recv_2_data_65; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_66 = recv_2_data_66; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_67 = recv_2_data_67; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_68 = recv_2_data_68; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_69 = recv_2_data_69; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_70 = recv_2_data_70; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_71 = recv_2_data_71; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_72 = recv_2_data_72; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_73 = recv_2_data_73; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_74 = recv_2_data_74; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_75 = recv_2_data_75; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_76 = recv_2_data_76; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_77 = recv_2_data_77; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_78 = recv_2_data_78; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_79 = recv_2_data_79; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_80 = recv_2_data_80; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_81 = recv_2_data_81; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_82 = recv_2_data_82; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_83 = recv_2_data_83; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_84 = recv_2_data_84; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_85 = recv_2_data_85; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_86 = recv_2_data_86; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_87 = recv_2_data_87; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_88 = recv_2_data_88; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_89 = recv_2_data_89; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_90 = recv_2_data_90; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_91 = recv_2_data_91; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_92 = recv_2_data_92; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_93 = recv_2_data_93; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_94 = recv_2_data_94; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_95 = recv_2_data_95; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_96 = recv_2_data_96; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_97 = recv_2_data_97; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_98 = recv_2_data_98; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_99 = recv_2_data_99; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_100 = recv_2_data_100; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_101 = recv_2_data_101; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_102 = recv_2_data_102; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_103 = recv_2_data_103; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_104 = recv_2_data_104; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_105 = recv_2_data_105; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_106 = recv_2_data_106; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_107 = recv_2_data_107; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_108 = recv_2_data_108; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_109 = recv_2_data_109; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_110 = recv_2_data_110; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_111 = recv_2_data_111; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_112 = recv_2_data_112; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_113 = recv_2_data_113; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_114 = recv_2_data_114; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_115 = recv_2_data_115; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_116 = recv_2_data_116; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_117 = recv_2_data_117; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_118 = recv_2_data_118; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_119 = recv_2_data_119; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_120 = recv_2_data_120; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_121 = recv_2_data_121; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_122 = recv_2_data_122; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_123 = recv_2_data_123; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_124 = recv_2_data_124; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_125 = recv_2_data_125; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_126 = recv_2_data_126; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_127 = recv_2_data_127; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_128 = recv_2_data_128; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_129 = recv_2_data_129; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_130 = recv_2_data_130; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_131 = recv_2_data_131; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_132 = recv_2_data_132; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_133 = recv_2_data_133; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_134 = recv_2_data_134; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_135 = recv_2_data_135; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_136 = recv_2_data_136; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_137 = recv_2_data_137; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_138 = recv_2_data_138; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_139 = recv_2_data_139; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_140 = recv_2_data_140; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_141 = recv_2_data_141; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_142 = recv_2_data_142; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_143 = recv_2_data_143; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_144 = recv_2_data_144; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_145 = recv_2_data_145; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_146 = recv_2_data_146; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_147 = recv_2_data_147; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_148 = recv_2_data_148; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_149 = recv_2_data_149; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_150 = recv_2_data_150; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_151 = recv_2_data_151; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_152 = recv_2_data_152; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_153 = recv_2_data_153; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_154 = recv_2_data_154; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_155 = recv_2_data_155; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_156 = recv_2_data_156; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_157 = recv_2_data_157; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_158 = recv_2_data_158; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_159 = recv_2_data_159; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_160 = recv_2_data_160; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_161 = recv_2_data_161; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_162 = recv_2_data_162; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_163 = recv_2_data_163; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_164 = recv_2_data_164; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_165 = recv_2_data_165; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_166 = recv_2_data_166; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_167 = recv_2_data_167; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_168 = recv_2_data_168; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_169 = recv_2_data_169; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_170 = recv_2_data_170; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_171 = recv_2_data_171; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_172 = recv_2_data_172; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_173 = recv_2_data_173; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_174 = recv_2_data_174; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_175 = recv_2_data_175; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_176 = recv_2_data_176; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_177 = recv_2_data_177; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_178 = recv_2_data_178; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_179 = recv_2_data_179; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_180 = recv_2_data_180; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_181 = recv_2_data_181; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_182 = recv_2_data_182; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_183 = recv_2_data_183; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_184 = recv_2_data_184; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_185 = recv_2_data_185; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_186 = recv_2_data_186; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_187 = recv_2_data_187; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_188 = recv_2_data_188; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_189 = recv_2_data_189; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_190 = recv_2_data_190; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_191 = recv_2_data_191; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_192 = recv_2_data_192; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_193 = recv_2_data_193; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_194 = recv_2_data_194; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_195 = recv_2_data_195; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_196 = recv_2_data_196; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_197 = recv_2_data_197; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_198 = recv_2_data_198; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_199 = recv_2_data_199; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_200 = recv_2_data_200; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_201 = recv_2_data_201; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_202 = recv_2_data_202; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_203 = recv_2_data_203; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_204 = recv_2_data_204; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_205 = recv_2_data_205; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_206 = recv_2_data_206; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_207 = recv_2_data_207; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_208 = recv_2_data_208; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_209 = recv_2_data_209; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_210 = recv_2_data_210; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_211 = recv_2_data_211; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_212 = recv_2_data_212; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_213 = recv_2_data_213; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_214 = recv_2_data_214; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_215 = recv_2_data_215; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_216 = recv_2_data_216; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_217 = recv_2_data_217; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_218 = recv_2_data_218; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_219 = recv_2_data_219; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_220 = recv_2_data_220; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_221 = recv_2_data_221; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_222 = recv_2_data_222; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_223 = recv_2_data_223; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_224 = recv_2_data_224; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_225 = recv_2_data_225; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_226 = recv_2_data_226; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_227 = recv_2_data_227; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_228 = recv_2_data_228; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_229 = recv_2_data_229; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_230 = recv_2_data_230; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_231 = recv_2_data_231; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_232 = recv_2_data_232; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_233 = recv_2_data_233; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_234 = recv_2_data_234; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_235 = recv_2_data_235; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_236 = recv_2_data_236; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_237 = recv_2_data_237; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_238 = recv_2_data_238; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_239 = recv_2_data_239; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_240 = recv_2_data_240; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_241 = recv_2_data_241; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_242 = recv_2_data_242; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_243 = recv_2_data_243; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_244 = recv_2_data_244; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_245 = recv_2_data_245; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_246 = recv_2_data_246; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_247 = recv_2_data_247; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_248 = recv_2_data_248; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_249 = recv_2_data_249; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_250 = recv_2_data_250; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_251 = recv_2_data_251; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_252 = recv_2_data_252; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_253 = recv_2_data_253; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_254 = recv_2_data_254; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_data_255 = recv_2_data_255; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_header_0 = recv_2_header_0; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_header_1 = recv_2_header_1; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_header_2 = recv_2_header_2; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_header_3 = recv_2_header_3; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_header_4 = recv_2_header_4; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_header_5 = recv_2_header_5; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_header_6 = recv_2_header_6; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_header_7 = recv_2_header_7; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_header_8 = recv_2_header_8; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_header_9 = recv_2_header_9; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_header_10 = recv_2_header_10; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_header_11 = recv_2_header_11; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_header_12 = recv_2_header_12; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_header_13 = recv_2_header_13; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_header_14 = recv_2_header_14; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_header_15 = recv_2_header_15; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_parse_current_state = recv_2_parse_current_state; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_parse_current_offset = recv_2_parse_current_offset; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_parse_transition_field = recv_2_parse_transition_field; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_next_processor_id = recv_2_next_processor_id; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_next_config_id = recv_2_next_config_id; // @[ipsa.scala 161:32]
  assign proc_2_io_pipe_phv_in_is_valid_processor = recv_2_is_valid_processor; // @[ipsa.scala 161:32]
  assign proc_2_io_mod_par_mod_en = io_mod_proc_mod_2_par_mod_en; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_par_mod_last_mau_id_mod = io_mod_proc_mod_2_par_mod_last_mau_id_mod; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_par_mod_last_mau_id = io_mod_proc_mod_2_par_mod_last_mau_id; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_par_mod_cs = io_mod_proc_mod_2_par_mod_cs; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_par_mod_module_mod_state_id_mod = io_mod_proc_mod_2_par_mod_module_mod_state_id_mod; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_par_mod_module_mod_state_id = io_mod_proc_mod_2_par_mod_module_mod_state_id; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_par_mod_module_mod_sram_w_cs = io_mod_proc_mod_2_par_mod_module_mod_sram_w_cs; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_par_mod_module_mod_sram_w_en = io_mod_proc_mod_2_par_mod_module_mod_sram_w_en; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_par_mod_module_mod_sram_w_addr = io_mod_proc_mod_2_par_mod_module_mod_sram_w_addr; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_par_mod_module_mod_sram_w_data = io_mod_proc_mod_2_par_mod_module_mod_sram_w_data; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_en = io_mod_proc_mod_2_mat_mod_en; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_config_id = io_mod_proc_mod_2_mat_mod_config_id; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_key_mod_header_id = io_mod_proc_mod_2_mat_mod_key_mod_header_id; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_key_mod_internal_offset = io_mod_proc_mod_2_mat_mod_key_mod_internal_offset; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_key_mod_key_length = io_mod_proc_mod_2_mat_mod_key_mod_key_length; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_0 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_0; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_1 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_1; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_2 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_2; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_3 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_3; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_4 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_4; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_5 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_5; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_6 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_6; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_7 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_7; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_8 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_8; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_9 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_9; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_10 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_10; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_11 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_11; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_12 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_12; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_13 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_13; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_14 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_14; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_15 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_15; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_16 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_16; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_17 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_17; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_18 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_18; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_19 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_19; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_20 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_20; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_21 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_21; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_22 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_22; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_23 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_23; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_24 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_24; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_25 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_25; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_26 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_26; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_27 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_27; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_28 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_28; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_29 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_29; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_30 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_30; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_31 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_31; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_32 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_32; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_33 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_33; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_34 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_34; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_35 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_35; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_36 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_36; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_37 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_37; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_38 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_38; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_39 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_39; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_40 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_40; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_41 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_41; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_42 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_42; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_43 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_43; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_44 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_44; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_45 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_45; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_46 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_46; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_47 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_47; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_48 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_48; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_49 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_49; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_50 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_50; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_51 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_51; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_52 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_52; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_53 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_53; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_54 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_54; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_55 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_55; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_56 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_56; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_57 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_57; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_58 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_58; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_59 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_59; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_60 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_60; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_61 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_61; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_62 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_62; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_sram_id_table_63 = io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_63; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_2_mat_mod_table_mod_table_width; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_2_mat_mod_table_mod_table_depth; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_act_mod_en_0 = io_mod_proc_mod_2_act_mod_en_0; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_act_mod_en_1 = io_mod_proc_mod_2_act_mod_en_1; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_act_mod_addr = io_mod_proc_mod_2_act_mod_addr; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_act_mod_data_0 = io_mod_proc_mod_2_act_mod_data_0; // @[ipsa.scala 63:20]
  assign proc_2_io_mod_act_mod_data_1 = io_mod_proc_mod_2_act_mod_data_1; // @[ipsa.scala 63:20]
  assign proc_2_io_mem_cluster_0_data = sram_cluster_0_io_r_2_cluster_0_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_1_data = sram_cluster_0_io_r_2_cluster_1_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_2_data = sram_cluster_0_io_r_2_cluster_2_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_3_data = sram_cluster_0_io_r_2_cluster_3_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_4_data = sram_cluster_0_io_r_2_cluster_4_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_5_data = sram_cluster_0_io_r_2_cluster_5_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_6_data = sram_cluster_0_io_r_2_cluster_6_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_7_data = sram_cluster_0_io_r_2_cluster_7_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_8_data = sram_cluster_0_io_r_2_cluster_8_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_9_data = sram_cluster_0_io_r_2_cluster_9_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_10_data = sram_cluster_0_io_r_2_cluster_10_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_11_data = sram_cluster_0_io_r_2_cluster_11_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_12_data = sram_cluster_0_io_r_2_cluster_12_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_13_data = sram_cluster_0_io_r_2_cluster_13_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_14_data = sram_cluster_0_io_r_2_cluster_14_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_15_data = sram_cluster_0_io_r_2_cluster_15_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_16_data = sram_cluster_0_io_r_2_cluster_16_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_17_data = sram_cluster_0_io_r_2_cluster_17_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_18_data = sram_cluster_0_io_r_2_cluster_18_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_19_data = sram_cluster_0_io_r_2_cluster_19_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_20_data = sram_cluster_0_io_r_2_cluster_20_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_21_data = sram_cluster_0_io_r_2_cluster_21_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_22_data = sram_cluster_0_io_r_2_cluster_22_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_23_data = sram_cluster_0_io_r_2_cluster_23_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_24_data = sram_cluster_0_io_r_2_cluster_24_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_25_data = sram_cluster_0_io_r_2_cluster_25_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_26_data = sram_cluster_0_io_r_2_cluster_26_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_27_data = sram_cluster_0_io_r_2_cluster_27_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_28_data = sram_cluster_0_io_r_2_cluster_28_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_29_data = sram_cluster_0_io_r_2_cluster_29_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_30_data = sram_cluster_0_io_r_2_cluster_30_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_31_data = sram_cluster_0_io_r_2_cluster_31_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_32_data = sram_cluster_0_io_r_2_cluster_32_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_33_data = sram_cluster_0_io_r_2_cluster_33_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_34_data = sram_cluster_0_io_r_2_cluster_34_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_35_data = sram_cluster_0_io_r_2_cluster_35_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_36_data = sram_cluster_0_io_r_2_cluster_36_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_37_data = sram_cluster_0_io_r_2_cluster_37_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_38_data = sram_cluster_0_io_r_2_cluster_38_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_39_data = sram_cluster_0_io_r_2_cluster_39_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_40_data = sram_cluster_0_io_r_2_cluster_40_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_41_data = sram_cluster_0_io_r_2_cluster_41_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_42_data = sram_cluster_0_io_r_2_cluster_42_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_43_data = sram_cluster_0_io_r_2_cluster_43_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_44_data = sram_cluster_0_io_r_2_cluster_44_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_45_data = sram_cluster_0_io_r_2_cluster_45_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_46_data = sram_cluster_0_io_r_2_cluster_46_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_47_data = sram_cluster_0_io_r_2_cluster_47_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_48_data = sram_cluster_0_io_r_2_cluster_48_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_49_data = sram_cluster_0_io_r_2_cluster_49_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_50_data = sram_cluster_0_io_r_2_cluster_50_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_51_data = sram_cluster_0_io_r_2_cluster_51_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_52_data = sram_cluster_0_io_r_2_cluster_52_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_53_data = sram_cluster_0_io_r_2_cluster_53_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_54_data = sram_cluster_0_io_r_2_cluster_54_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_55_data = sram_cluster_0_io_r_2_cluster_55_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_56_data = sram_cluster_0_io_r_2_cluster_56_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_57_data = sram_cluster_0_io_r_2_cluster_57_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_58_data = sram_cluster_0_io_r_2_cluster_58_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_59_data = sram_cluster_0_io_r_2_cluster_59_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_60_data = sram_cluster_0_io_r_2_cluster_60_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_61_data = sram_cluster_0_io_r_2_cluster_61_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_62_data = sram_cluster_0_io_r_2_cluster_62_data; // @[ipsa.scala 76:37]
  assign proc_2_io_mem_cluster_63_data = sram_cluster_0_io_r_2_cluster_63_data; // @[ipsa.scala 76:37]
  assign proc_3_clock = clock;
  assign proc_3_io_pipe_phv_in_data_0 = recv_3_data_0; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_1 = recv_3_data_1; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_2 = recv_3_data_2; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_3 = recv_3_data_3; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_4 = recv_3_data_4; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_5 = recv_3_data_5; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_6 = recv_3_data_6; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_7 = recv_3_data_7; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_8 = recv_3_data_8; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_9 = recv_3_data_9; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_10 = recv_3_data_10; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_11 = recv_3_data_11; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_12 = recv_3_data_12; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_13 = recv_3_data_13; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_14 = recv_3_data_14; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_15 = recv_3_data_15; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_16 = recv_3_data_16; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_17 = recv_3_data_17; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_18 = recv_3_data_18; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_19 = recv_3_data_19; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_20 = recv_3_data_20; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_21 = recv_3_data_21; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_22 = recv_3_data_22; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_23 = recv_3_data_23; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_24 = recv_3_data_24; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_25 = recv_3_data_25; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_26 = recv_3_data_26; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_27 = recv_3_data_27; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_28 = recv_3_data_28; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_29 = recv_3_data_29; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_30 = recv_3_data_30; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_31 = recv_3_data_31; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_32 = recv_3_data_32; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_33 = recv_3_data_33; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_34 = recv_3_data_34; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_35 = recv_3_data_35; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_36 = recv_3_data_36; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_37 = recv_3_data_37; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_38 = recv_3_data_38; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_39 = recv_3_data_39; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_40 = recv_3_data_40; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_41 = recv_3_data_41; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_42 = recv_3_data_42; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_43 = recv_3_data_43; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_44 = recv_3_data_44; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_45 = recv_3_data_45; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_46 = recv_3_data_46; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_47 = recv_3_data_47; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_48 = recv_3_data_48; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_49 = recv_3_data_49; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_50 = recv_3_data_50; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_51 = recv_3_data_51; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_52 = recv_3_data_52; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_53 = recv_3_data_53; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_54 = recv_3_data_54; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_55 = recv_3_data_55; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_56 = recv_3_data_56; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_57 = recv_3_data_57; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_58 = recv_3_data_58; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_59 = recv_3_data_59; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_60 = recv_3_data_60; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_61 = recv_3_data_61; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_62 = recv_3_data_62; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_63 = recv_3_data_63; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_64 = recv_3_data_64; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_65 = recv_3_data_65; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_66 = recv_3_data_66; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_67 = recv_3_data_67; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_68 = recv_3_data_68; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_69 = recv_3_data_69; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_70 = recv_3_data_70; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_71 = recv_3_data_71; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_72 = recv_3_data_72; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_73 = recv_3_data_73; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_74 = recv_3_data_74; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_75 = recv_3_data_75; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_76 = recv_3_data_76; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_77 = recv_3_data_77; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_78 = recv_3_data_78; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_79 = recv_3_data_79; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_80 = recv_3_data_80; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_81 = recv_3_data_81; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_82 = recv_3_data_82; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_83 = recv_3_data_83; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_84 = recv_3_data_84; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_85 = recv_3_data_85; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_86 = recv_3_data_86; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_87 = recv_3_data_87; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_88 = recv_3_data_88; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_89 = recv_3_data_89; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_90 = recv_3_data_90; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_91 = recv_3_data_91; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_92 = recv_3_data_92; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_93 = recv_3_data_93; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_94 = recv_3_data_94; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_95 = recv_3_data_95; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_96 = recv_3_data_96; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_97 = recv_3_data_97; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_98 = recv_3_data_98; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_99 = recv_3_data_99; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_100 = recv_3_data_100; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_101 = recv_3_data_101; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_102 = recv_3_data_102; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_103 = recv_3_data_103; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_104 = recv_3_data_104; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_105 = recv_3_data_105; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_106 = recv_3_data_106; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_107 = recv_3_data_107; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_108 = recv_3_data_108; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_109 = recv_3_data_109; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_110 = recv_3_data_110; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_111 = recv_3_data_111; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_112 = recv_3_data_112; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_113 = recv_3_data_113; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_114 = recv_3_data_114; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_115 = recv_3_data_115; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_116 = recv_3_data_116; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_117 = recv_3_data_117; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_118 = recv_3_data_118; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_119 = recv_3_data_119; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_120 = recv_3_data_120; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_121 = recv_3_data_121; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_122 = recv_3_data_122; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_123 = recv_3_data_123; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_124 = recv_3_data_124; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_125 = recv_3_data_125; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_126 = recv_3_data_126; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_127 = recv_3_data_127; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_128 = recv_3_data_128; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_129 = recv_3_data_129; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_130 = recv_3_data_130; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_131 = recv_3_data_131; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_132 = recv_3_data_132; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_133 = recv_3_data_133; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_134 = recv_3_data_134; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_135 = recv_3_data_135; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_136 = recv_3_data_136; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_137 = recv_3_data_137; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_138 = recv_3_data_138; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_139 = recv_3_data_139; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_140 = recv_3_data_140; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_141 = recv_3_data_141; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_142 = recv_3_data_142; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_143 = recv_3_data_143; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_144 = recv_3_data_144; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_145 = recv_3_data_145; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_146 = recv_3_data_146; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_147 = recv_3_data_147; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_148 = recv_3_data_148; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_149 = recv_3_data_149; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_150 = recv_3_data_150; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_151 = recv_3_data_151; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_152 = recv_3_data_152; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_153 = recv_3_data_153; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_154 = recv_3_data_154; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_155 = recv_3_data_155; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_156 = recv_3_data_156; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_157 = recv_3_data_157; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_158 = recv_3_data_158; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_159 = recv_3_data_159; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_160 = recv_3_data_160; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_161 = recv_3_data_161; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_162 = recv_3_data_162; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_163 = recv_3_data_163; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_164 = recv_3_data_164; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_165 = recv_3_data_165; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_166 = recv_3_data_166; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_167 = recv_3_data_167; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_168 = recv_3_data_168; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_169 = recv_3_data_169; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_170 = recv_3_data_170; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_171 = recv_3_data_171; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_172 = recv_3_data_172; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_173 = recv_3_data_173; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_174 = recv_3_data_174; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_175 = recv_3_data_175; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_176 = recv_3_data_176; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_177 = recv_3_data_177; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_178 = recv_3_data_178; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_179 = recv_3_data_179; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_180 = recv_3_data_180; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_181 = recv_3_data_181; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_182 = recv_3_data_182; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_183 = recv_3_data_183; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_184 = recv_3_data_184; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_185 = recv_3_data_185; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_186 = recv_3_data_186; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_187 = recv_3_data_187; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_188 = recv_3_data_188; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_189 = recv_3_data_189; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_190 = recv_3_data_190; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_191 = recv_3_data_191; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_192 = recv_3_data_192; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_193 = recv_3_data_193; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_194 = recv_3_data_194; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_195 = recv_3_data_195; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_196 = recv_3_data_196; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_197 = recv_3_data_197; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_198 = recv_3_data_198; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_199 = recv_3_data_199; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_200 = recv_3_data_200; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_201 = recv_3_data_201; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_202 = recv_3_data_202; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_203 = recv_3_data_203; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_204 = recv_3_data_204; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_205 = recv_3_data_205; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_206 = recv_3_data_206; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_207 = recv_3_data_207; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_208 = recv_3_data_208; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_209 = recv_3_data_209; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_210 = recv_3_data_210; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_211 = recv_3_data_211; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_212 = recv_3_data_212; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_213 = recv_3_data_213; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_214 = recv_3_data_214; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_215 = recv_3_data_215; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_216 = recv_3_data_216; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_217 = recv_3_data_217; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_218 = recv_3_data_218; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_219 = recv_3_data_219; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_220 = recv_3_data_220; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_221 = recv_3_data_221; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_222 = recv_3_data_222; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_223 = recv_3_data_223; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_224 = recv_3_data_224; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_225 = recv_3_data_225; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_226 = recv_3_data_226; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_227 = recv_3_data_227; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_228 = recv_3_data_228; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_229 = recv_3_data_229; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_230 = recv_3_data_230; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_231 = recv_3_data_231; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_232 = recv_3_data_232; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_233 = recv_3_data_233; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_234 = recv_3_data_234; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_235 = recv_3_data_235; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_236 = recv_3_data_236; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_237 = recv_3_data_237; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_238 = recv_3_data_238; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_239 = recv_3_data_239; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_240 = recv_3_data_240; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_241 = recv_3_data_241; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_242 = recv_3_data_242; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_243 = recv_3_data_243; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_244 = recv_3_data_244; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_245 = recv_3_data_245; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_246 = recv_3_data_246; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_247 = recv_3_data_247; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_248 = recv_3_data_248; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_249 = recv_3_data_249; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_250 = recv_3_data_250; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_251 = recv_3_data_251; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_252 = recv_3_data_252; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_253 = recv_3_data_253; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_254 = recv_3_data_254; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_data_255 = recv_3_data_255; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_header_0 = recv_3_header_0; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_header_1 = recv_3_header_1; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_header_2 = recv_3_header_2; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_header_3 = recv_3_header_3; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_header_4 = recv_3_header_4; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_header_5 = recv_3_header_5; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_header_6 = recv_3_header_6; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_header_7 = recv_3_header_7; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_header_8 = recv_3_header_8; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_header_9 = recv_3_header_9; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_header_10 = recv_3_header_10; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_header_11 = recv_3_header_11; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_header_12 = recv_3_header_12; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_header_13 = recv_3_header_13; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_header_14 = recv_3_header_14; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_header_15 = recv_3_header_15; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_parse_current_state = recv_3_parse_current_state; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_parse_current_offset = recv_3_parse_current_offset; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_parse_transition_field = recv_3_parse_transition_field; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_next_processor_id = recv_3_next_processor_id; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_next_config_id = recv_3_next_config_id; // @[ipsa.scala 161:32]
  assign proc_3_io_pipe_phv_in_is_valid_processor = recv_3_is_valid_processor; // @[ipsa.scala 161:32]
  assign proc_3_io_mod_par_mod_en = io_mod_proc_mod_3_par_mod_en; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_par_mod_last_mau_id_mod = io_mod_proc_mod_3_par_mod_last_mau_id_mod; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_par_mod_last_mau_id = io_mod_proc_mod_3_par_mod_last_mau_id; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_par_mod_cs = io_mod_proc_mod_3_par_mod_cs; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_par_mod_module_mod_state_id_mod = io_mod_proc_mod_3_par_mod_module_mod_state_id_mod; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_par_mod_module_mod_state_id = io_mod_proc_mod_3_par_mod_module_mod_state_id; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_par_mod_module_mod_sram_w_cs = io_mod_proc_mod_3_par_mod_module_mod_sram_w_cs; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_par_mod_module_mod_sram_w_en = io_mod_proc_mod_3_par_mod_module_mod_sram_w_en; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_par_mod_module_mod_sram_w_addr = io_mod_proc_mod_3_par_mod_module_mod_sram_w_addr; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_par_mod_module_mod_sram_w_data = io_mod_proc_mod_3_par_mod_module_mod_sram_w_data; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_en = io_mod_proc_mod_3_mat_mod_en; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_config_id = io_mod_proc_mod_3_mat_mod_config_id; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_key_mod_header_id = io_mod_proc_mod_3_mat_mod_key_mod_header_id; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_key_mod_internal_offset = io_mod_proc_mod_3_mat_mod_key_mod_internal_offset; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_key_mod_key_length = io_mod_proc_mod_3_mat_mod_key_mod_key_length; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_0 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_0; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_1 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_1; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_2 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_2; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_3 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_3; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_4 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_4; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_5 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_5; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_6 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_6; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_7 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_7; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_8 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_8; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_9 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_9; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_10 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_10; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_11 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_11; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_12 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_12; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_13 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_13; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_14 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_14; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_15 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_15; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_16 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_16; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_17 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_17; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_18 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_18; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_19 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_19; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_20 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_20; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_21 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_21; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_22 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_22; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_23 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_23; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_24 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_24; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_25 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_25; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_26 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_26; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_27 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_27; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_28 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_28; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_29 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_29; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_30 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_30; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_31 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_31; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_32 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_32; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_33 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_33; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_34 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_34; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_35 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_35; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_36 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_36; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_37 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_37; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_38 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_38; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_39 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_39; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_40 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_40; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_41 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_41; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_42 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_42; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_43 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_43; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_44 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_44; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_45 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_45; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_46 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_46; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_47 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_47; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_48 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_48; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_49 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_49; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_50 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_50; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_51 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_51; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_52 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_52; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_53 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_53; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_54 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_54; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_55 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_55; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_56 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_56; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_57 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_57; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_58 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_58; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_59 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_59; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_60 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_60; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_61 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_61; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_62 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_62; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_sram_id_table_63 = io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_63; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_3_mat_mod_table_mod_table_width; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_3_mat_mod_table_mod_table_depth; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_act_mod_en_0 = io_mod_proc_mod_3_act_mod_en_0; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_act_mod_en_1 = io_mod_proc_mod_3_act_mod_en_1; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_act_mod_addr = io_mod_proc_mod_3_act_mod_addr; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_act_mod_data_0 = io_mod_proc_mod_3_act_mod_data_0; // @[ipsa.scala 63:20]
  assign proc_3_io_mod_act_mod_data_1 = io_mod_proc_mod_3_act_mod_data_1; // @[ipsa.scala 63:20]
  assign proc_3_io_mem_cluster_0_data = sram_cluster_0_io_r_3_cluster_0_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_1_data = sram_cluster_0_io_r_3_cluster_1_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_2_data = sram_cluster_0_io_r_3_cluster_2_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_3_data = sram_cluster_0_io_r_3_cluster_3_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_4_data = sram_cluster_0_io_r_3_cluster_4_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_5_data = sram_cluster_0_io_r_3_cluster_5_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_6_data = sram_cluster_0_io_r_3_cluster_6_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_7_data = sram_cluster_0_io_r_3_cluster_7_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_8_data = sram_cluster_0_io_r_3_cluster_8_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_9_data = sram_cluster_0_io_r_3_cluster_9_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_10_data = sram_cluster_0_io_r_3_cluster_10_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_11_data = sram_cluster_0_io_r_3_cluster_11_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_12_data = sram_cluster_0_io_r_3_cluster_12_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_13_data = sram_cluster_0_io_r_3_cluster_13_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_14_data = sram_cluster_0_io_r_3_cluster_14_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_15_data = sram_cluster_0_io_r_3_cluster_15_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_16_data = sram_cluster_0_io_r_3_cluster_16_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_17_data = sram_cluster_0_io_r_3_cluster_17_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_18_data = sram_cluster_0_io_r_3_cluster_18_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_19_data = sram_cluster_0_io_r_3_cluster_19_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_20_data = sram_cluster_0_io_r_3_cluster_20_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_21_data = sram_cluster_0_io_r_3_cluster_21_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_22_data = sram_cluster_0_io_r_3_cluster_22_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_23_data = sram_cluster_0_io_r_3_cluster_23_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_24_data = sram_cluster_0_io_r_3_cluster_24_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_25_data = sram_cluster_0_io_r_3_cluster_25_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_26_data = sram_cluster_0_io_r_3_cluster_26_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_27_data = sram_cluster_0_io_r_3_cluster_27_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_28_data = sram_cluster_0_io_r_3_cluster_28_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_29_data = sram_cluster_0_io_r_3_cluster_29_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_30_data = sram_cluster_0_io_r_3_cluster_30_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_31_data = sram_cluster_0_io_r_3_cluster_31_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_32_data = sram_cluster_0_io_r_3_cluster_32_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_33_data = sram_cluster_0_io_r_3_cluster_33_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_34_data = sram_cluster_0_io_r_3_cluster_34_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_35_data = sram_cluster_0_io_r_3_cluster_35_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_36_data = sram_cluster_0_io_r_3_cluster_36_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_37_data = sram_cluster_0_io_r_3_cluster_37_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_38_data = sram_cluster_0_io_r_3_cluster_38_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_39_data = sram_cluster_0_io_r_3_cluster_39_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_40_data = sram_cluster_0_io_r_3_cluster_40_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_41_data = sram_cluster_0_io_r_3_cluster_41_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_42_data = sram_cluster_0_io_r_3_cluster_42_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_43_data = sram_cluster_0_io_r_3_cluster_43_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_44_data = sram_cluster_0_io_r_3_cluster_44_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_45_data = sram_cluster_0_io_r_3_cluster_45_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_46_data = sram_cluster_0_io_r_3_cluster_46_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_47_data = sram_cluster_0_io_r_3_cluster_47_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_48_data = sram_cluster_0_io_r_3_cluster_48_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_49_data = sram_cluster_0_io_r_3_cluster_49_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_50_data = sram_cluster_0_io_r_3_cluster_50_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_51_data = sram_cluster_0_io_r_3_cluster_51_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_52_data = sram_cluster_0_io_r_3_cluster_52_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_53_data = sram_cluster_0_io_r_3_cluster_53_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_54_data = sram_cluster_0_io_r_3_cluster_54_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_55_data = sram_cluster_0_io_r_3_cluster_55_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_56_data = sram_cluster_0_io_r_3_cluster_56_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_57_data = sram_cluster_0_io_r_3_cluster_57_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_58_data = sram_cluster_0_io_r_3_cluster_58_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_59_data = sram_cluster_0_io_r_3_cluster_59_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_60_data = sram_cluster_0_io_r_3_cluster_60_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_61_data = sram_cluster_0_io_r_3_cluster_61_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_62_data = sram_cluster_0_io_r_3_cluster_62_data; // @[ipsa.scala 76:37]
  assign proc_3_io_mem_cluster_63_data = sram_cluster_0_io_r_3_cluster_63_data; // @[ipsa.scala 76:37]
  assign sram_cluster_0_clock = clock;
  assign sram_cluster_0_io_w_wcs = io_w_0_wcs; // @[ipsa.scala 69:18]
  assign sram_cluster_0_io_w_w_en = io_w_0_w_en; // @[ipsa.scala 69:18]
  assign sram_cluster_0_io_w_w_addr = io_w_0_w_addr; // @[ipsa.scala 69:18]
  assign sram_cluster_0_io_w_w_data = io_w_0_w_data; // @[ipsa.scala 69:18]
  assign sram_cluster_0_io_r_0_cluster_0_en = proc_0_io_mem_cluster_0_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_0_addr = proc_0_io_mem_cluster_0_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_1_en = proc_0_io_mem_cluster_1_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_1_addr = proc_0_io_mem_cluster_1_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_2_en = proc_0_io_mem_cluster_2_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_2_addr = proc_0_io_mem_cluster_2_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_3_en = proc_0_io_mem_cluster_3_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_3_addr = proc_0_io_mem_cluster_3_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_4_en = proc_0_io_mem_cluster_4_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_4_addr = proc_0_io_mem_cluster_4_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_5_en = proc_0_io_mem_cluster_5_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_5_addr = proc_0_io_mem_cluster_5_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_6_en = proc_0_io_mem_cluster_6_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_6_addr = proc_0_io_mem_cluster_6_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_7_en = proc_0_io_mem_cluster_7_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_7_addr = proc_0_io_mem_cluster_7_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_8_en = proc_0_io_mem_cluster_8_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_8_addr = proc_0_io_mem_cluster_8_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_9_en = proc_0_io_mem_cluster_9_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_9_addr = proc_0_io_mem_cluster_9_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_10_en = proc_0_io_mem_cluster_10_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_10_addr = proc_0_io_mem_cluster_10_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_11_en = proc_0_io_mem_cluster_11_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_11_addr = proc_0_io_mem_cluster_11_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_12_en = proc_0_io_mem_cluster_12_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_12_addr = proc_0_io_mem_cluster_12_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_13_en = proc_0_io_mem_cluster_13_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_13_addr = proc_0_io_mem_cluster_13_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_14_en = proc_0_io_mem_cluster_14_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_14_addr = proc_0_io_mem_cluster_14_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_15_en = proc_0_io_mem_cluster_15_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_15_addr = proc_0_io_mem_cluster_15_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_16_en = proc_0_io_mem_cluster_16_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_16_addr = proc_0_io_mem_cluster_16_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_17_en = proc_0_io_mem_cluster_17_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_17_addr = proc_0_io_mem_cluster_17_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_18_en = proc_0_io_mem_cluster_18_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_18_addr = proc_0_io_mem_cluster_18_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_19_en = proc_0_io_mem_cluster_19_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_19_addr = proc_0_io_mem_cluster_19_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_20_en = proc_0_io_mem_cluster_20_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_20_addr = proc_0_io_mem_cluster_20_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_21_en = proc_0_io_mem_cluster_21_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_21_addr = proc_0_io_mem_cluster_21_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_22_en = proc_0_io_mem_cluster_22_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_22_addr = proc_0_io_mem_cluster_22_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_23_en = proc_0_io_mem_cluster_23_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_23_addr = proc_0_io_mem_cluster_23_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_24_en = proc_0_io_mem_cluster_24_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_24_addr = proc_0_io_mem_cluster_24_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_25_en = proc_0_io_mem_cluster_25_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_25_addr = proc_0_io_mem_cluster_25_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_26_en = proc_0_io_mem_cluster_26_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_26_addr = proc_0_io_mem_cluster_26_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_27_en = proc_0_io_mem_cluster_27_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_27_addr = proc_0_io_mem_cluster_27_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_28_en = proc_0_io_mem_cluster_28_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_28_addr = proc_0_io_mem_cluster_28_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_29_en = proc_0_io_mem_cluster_29_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_29_addr = proc_0_io_mem_cluster_29_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_30_en = proc_0_io_mem_cluster_30_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_30_addr = proc_0_io_mem_cluster_30_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_31_en = proc_0_io_mem_cluster_31_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_31_addr = proc_0_io_mem_cluster_31_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_32_en = proc_0_io_mem_cluster_32_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_32_addr = proc_0_io_mem_cluster_32_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_33_en = proc_0_io_mem_cluster_33_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_33_addr = proc_0_io_mem_cluster_33_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_34_en = proc_0_io_mem_cluster_34_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_34_addr = proc_0_io_mem_cluster_34_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_35_en = proc_0_io_mem_cluster_35_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_35_addr = proc_0_io_mem_cluster_35_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_36_en = proc_0_io_mem_cluster_36_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_36_addr = proc_0_io_mem_cluster_36_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_37_en = proc_0_io_mem_cluster_37_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_37_addr = proc_0_io_mem_cluster_37_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_38_en = proc_0_io_mem_cluster_38_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_38_addr = proc_0_io_mem_cluster_38_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_39_en = proc_0_io_mem_cluster_39_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_39_addr = proc_0_io_mem_cluster_39_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_40_en = proc_0_io_mem_cluster_40_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_40_addr = proc_0_io_mem_cluster_40_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_41_en = proc_0_io_mem_cluster_41_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_41_addr = proc_0_io_mem_cluster_41_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_42_en = proc_0_io_mem_cluster_42_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_42_addr = proc_0_io_mem_cluster_42_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_43_en = proc_0_io_mem_cluster_43_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_43_addr = proc_0_io_mem_cluster_43_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_44_en = proc_0_io_mem_cluster_44_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_44_addr = proc_0_io_mem_cluster_44_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_45_en = proc_0_io_mem_cluster_45_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_45_addr = proc_0_io_mem_cluster_45_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_46_en = proc_0_io_mem_cluster_46_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_46_addr = proc_0_io_mem_cluster_46_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_47_en = proc_0_io_mem_cluster_47_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_47_addr = proc_0_io_mem_cluster_47_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_48_en = proc_0_io_mem_cluster_48_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_48_addr = proc_0_io_mem_cluster_48_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_49_en = proc_0_io_mem_cluster_49_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_49_addr = proc_0_io_mem_cluster_49_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_50_en = proc_0_io_mem_cluster_50_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_50_addr = proc_0_io_mem_cluster_50_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_51_en = proc_0_io_mem_cluster_51_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_51_addr = proc_0_io_mem_cluster_51_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_52_en = proc_0_io_mem_cluster_52_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_52_addr = proc_0_io_mem_cluster_52_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_53_en = proc_0_io_mem_cluster_53_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_53_addr = proc_0_io_mem_cluster_53_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_54_en = proc_0_io_mem_cluster_54_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_54_addr = proc_0_io_mem_cluster_54_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_55_en = proc_0_io_mem_cluster_55_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_55_addr = proc_0_io_mem_cluster_55_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_56_en = proc_0_io_mem_cluster_56_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_56_addr = proc_0_io_mem_cluster_56_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_57_en = proc_0_io_mem_cluster_57_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_57_addr = proc_0_io_mem_cluster_57_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_58_en = proc_0_io_mem_cluster_58_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_58_addr = proc_0_io_mem_cluster_58_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_59_en = proc_0_io_mem_cluster_59_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_59_addr = proc_0_io_mem_cluster_59_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_60_en = proc_0_io_mem_cluster_60_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_60_addr = proc_0_io_mem_cluster_60_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_61_en = proc_0_io_mem_cluster_61_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_61_addr = proc_0_io_mem_cluster_61_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_62_en = proc_0_io_mem_cluster_62_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_62_addr = proc_0_io_mem_cluster_62_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_63_en = proc_0_io_mem_cluster_63_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_0_cluster_63_addr = proc_0_io_mem_cluster_63_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_0_en = proc_1_io_mem_cluster_0_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_0_addr = proc_1_io_mem_cluster_0_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_1_en = proc_1_io_mem_cluster_1_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_1_addr = proc_1_io_mem_cluster_1_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_2_en = proc_1_io_mem_cluster_2_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_2_addr = proc_1_io_mem_cluster_2_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_3_en = proc_1_io_mem_cluster_3_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_3_addr = proc_1_io_mem_cluster_3_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_4_en = proc_1_io_mem_cluster_4_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_4_addr = proc_1_io_mem_cluster_4_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_5_en = proc_1_io_mem_cluster_5_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_5_addr = proc_1_io_mem_cluster_5_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_6_en = proc_1_io_mem_cluster_6_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_6_addr = proc_1_io_mem_cluster_6_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_7_en = proc_1_io_mem_cluster_7_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_7_addr = proc_1_io_mem_cluster_7_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_8_en = proc_1_io_mem_cluster_8_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_8_addr = proc_1_io_mem_cluster_8_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_9_en = proc_1_io_mem_cluster_9_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_9_addr = proc_1_io_mem_cluster_9_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_10_en = proc_1_io_mem_cluster_10_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_10_addr = proc_1_io_mem_cluster_10_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_11_en = proc_1_io_mem_cluster_11_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_11_addr = proc_1_io_mem_cluster_11_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_12_en = proc_1_io_mem_cluster_12_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_12_addr = proc_1_io_mem_cluster_12_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_13_en = proc_1_io_mem_cluster_13_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_13_addr = proc_1_io_mem_cluster_13_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_14_en = proc_1_io_mem_cluster_14_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_14_addr = proc_1_io_mem_cluster_14_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_15_en = proc_1_io_mem_cluster_15_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_15_addr = proc_1_io_mem_cluster_15_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_16_en = proc_1_io_mem_cluster_16_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_16_addr = proc_1_io_mem_cluster_16_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_17_en = proc_1_io_mem_cluster_17_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_17_addr = proc_1_io_mem_cluster_17_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_18_en = proc_1_io_mem_cluster_18_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_18_addr = proc_1_io_mem_cluster_18_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_19_en = proc_1_io_mem_cluster_19_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_19_addr = proc_1_io_mem_cluster_19_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_20_en = proc_1_io_mem_cluster_20_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_20_addr = proc_1_io_mem_cluster_20_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_21_en = proc_1_io_mem_cluster_21_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_21_addr = proc_1_io_mem_cluster_21_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_22_en = proc_1_io_mem_cluster_22_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_22_addr = proc_1_io_mem_cluster_22_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_23_en = proc_1_io_mem_cluster_23_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_23_addr = proc_1_io_mem_cluster_23_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_24_en = proc_1_io_mem_cluster_24_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_24_addr = proc_1_io_mem_cluster_24_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_25_en = proc_1_io_mem_cluster_25_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_25_addr = proc_1_io_mem_cluster_25_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_26_en = proc_1_io_mem_cluster_26_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_26_addr = proc_1_io_mem_cluster_26_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_27_en = proc_1_io_mem_cluster_27_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_27_addr = proc_1_io_mem_cluster_27_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_28_en = proc_1_io_mem_cluster_28_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_28_addr = proc_1_io_mem_cluster_28_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_29_en = proc_1_io_mem_cluster_29_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_29_addr = proc_1_io_mem_cluster_29_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_30_en = proc_1_io_mem_cluster_30_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_30_addr = proc_1_io_mem_cluster_30_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_31_en = proc_1_io_mem_cluster_31_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_31_addr = proc_1_io_mem_cluster_31_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_32_en = proc_1_io_mem_cluster_32_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_32_addr = proc_1_io_mem_cluster_32_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_33_en = proc_1_io_mem_cluster_33_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_33_addr = proc_1_io_mem_cluster_33_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_34_en = proc_1_io_mem_cluster_34_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_34_addr = proc_1_io_mem_cluster_34_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_35_en = proc_1_io_mem_cluster_35_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_35_addr = proc_1_io_mem_cluster_35_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_36_en = proc_1_io_mem_cluster_36_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_36_addr = proc_1_io_mem_cluster_36_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_37_en = proc_1_io_mem_cluster_37_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_37_addr = proc_1_io_mem_cluster_37_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_38_en = proc_1_io_mem_cluster_38_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_38_addr = proc_1_io_mem_cluster_38_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_39_en = proc_1_io_mem_cluster_39_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_39_addr = proc_1_io_mem_cluster_39_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_40_en = proc_1_io_mem_cluster_40_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_40_addr = proc_1_io_mem_cluster_40_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_41_en = proc_1_io_mem_cluster_41_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_41_addr = proc_1_io_mem_cluster_41_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_42_en = proc_1_io_mem_cluster_42_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_42_addr = proc_1_io_mem_cluster_42_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_43_en = proc_1_io_mem_cluster_43_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_43_addr = proc_1_io_mem_cluster_43_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_44_en = proc_1_io_mem_cluster_44_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_44_addr = proc_1_io_mem_cluster_44_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_45_en = proc_1_io_mem_cluster_45_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_45_addr = proc_1_io_mem_cluster_45_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_46_en = proc_1_io_mem_cluster_46_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_46_addr = proc_1_io_mem_cluster_46_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_47_en = proc_1_io_mem_cluster_47_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_47_addr = proc_1_io_mem_cluster_47_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_48_en = proc_1_io_mem_cluster_48_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_48_addr = proc_1_io_mem_cluster_48_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_49_en = proc_1_io_mem_cluster_49_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_49_addr = proc_1_io_mem_cluster_49_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_50_en = proc_1_io_mem_cluster_50_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_50_addr = proc_1_io_mem_cluster_50_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_51_en = proc_1_io_mem_cluster_51_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_51_addr = proc_1_io_mem_cluster_51_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_52_en = proc_1_io_mem_cluster_52_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_52_addr = proc_1_io_mem_cluster_52_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_53_en = proc_1_io_mem_cluster_53_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_53_addr = proc_1_io_mem_cluster_53_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_54_en = proc_1_io_mem_cluster_54_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_54_addr = proc_1_io_mem_cluster_54_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_55_en = proc_1_io_mem_cluster_55_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_55_addr = proc_1_io_mem_cluster_55_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_56_en = proc_1_io_mem_cluster_56_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_56_addr = proc_1_io_mem_cluster_56_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_57_en = proc_1_io_mem_cluster_57_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_57_addr = proc_1_io_mem_cluster_57_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_58_en = proc_1_io_mem_cluster_58_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_58_addr = proc_1_io_mem_cluster_58_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_59_en = proc_1_io_mem_cluster_59_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_59_addr = proc_1_io_mem_cluster_59_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_60_en = proc_1_io_mem_cluster_60_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_60_addr = proc_1_io_mem_cluster_60_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_61_en = proc_1_io_mem_cluster_61_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_61_addr = proc_1_io_mem_cluster_61_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_62_en = proc_1_io_mem_cluster_62_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_62_addr = proc_1_io_mem_cluster_62_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_63_en = proc_1_io_mem_cluster_63_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_1_cluster_63_addr = proc_1_io_mem_cluster_63_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_0_en = proc_2_io_mem_cluster_0_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_0_addr = proc_2_io_mem_cluster_0_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_1_en = proc_2_io_mem_cluster_1_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_1_addr = proc_2_io_mem_cluster_1_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_2_en = proc_2_io_mem_cluster_2_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_2_addr = proc_2_io_mem_cluster_2_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_3_en = proc_2_io_mem_cluster_3_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_3_addr = proc_2_io_mem_cluster_3_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_4_en = proc_2_io_mem_cluster_4_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_4_addr = proc_2_io_mem_cluster_4_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_5_en = proc_2_io_mem_cluster_5_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_5_addr = proc_2_io_mem_cluster_5_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_6_en = proc_2_io_mem_cluster_6_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_6_addr = proc_2_io_mem_cluster_6_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_7_en = proc_2_io_mem_cluster_7_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_7_addr = proc_2_io_mem_cluster_7_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_8_en = proc_2_io_mem_cluster_8_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_8_addr = proc_2_io_mem_cluster_8_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_9_en = proc_2_io_mem_cluster_9_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_9_addr = proc_2_io_mem_cluster_9_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_10_en = proc_2_io_mem_cluster_10_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_10_addr = proc_2_io_mem_cluster_10_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_11_en = proc_2_io_mem_cluster_11_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_11_addr = proc_2_io_mem_cluster_11_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_12_en = proc_2_io_mem_cluster_12_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_12_addr = proc_2_io_mem_cluster_12_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_13_en = proc_2_io_mem_cluster_13_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_13_addr = proc_2_io_mem_cluster_13_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_14_en = proc_2_io_mem_cluster_14_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_14_addr = proc_2_io_mem_cluster_14_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_15_en = proc_2_io_mem_cluster_15_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_15_addr = proc_2_io_mem_cluster_15_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_16_en = proc_2_io_mem_cluster_16_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_16_addr = proc_2_io_mem_cluster_16_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_17_en = proc_2_io_mem_cluster_17_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_17_addr = proc_2_io_mem_cluster_17_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_18_en = proc_2_io_mem_cluster_18_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_18_addr = proc_2_io_mem_cluster_18_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_19_en = proc_2_io_mem_cluster_19_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_19_addr = proc_2_io_mem_cluster_19_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_20_en = proc_2_io_mem_cluster_20_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_20_addr = proc_2_io_mem_cluster_20_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_21_en = proc_2_io_mem_cluster_21_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_21_addr = proc_2_io_mem_cluster_21_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_22_en = proc_2_io_mem_cluster_22_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_22_addr = proc_2_io_mem_cluster_22_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_23_en = proc_2_io_mem_cluster_23_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_23_addr = proc_2_io_mem_cluster_23_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_24_en = proc_2_io_mem_cluster_24_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_24_addr = proc_2_io_mem_cluster_24_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_25_en = proc_2_io_mem_cluster_25_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_25_addr = proc_2_io_mem_cluster_25_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_26_en = proc_2_io_mem_cluster_26_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_26_addr = proc_2_io_mem_cluster_26_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_27_en = proc_2_io_mem_cluster_27_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_27_addr = proc_2_io_mem_cluster_27_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_28_en = proc_2_io_mem_cluster_28_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_28_addr = proc_2_io_mem_cluster_28_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_29_en = proc_2_io_mem_cluster_29_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_29_addr = proc_2_io_mem_cluster_29_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_30_en = proc_2_io_mem_cluster_30_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_30_addr = proc_2_io_mem_cluster_30_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_31_en = proc_2_io_mem_cluster_31_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_31_addr = proc_2_io_mem_cluster_31_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_32_en = proc_2_io_mem_cluster_32_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_32_addr = proc_2_io_mem_cluster_32_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_33_en = proc_2_io_mem_cluster_33_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_33_addr = proc_2_io_mem_cluster_33_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_34_en = proc_2_io_mem_cluster_34_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_34_addr = proc_2_io_mem_cluster_34_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_35_en = proc_2_io_mem_cluster_35_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_35_addr = proc_2_io_mem_cluster_35_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_36_en = proc_2_io_mem_cluster_36_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_36_addr = proc_2_io_mem_cluster_36_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_37_en = proc_2_io_mem_cluster_37_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_37_addr = proc_2_io_mem_cluster_37_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_38_en = proc_2_io_mem_cluster_38_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_38_addr = proc_2_io_mem_cluster_38_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_39_en = proc_2_io_mem_cluster_39_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_39_addr = proc_2_io_mem_cluster_39_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_40_en = proc_2_io_mem_cluster_40_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_40_addr = proc_2_io_mem_cluster_40_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_41_en = proc_2_io_mem_cluster_41_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_41_addr = proc_2_io_mem_cluster_41_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_42_en = proc_2_io_mem_cluster_42_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_42_addr = proc_2_io_mem_cluster_42_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_43_en = proc_2_io_mem_cluster_43_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_43_addr = proc_2_io_mem_cluster_43_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_44_en = proc_2_io_mem_cluster_44_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_44_addr = proc_2_io_mem_cluster_44_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_45_en = proc_2_io_mem_cluster_45_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_45_addr = proc_2_io_mem_cluster_45_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_46_en = proc_2_io_mem_cluster_46_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_46_addr = proc_2_io_mem_cluster_46_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_47_en = proc_2_io_mem_cluster_47_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_47_addr = proc_2_io_mem_cluster_47_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_48_en = proc_2_io_mem_cluster_48_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_48_addr = proc_2_io_mem_cluster_48_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_49_en = proc_2_io_mem_cluster_49_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_49_addr = proc_2_io_mem_cluster_49_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_50_en = proc_2_io_mem_cluster_50_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_50_addr = proc_2_io_mem_cluster_50_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_51_en = proc_2_io_mem_cluster_51_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_51_addr = proc_2_io_mem_cluster_51_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_52_en = proc_2_io_mem_cluster_52_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_52_addr = proc_2_io_mem_cluster_52_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_53_en = proc_2_io_mem_cluster_53_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_53_addr = proc_2_io_mem_cluster_53_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_54_en = proc_2_io_mem_cluster_54_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_54_addr = proc_2_io_mem_cluster_54_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_55_en = proc_2_io_mem_cluster_55_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_55_addr = proc_2_io_mem_cluster_55_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_56_en = proc_2_io_mem_cluster_56_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_56_addr = proc_2_io_mem_cluster_56_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_57_en = proc_2_io_mem_cluster_57_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_57_addr = proc_2_io_mem_cluster_57_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_58_en = proc_2_io_mem_cluster_58_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_58_addr = proc_2_io_mem_cluster_58_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_59_en = proc_2_io_mem_cluster_59_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_59_addr = proc_2_io_mem_cluster_59_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_60_en = proc_2_io_mem_cluster_60_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_60_addr = proc_2_io_mem_cluster_60_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_61_en = proc_2_io_mem_cluster_61_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_61_addr = proc_2_io_mem_cluster_61_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_62_en = proc_2_io_mem_cluster_62_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_62_addr = proc_2_io_mem_cluster_62_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_63_en = proc_2_io_mem_cluster_63_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_2_cluster_63_addr = proc_2_io_mem_cluster_63_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_0_en = proc_3_io_mem_cluster_0_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_0_addr = proc_3_io_mem_cluster_0_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_1_en = proc_3_io_mem_cluster_1_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_1_addr = proc_3_io_mem_cluster_1_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_2_en = proc_3_io_mem_cluster_2_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_2_addr = proc_3_io_mem_cluster_2_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_3_en = proc_3_io_mem_cluster_3_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_3_addr = proc_3_io_mem_cluster_3_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_4_en = proc_3_io_mem_cluster_4_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_4_addr = proc_3_io_mem_cluster_4_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_5_en = proc_3_io_mem_cluster_5_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_5_addr = proc_3_io_mem_cluster_5_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_6_en = proc_3_io_mem_cluster_6_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_6_addr = proc_3_io_mem_cluster_6_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_7_en = proc_3_io_mem_cluster_7_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_7_addr = proc_3_io_mem_cluster_7_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_8_en = proc_3_io_mem_cluster_8_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_8_addr = proc_3_io_mem_cluster_8_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_9_en = proc_3_io_mem_cluster_9_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_9_addr = proc_3_io_mem_cluster_9_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_10_en = proc_3_io_mem_cluster_10_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_10_addr = proc_3_io_mem_cluster_10_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_11_en = proc_3_io_mem_cluster_11_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_11_addr = proc_3_io_mem_cluster_11_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_12_en = proc_3_io_mem_cluster_12_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_12_addr = proc_3_io_mem_cluster_12_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_13_en = proc_3_io_mem_cluster_13_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_13_addr = proc_3_io_mem_cluster_13_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_14_en = proc_3_io_mem_cluster_14_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_14_addr = proc_3_io_mem_cluster_14_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_15_en = proc_3_io_mem_cluster_15_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_15_addr = proc_3_io_mem_cluster_15_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_16_en = proc_3_io_mem_cluster_16_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_16_addr = proc_3_io_mem_cluster_16_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_17_en = proc_3_io_mem_cluster_17_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_17_addr = proc_3_io_mem_cluster_17_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_18_en = proc_3_io_mem_cluster_18_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_18_addr = proc_3_io_mem_cluster_18_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_19_en = proc_3_io_mem_cluster_19_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_19_addr = proc_3_io_mem_cluster_19_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_20_en = proc_3_io_mem_cluster_20_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_20_addr = proc_3_io_mem_cluster_20_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_21_en = proc_3_io_mem_cluster_21_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_21_addr = proc_3_io_mem_cluster_21_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_22_en = proc_3_io_mem_cluster_22_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_22_addr = proc_3_io_mem_cluster_22_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_23_en = proc_3_io_mem_cluster_23_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_23_addr = proc_3_io_mem_cluster_23_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_24_en = proc_3_io_mem_cluster_24_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_24_addr = proc_3_io_mem_cluster_24_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_25_en = proc_3_io_mem_cluster_25_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_25_addr = proc_3_io_mem_cluster_25_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_26_en = proc_3_io_mem_cluster_26_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_26_addr = proc_3_io_mem_cluster_26_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_27_en = proc_3_io_mem_cluster_27_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_27_addr = proc_3_io_mem_cluster_27_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_28_en = proc_3_io_mem_cluster_28_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_28_addr = proc_3_io_mem_cluster_28_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_29_en = proc_3_io_mem_cluster_29_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_29_addr = proc_3_io_mem_cluster_29_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_30_en = proc_3_io_mem_cluster_30_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_30_addr = proc_3_io_mem_cluster_30_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_31_en = proc_3_io_mem_cluster_31_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_31_addr = proc_3_io_mem_cluster_31_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_32_en = proc_3_io_mem_cluster_32_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_32_addr = proc_3_io_mem_cluster_32_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_33_en = proc_3_io_mem_cluster_33_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_33_addr = proc_3_io_mem_cluster_33_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_34_en = proc_3_io_mem_cluster_34_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_34_addr = proc_3_io_mem_cluster_34_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_35_en = proc_3_io_mem_cluster_35_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_35_addr = proc_3_io_mem_cluster_35_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_36_en = proc_3_io_mem_cluster_36_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_36_addr = proc_3_io_mem_cluster_36_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_37_en = proc_3_io_mem_cluster_37_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_37_addr = proc_3_io_mem_cluster_37_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_38_en = proc_3_io_mem_cluster_38_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_38_addr = proc_3_io_mem_cluster_38_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_39_en = proc_3_io_mem_cluster_39_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_39_addr = proc_3_io_mem_cluster_39_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_40_en = proc_3_io_mem_cluster_40_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_40_addr = proc_3_io_mem_cluster_40_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_41_en = proc_3_io_mem_cluster_41_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_41_addr = proc_3_io_mem_cluster_41_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_42_en = proc_3_io_mem_cluster_42_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_42_addr = proc_3_io_mem_cluster_42_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_43_en = proc_3_io_mem_cluster_43_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_43_addr = proc_3_io_mem_cluster_43_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_44_en = proc_3_io_mem_cluster_44_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_44_addr = proc_3_io_mem_cluster_44_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_45_en = proc_3_io_mem_cluster_45_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_45_addr = proc_3_io_mem_cluster_45_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_46_en = proc_3_io_mem_cluster_46_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_46_addr = proc_3_io_mem_cluster_46_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_47_en = proc_3_io_mem_cluster_47_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_47_addr = proc_3_io_mem_cluster_47_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_48_en = proc_3_io_mem_cluster_48_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_48_addr = proc_3_io_mem_cluster_48_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_49_en = proc_3_io_mem_cluster_49_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_49_addr = proc_3_io_mem_cluster_49_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_50_en = proc_3_io_mem_cluster_50_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_50_addr = proc_3_io_mem_cluster_50_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_51_en = proc_3_io_mem_cluster_51_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_51_addr = proc_3_io_mem_cluster_51_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_52_en = proc_3_io_mem_cluster_52_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_52_addr = proc_3_io_mem_cluster_52_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_53_en = proc_3_io_mem_cluster_53_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_53_addr = proc_3_io_mem_cluster_53_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_54_en = proc_3_io_mem_cluster_54_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_54_addr = proc_3_io_mem_cluster_54_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_55_en = proc_3_io_mem_cluster_55_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_55_addr = proc_3_io_mem_cluster_55_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_56_en = proc_3_io_mem_cluster_56_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_56_addr = proc_3_io_mem_cluster_56_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_57_en = proc_3_io_mem_cluster_57_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_57_addr = proc_3_io_mem_cluster_57_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_58_en = proc_3_io_mem_cluster_58_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_58_addr = proc_3_io_mem_cluster_58_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_59_en = proc_3_io_mem_cluster_59_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_59_addr = proc_3_io_mem_cluster_59_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_60_en = proc_3_io_mem_cluster_60_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_60_addr = proc_3_io_mem_cluster_60_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_61_en = proc_3_io_mem_cluster_61_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_61_addr = proc_3_io_mem_cluster_61_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_62_en = proc_3_io_mem_cluster_62_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_62_addr = proc_3_io_mem_cluster_62_addr; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_63_en = proc_3_io_mem_cluster_63_en; // @[ipsa.scala 76:37]
  assign sram_cluster_0_io_r_3_cluster_63_addr = proc_3_io_mem_cluster_63_addr; // @[ipsa.scala 76:37]
  assign init_clock = clock;
  assign init_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_160 = io_pipe_phv_in_data_160; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_161 = io_pipe_phv_in_data_161; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_162 = io_pipe_phv_in_data_162; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_163 = io_pipe_phv_in_data_163; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_164 = io_pipe_phv_in_data_164; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_165 = io_pipe_phv_in_data_165; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_166 = io_pipe_phv_in_data_166; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_167 = io_pipe_phv_in_data_167; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_168 = io_pipe_phv_in_data_168; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_169 = io_pipe_phv_in_data_169; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_170 = io_pipe_phv_in_data_170; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_171 = io_pipe_phv_in_data_171; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_172 = io_pipe_phv_in_data_172; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_173 = io_pipe_phv_in_data_173; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_174 = io_pipe_phv_in_data_174; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_175 = io_pipe_phv_in_data_175; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_176 = io_pipe_phv_in_data_176; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_177 = io_pipe_phv_in_data_177; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_178 = io_pipe_phv_in_data_178; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_179 = io_pipe_phv_in_data_179; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_180 = io_pipe_phv_in_data_180; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_181 = io_pipe_phv_in_data_181; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_182 = io_pipe_phv_in_data_182; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_183 = io_pipe_phv_in_data_183; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_184 = io_pipe_phv_in_data_184; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_185 = io_pipe_phv_in_data_185; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_186 = io_pipe_phv_in_data_186; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_187 = io_pipe_phv_in_data_187; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_188 = io_pipe_phv_in_data_188; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_189 = io_pipe_phv_in_data_189; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_190 = io_pipe_phv_in_data_190; // @[ipsa.scala 81:25]
  assign init_io_pipe_phv_in_data_191 = io_pipe_phv_in_data_191; // @[ipsa.scala 81:25]
  assign init_io_first_proc_id = first_proc_id; // @[ipsa.scala 82:27]
  assign trans_0_clock = clock;
  assign trans_0_io_pipe_phv_in_data_0 = proc_0_io_pipe_phv_out_data_0; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_1 = proc_0_io_pipe_phv_out_data_1; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_2 = proc_0_io_pipe_phv_out_data_2; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_3 = proc_0_io_pipe_phv_out_data_3; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_4 = proc_0_io_pipe_phv_out_data_4; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_5 = proc_0_io_pipe_phv_out_data_5; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_6 = proc_0_io_pipe_phv_out_data_6; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_7 = proc_0_io_pipe_phv_out_data_7; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_8 = proc_0_io_pipe_phv_out_data_8; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_9 = proc_0_io_pipe_phv_out_data_9; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_10 = proc_0_io_pipe_phv_out_data_10; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_11 = proc_0_io_pipe_phv_out_data_11; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_12 = proc_0_io_pipe_phv_out_data_12; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_13 = proc_0_io_pipe_phv_out_data_13; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_14 = proc_0_io_pipe_phv_out_data_14; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_15 = proc_0_io_pipe_phv_out_data_15; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_16 = proc_0_io_pipe_phv_out_data_16; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_17 = proc_0_io_pipe_phv_out_data_17; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_18 = proc_0_io_pipe_phv_out_data_18; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_19 = proc_0_io_pipe_phv_out_data_19; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_20 = proc_0_io_pipe_phv_out_data_20; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_21 = proc_0_io_pipe_phv_out_data_21; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_22 = proc_0_io_pipe_phv_out_data_22; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_23 = proc_0_io_pipe_phv_out_data_23; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_24 = proc_0_io_pipe_phv_out_data_24; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_25 = proc_0_io_pipe_phv_out_data_25; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_26 = proc_0_io_pipe_phv_out_data_26; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_27 = proc_0_io_pipe_phv_out_data_27; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_28 = proc_0_io_pipe_phv_out_data_28; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_29 = proc_0_io_pipe_phv_out_data_29; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_30 = proc_0_io_pipe_phv_out_data_30; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_31 = proc_0_io_pipe_phv_out_data_31; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_32 = proc_0_io_pipe_phv_out_data_32; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_33 = proc_0_io_pipe_phv_out_data_33; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_34 = proc_0_io_pipe_phv_out_data_34; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_35 = proc_0_io_pipe_phv_out_data_35; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_36 = proc_0_io_pipe_phv_out_data_36; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_37 = proc_0_io_pipe_phv_out_data_37; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_38 = proc_0_io_pipe_phv_out_data_38; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_39 = proc_0_io_pipe_phv_out_data_39; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_40 = proc_0_io_pipe_phv_out_data_40; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_41 = proc_0_io_pipe_phv_out_data_41; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_42 = proc_0_io_pipe_phv_out_data_42; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_43 = proc_0_io_pipe_phv_out_data_43; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_44 = proc_0_io_pipe_phv_out_data_44; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_45 = proc_0_io_pipe_phv_out_data_45; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_46 = proc_0_io_pipe_phv_out_data_46; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_47 = proc_0_io_pipe_phv_out_data_47; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_48 = proc_0_io_pipe_phv_out_data_48; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_49 = proc_0_io_pipe_phv_out_data_49; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_50 = proc_0_io_pipe_phv_out_data_50; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_51 = proc_0_io_pipe_phv_out_data_51; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_52 = proc_0_io_pipe_phv_out_data_52; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_53 = proc_0_io_pipe_phv_out_data_53; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_54 = proc_0_io_pipe_phv_out_data_54; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_55 = proc_0_io_pipe_phv_out_data_55; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_56 = proc_0_io_pipe_phv_out_data_56; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_57 = proc_0_io_pipe_phv_out_data_57; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_58 = proc_0_io_pipe_phv_out_data_58; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_59 = proc_0_io_pipe_phv_out_data_59; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_60 = proc_0_io_pipe_phv_out_data_60; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_61 = proc_0_io_pipe_phv_out_data_61; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_62 = proc_0_io_pipe_phv_out_data_62; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_63 = proc_0_io_pipe_phv_out_data_63; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_64 = proc_0_io_pipe_phv_out_data_64; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_65 = proc_0_io_pipe_phv_out_data_65; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_66 = proc_0_io_pipe_phv_out_data_66; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_67 = proc_0_io_pipe_phv_out_data_67; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_68 = proc_0_io_pipe_phv_out_data_68; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_69 = proc_0_io_pipe_phv_out_data_69; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_70 = proc_0_io_pipe_phv_out_data_70; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_71 = proc_0_io_pipe_phv_out_data_71; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_72 = proc_0_io_pipe_phv_out_data_72; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_73 = proc_0_io_pipe_phv_out_data_73; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_74 = proc_0_io_pipe_phv_out_data_74; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_75 = proc_0_io_pipe_phv_out_data_75; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_76 = proc_0_io_pipe_phv_out_data_76; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_77 = proc_0_io_pipe_phv_out_data_77; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_78 = proc_0_io_pipe_phv_out_data_78; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_79 = proc_0_io_pipe_phv_out_data_79; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_80 = proc_0_io_pipe_phv_out_data_80; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_81 = proc_0_io_pipe_phv_out_data_81; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_82 = proc_0_io_pipe_phv_out_data_82; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_83 = proc_0_io_pipe_phv_out_data_83; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_84 = proc_0_io_pipe_phv_out_data_84; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_85 = proc_0_io_pipe_phv_out_data_85; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_86 = proc_0_io_pipe_phv_out_data_86; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_87 = proc_0_io_pipe_phv_out_data_87; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_88 = proc_0_io_pipe_phv_out_data_88; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_89 = proc_0_io_pipe_phv_out_data_89; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_90 = proc_0_io_pipe_phv_out_data_90; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_91 = proc_0_io_pipe_phv_out_data_91; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_92 = proc_0_io_pipe_phv_out_data_92; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_93 = proc_0_io_pipe_phv_out_data_93; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_94 = proc_0_io_pipe_phv_out_data_94; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_95 = proc_0_io_pipe_phv_out_data_95; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_96 = proc_0_io_pipe_phv_out_data_96; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_97 = proc_0_io_pipe_phv_out_data_97; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_98 = proc_0_io_pipe_phv_out_data_98; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_99 = proc_0_io_pipe_phv_out_data_99; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_100 = proc_0_io_pipe_phv_out_data_100; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_101 = proc_0_io_pipe_phv_out_data_101; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_102 = proc_0_io_pipe_phv_out_data_102; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_103 = proc_0_io_pipe_phv_out_data_103; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_104 = proc_0_io_pipe_phv_out_data_104; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_105 = proc_0_io_pipe_phv_out_data_105; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_106 = proc_0_io_pipe_phv_out_data_106; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_107 = proc_0_io_pipe_phv_out_data_107; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_108 = proc_0_io_pipe_phv_out_data_108; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_109 = proc_0_io_pipe_phv_out_data_109; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_110 = proc_0_io_pipe_phv_out_data_110; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_111 = proc_0_io_pipe_phv_out_data_111; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_112 = proc_0_io_pipe_phv_out_data_112; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_113 = proc_0_io_pipe_phv_out_data_113; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_114 = proc_0_io_pipe_phv_out_data_114; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_115 = proc_0_io_pipe_phv_out_data_115; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_116 = proc_0_io_pipe_phv_out_data_116; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_117 = proc_0_io_pipe_phv_out_data_117; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_118 = proc_0_io_pipe_phv_out_data_118; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_119 = proc_0_io_pipe_phv_out_data_119; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_120 = proc_0_io_pipe_phv_out_data_120; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_121 = proc_0_io_pipe_phv_out_data_121; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_122 = proc_0_io_pipe_phv_out_data_122; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_123 = proc_0_io_pipe_phv_out_data_123; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_124 = proc_0_io_pipe_phv_out_data_124; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_125 = proc_0_io_pipe_phv_out_data_125; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_126 = proc_0_io_pipe_phv_out_data_126; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_127 = proc_0_io_pipe_phv_out_data_127; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_128 = proc_0_io_pipe_phv_out_data_128; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_129 = proc_0_io_pipe_phv_out_data_129; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_130 = proc_0_io_pipe_phv_out_data_130; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_131 = proc_0_io_pipe_phv_out_data_131; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_132 = proc_0_io_pipe_phv_out_data_132; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_133 = proc_0_io_pipe_phv_out_data_133; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_134 = proc_0_io_pipe_phv_out_data_134; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_135 = proc_0_io_pipe_phv_out_data_135; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_136 = proc_0_io_pipe_phv_out_data_136; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_137 = proc_0_io_pipe_phv_out_data_137; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_138 = proc_0_io_pipe_phv_out_data_138; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_139 = proc_0_io_pipe_phv_out_data_139; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_140 = proc_0_io_pipe_phv_out_data_140; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_141 = proc_0_io_pipe_phv_out_data_141; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_142 = proc_0_io_pipe_phv_out_data_142; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_143 = proc_0_io_pipe_phv_out_data_143; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_144 = proc_0_io_pipe_phv_out_data_144; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_145 = proc_0_io_pipe_phv_out_data_145; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_146 = proc_0_io_pipe_phv_out_data_146; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_147 = proc_0_io_pipe_phv_out_data_147; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_148 = proc_0_io_pipe_phv_out_data_148; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_149 = proc_0_io_pipe_phv_out_data_149; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_150 = proc_0_io_pipe_phv_out_data_150; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_151 = proc_0_io_pipe_phv_out_data_151; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_152 = proc_0_io_pipe_phv_out_data_152; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_153 = proc_0_io_pipe_phv_out_data_153; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_154 = proc_0_io_pipe_phv_out_data_154; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_155 = proc_0_io_pipe_phv_out_data_155; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_156 = proc_0_io_pipe_phv_out_data_156; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_157 = proc_0_io_pipe_phv_out_data_157; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_158 = proc_0_io_pipe_phv_out_data_158; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_159 = proc_0_io_pipe_phv_out_data_159; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_160 = proc_0_io_pipe_phv_out_data_160; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_161 = proc_0_io_pipe_phv_out_data_161; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_162 = proc_0_io_pipe_phv_out_data_162; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_163 = proc_0_io_pipe_phv_out_data_163; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_164 = proc_0_io_pipe_phv_out_data_164; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_165 = proc_0_io_pipe_phv_out_data_165; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_166 = proc_0_io_pipe_phv_out_data_166; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_167 = proc_0_io_pipe_phv_out_data_167; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_168 = proc_0_io_pipe_phv_out_data_168; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_169 = proc_0_io_pipe_phv_out_data_169; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_170 = proc_0_io_pipe_phv_out_data_170; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_171 = proc_0_io_pipe_phv_out_data_171; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_172 = proc_0_io_pipe_phv_out_data_172; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_173 = proc_0_io_pipe_phv_out_data_173; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_174 = proc_0_io_pipe_phv_out_data_174; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_175 = proc_0_io_pipe_phv_out_data_175; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_176 = proc_0_io_pipe_phv_out_data_176; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_177 = proc_0_io_pipe_phv_out_data_177; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_178 = proc_0_io_pipe_phv_out_data_178; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_179 = proc_0_io_pipe_phv_out_data_179; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_180 = proc_0_io_pipe_phv_out_data_180; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_181 = proc_0_io_pipe_phv_out_data_181; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_182 = proc_0_io_pipe_phv_out_data_182; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_183 = proc_0_io_pipe_phv_out_data_183; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_184 = proc_0_io_pipe_phv_out_data_184; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_185 = proc_0_io_pipe_phv_out_data_185; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_186 = proc_0_io_pipe_phv_out_data_186; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_187 = proc_0_io_pipe_phv_out_data_187; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_188 = proc_0_io_pipe_phv_out_data_188; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_189 = proc_0_io_pipe_phv_out_data_189; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_190 = proc_0_io_pipe_phv_out_data_190; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_191 = proc_0_io_pipe_phv_out_data_191; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_192 = proc_0_io_pipe_phv_out_data_192; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_193 = proc_0_io_pipe_phv_out_data_193; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_194 = proc_0_io_pipe_phv_out_data_194; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_195 = proc_0_io_pipe_phv_out_data_195; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_196 = proc_0_io_pipe_phv_out_data_196; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_197 = proc_0_io_pipe_phv_out_data_197; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_198 = proc_0_io_pipe_phv_out_data_198; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_199 = proc_0_io_pipe_phv_out_data_199; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_200 = proc_0_io_pipe_phv_out_data_200; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_201 = proc_0_io_pipe_phv_out_data_201; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_202 = proc_0_io_pipe_phv_out_data_202; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_203 = proc_0_io_pipe_phv_out_data_203; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_204 = proc_0_io_pipe_phv_out_data_204; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_205 = proc_0_io_pipe_phv_out_data_205; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_206 = proc_0_io_pipe_phv_out_data_206; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_207 = proc_0_io_pipe_phv_out_data_207; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_208 = proc_0_io_pipe_phv_out_data_208; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_209 = proc_0_io_pipe_phv_out_data_209; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_210 = proc_0_io_pipe_phv_out_data_210; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_211 = proc_0_io_pipe_phv_out_data_211; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_212 = proc_0_io_pipe_phv_out_data_212; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_213 = proc_0_io_pipe_phv_out_data_213; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_214 = proc_0_io_pipe_phv_out_data_214; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_215 = proc_0_io_pipe_phv_out_data_215; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_216 = proc_0_io_pipe_phv_out_data_216; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_217 = proc_0_io_pipe_phv_out_data_217; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_218 = proc_0_io_pipe_phv_out_data_218; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_219 = proc_0_io_pipe_phv_out_data_219; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_220 = proc_0_io_pipe_phv_out_data_220; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_221 = proc_0_io_pipe_phv_out_data_221; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_222 = proc_0_io_pipe_phv_out_data_222; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_223 = proc_0_io_pipe_phv_out_data_223; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_224 = proc_0_io_pipe_phv_out_data_224; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_225 = proc_0_io_pipe_phv_out_data_225; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_226 = proc_0_io_pipe_phv_out_data_226; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_227 = proc_0_io_pipe_phv_out_data_227; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_228 = proc_0_io_pipe_phv_out_data_228; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_229 = proc_0_io_pipe_phv_out_data_229; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_230 = proc_0_io_pipe_phv_out_data_230; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_231 = proc_0_io_pipe_phv_out_data_231; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_232 = proc_0_io_pipe_phv_out_data_232; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_233 = proc_0_io_pipe_phv_out_data_233; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_234 = proc_0_io_pipe_phv_out_data_234; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_235 = proc_0_io_pipe_phv_out_data_235; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_236 = proc_0_io_pipe_phv_out_data_236; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_237 = proc_0_io_pipe_phv_out_data_237; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_238 = proc_0_io_pipe_phv_out_data_238; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_239 = proc_0_io_pipe_phv_out_data_239; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_240 = proc_0_io_pipe_phv_out_data_240; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_241 = proc_0_io_pipe_phv_out_data_241; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_242 = proc_0_io_pipe_phv_out_data_242; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_243 = proc_0_io_pipe_phv_out_data_243; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_244 = proc_0_io_pipe_phv_out_data_244; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_245 = proc_0_io_pipe_phv_out_data_245; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_246 = proc_0_io_pipe_phv_out_data_246; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_247 = proc_0_io_pipe_phv_out_data_247; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_248 = proc_0_io_pipe_phv_out_data_248; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_249 = proc_0_io_pipe_phv_out_data_249; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_250 = proc_0_io_pipe_phv_out_data_250; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_251 = proc_0_io_pipe_phv_out_data_251; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_252 = proc_0_io_pipe_phv_out_data_252; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_253 = proc_0_io_pipe_phv_out_data_253; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_254 = proc_0_io_pipe_phv_out_data_254; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_data_255 = proc_0_io_pipe_phv_out_data_255; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_header_0 = proc_0_io_pipe_phv_out_header_0; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_header_1 = proc_0_io_pipe_phv_out_header_1; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_header_2 = proc_0_io_pipe_phv_out_header_2; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_header_3 = proc_0_io_pipe_phv_out_header_3; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_header_4 = proc_0_io_pipe_phv_out_header_4; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_header_5 = proc_0_io_pipe_phv_out_header_5; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_header_6 = proc_0_io_pipe_phv_out_header_6; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_header_7 = proc_0_io_pipe_phv_out_header_7; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_header_8 = proc_0_io_pipe_phv_out_header_8; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_header_9 = proc_0_io_pipe_phv_out_header_9; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_header_10 = proc_0_io_pipe_phv_out_header_10; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_header_11 = proc_0_io_pipe_phv_out_header_11; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_header_12 = proc_0_io_pipe_phv_out_header_12; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_header_13 = proc_0_io_pipe_phv_out_header_13; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_header_14 = proc_0_io_pipe_phv_out_header_14; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_header_15 = proc_0_io_pipe_phv_out_header_15; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_parse_current_state = proc_0_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_parse_current_offset = proc_0_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_parse_transition_field = proc_0_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_next_processor_id = proc_0_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 88:32]
  assign trans_0_io_pipe_phv_in_next_config_id = proc_0_io_pipe_phv_out_next_config_id; // @[ipsa.scala 88:32]
  assign trans_0_io_next_proc_exist = last_proc_id != 2'h0; // @[ipsa.scala 86:48]
  assign trans_0_io_next_proc_id_in = next_proc_id_0; // @[ipsa.scala 87:32]
  assign trans_1_clock = clock;
  assign trans_1_io_pipe_phv_in_data_0 = proc_1_io_pipe_phv_out_data_0; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_1 = proc_1_io_pipe_phv_out_data_1; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_2 = proc_1_io_pipe_phv_out_data_2; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_3 = proc_1_io_pipe_phv_out_data_3; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_4 = proc_1_io_pipe_phv_out_data_4; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_5 = proc_1_io_pipe_phv_out_data_5; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_6 = proc_1_io_pipe_phv_out_data_6; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_7 = proc_1_io_pipe_phv_out_data_7; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_8 = proc_1_io_pipe_phv_out_data_8; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_9 = proc_1_io_pipe_phv_out_data_9; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_10 = proc_1_io_pipe_phv_out_data_10; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_11 = proc_1_io_pipe_phv_out_data_11; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_12 = proc_1_io_pipe_phv_out_data_12; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_13 = proc_1_io_pipe_phv_out_data_13; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_14 = proc_1_io_pipe_phv_out_data_14; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_15 = proc_1_io_pipe_phv_out_data_15; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_16 = proc_1_io_pipe_phv_out_data_16; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_17 = proc_1_io_pipe_phv_out_data_17; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_18 = proc_1_io_pipe_phv_out_data_18; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_19 = proc_1_io_pipe_phv_out_data_19; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_20 = proc_1_io_pipe_phv_out_data_20; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_21 = proc_1_io_pipe_phv_out_data_21; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_22 = proc_1_io_pipe_phv_out_data_22; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_23 = proc_1_io_pipe_phv_out_data_23; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_24 = proc_1_io_pipe_phv_out_data_24; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_25 = proc_1_io_pipe_phv_out_data_25; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_26 = proc_1_io_pipe_phv_out_data_26; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_27 = proc_1_io_pipe_phv_out_data_27; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_28 = proc_1_io_pipe_phv_out_data_28; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_29 = proc_1_io_pipe_phv_out_data_29; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_30 = proc_1_io_pipe_phv_out_data_30; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_31 = proc_1_io_pipe_phv_out_data_31; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_32 = proc_1_io_pipe_phv_out_data_32; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_33 = proc_1_io_pipe_phv_out_data_33; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_34 = proc_1_io_pipe_phv_out_data_34; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_35 = proc_1_io_pipe_phv_out_data_35; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_36 = proc_1_io_pipe_phv_out_data_36; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_37 = proc_1_io_pipe_phv_out_data_37; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_38 = proc_1_io_pipe_phv_out_data_38; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_39 = proc_1_io_pipe_phv_out_data_39; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_40 = proc_1_io_pipe_phv_out_data_40; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_41 = proc_1_io_pipe_phv_out_data_41; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_42 = proc_1_io_pipe_phv_out_data_42; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_43 = proc_1_io_pipe_phv_out_data_43; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_44 = proc_1_io_pipe_phv_out_data_44; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_45 = proc_1_io_pipe_phv_out_data_45; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_46 = proc_1_io_pipe_phv_out_data_46; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_47 = proc_1_io_pipe_phv_out_data_47; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_48 = proc_1_io_pipe_phv_out_data_48; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_49 = proc_1_io_pipe_phv_out_data_49; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_50 = proc_1_io_pipe_phv_out_data_50; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_51 = proc_1_io_pipe_phv_out_data_51; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_52 = proc_1_io_pipe_phv_out_data_52; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_53 = proc_1_io_pipe_phv_out_data_53; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_54 = proc_1_io_pipe_phv_out_data_54; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_55 = proc_1_io_pipe_phv_out_data_55; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_56 = proc_1_io_pipe_phv_out_data_56; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_57 = proc_1_io_pipe_phv_out_data_57; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_58 = proc_1_io_pipe_phv_out_data_58; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_59 = proc_1_io_pipe_phv_out_data_59; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_60 = proc_1_io_pipe_phv_out_data_60; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_61 = proc_1_io_pipe_phv_out_data_61; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_62 = proc_1_io_pipe_phv_out_data_62; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_63 = proc_1_io_pipe_phv_out_data_63; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_64 = proc_1_io_pipe_phv_out_data_64; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_65 = proc_1_io_pipe_phv_out_data_65; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_66 = proc_1_io_pipe_phv_out_data_66; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_67 = proc_1_io_pipe_phv_out_data_67; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_68 = proc_1_io_pipe_phv_out_data_68; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_69 = proc_1_io_pipe_phv_out_data_69; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_70 = proc_1_io_pipe_phv_out_data_70; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_71 = proc_1_io_pipe_phv_out_data_71; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_72 = proc_1_io_pipe_phv_out_data_72; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_73 = proc_1_io_pipe_phv_out_data_73; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_74 = proc_1_io_pipe_phv_out_data_74; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_75 = proc_1_io_pipe_phv_out_data_75; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_76 = proc_1_io_pipe_phv_out_data_76; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_77 = proc_1_io_pipe_phv_out_data_77; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_78 = proc_1_io_pipe_phv_out_data_78; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_79 = proc_1_io_pipe_phv_out_data_79; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_80 = proc_1_io_pipe_phv_out_data_80; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_81 = proc_1_io_pipe_phv_out_data_81; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_82 = proc_1_io_pipe_phv_out_data_82; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_83 = proc_1_io_pipe_phv_out_data_83; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_84 = proc_1_io_pipe_phv_out_data_84; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_85 = proc_1_io_pipe_phv_out_data_85; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_86 = proc_1_io_pipe_phv_out_data_86; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_87 = proc_1_io_pipe_phv_out_data_87; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_88 = proc_1_io_pipe_phv_out_data_88; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_89 = proc_1_io_pipe_phv_out_data_89; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_90 = proc_1_io_pipe_phv_out_data_90; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_91 = proc_1_io_pipe_phv_out_data_91; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_92 = proc_1_io_pipe_phv_out_data_92; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_93 = proc_1_io_pipe_phv_out_data_93; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_94 = proc_1_io_pipe_phv_out_data_94; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_95 = proc_1_io_pipe_phv_out_data_95; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_96 = proc_1_io_pipe_phv_out_data_96; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_97 = proc_1_io_pipe_phv_out_data_97; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_98 = proc_1_io_pipe_phv_out_data_98; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_99 = proc_1_io_pipe_phv_out_data_99; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_100 = proc_1_io_pipe_phv_out_data_100; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_101 = proc_1_io_pipe_phv_out_data_101; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_102 = proc_1_io_pipe_phv_out_data_102; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_103 = proc_1_io_pipe_phv_out_data_103; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_104 = proc_1_io_pipe_phv_out_data_104; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_105 = proc_1_io_pipe_phv_out_data_105; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_106 = proc_1_io_pipe_phv_out_data_106; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_107 = proc_1_io_pipe_phv_out_data_107; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_108 = proc_1_io_pipe_phv_out_data_108; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_109 = proc_1_io_pipe_phv_out_data_109; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_110 = proc_1_io_pipe_phv_out_data_110; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_111 = proc_1_io_pipe_phv_out_data_111; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_112 = proc_1_io_pipe_phv_out_data_112; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_113 = proc_1_io_pipe_phv_out_data_113; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_114 = proc_1_io_pipe_phv_out_data_114; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_115 = proc_1_io_pipe_phv_out_data_115; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_116 = proc_1_io_pipe_phv_out_data_116; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_117 = proc_1_io_pipe_phv_out_data_117; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_118 = proc_1_io_pipe_phv_out_data_118; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_119 = proc_1_io_pipe_phv_out_data_119; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_120 = proc_1_io_pipe_phv_out_data_120; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_121 = proc_1_io_pipe_phv_out_data_121; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_122 = proc_1_io_pipe_phv_out_data_122; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_123 = proc_1_io_pipe_phv_out_data_123; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_124 = proc_1_io_pipe_phv_out_data_124; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_125 = proc_1_io_pipe_phv_out_data_125; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_126 = proc_1_io_pipe_phv_out_data_126; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_127 = proc_1_io_pipe_phv_out_data_127; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_128 = proc_1_io_pipe_phv_out_data_128; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_129 = proc_1_io_pipe_phv_out_data_129; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_130 = proc_1_io_pipe_phv_out_data_130; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_131 = proc_1_io_pipe_phv_out_data_131; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_132 = proc_1_io_pipe_phv_out_data_132; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_133 = proc_1_io_pipe_phv_out_data_133; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_134 = proc_1_io_pipe_phv_out_data_134; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_135 = proc_1_io_pipe_phv_out_data_135; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_136 = proc_1_io_pipe_phv_out_data_136; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_137 = proc_1_io_pipe_phv_out_data_137; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_138 = proc_1_io_pipe_phv_out_data_138; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_139 = proc_1_io_pipe_phv_out_data_139; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_140 = proc_1_io_pipe_phv_out_data_140; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_141 = proc_1_io_pipe_phv_out_data_141; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_142 = proc_1_io_pipe_phv_out_data_142; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_143 = proc_1_io_pipe_phv_out_data_143; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_144 = proc_1_io_pipe_phv_out_data_144; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_145 = proc_1_io_pipe_phv_out_data_145; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_146 = proc_1_io_pipe_phv_out_data_146; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_147 = proc_1_io_pipe_phv_out_data_147; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_148 = proc_1_io_pipe_phv_out_data_148; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_149 = proc_1_io_pipe_phv_out_data_149; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_150 = proc_1_io_pipe_phv_out_data_150; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_151 = proc_1_io_pipe_phv_out_data_151; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_152 = proc_1_io_pipe_phv_out_data_152; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_153 = proc_1_io_pipe_phv_out_data_153; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_154 = proc_1_io_pipe_phv_out_data_154; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_155 = proc_1_io_pipe_phv_out_data_155; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_156 = proc_1_io_pipe_phv_out_data_156; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_157 = proc_1_io_pipe_phv_out_data_157; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_158 = proc_1_io_pipe_phv_out_data_158; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_159 = proc_1_io_pipe_phv_out_data_159; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_160 = proc_1_io_pipe_phv_out_data_160; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_161 = proc_1_io_pipe_phv_out_data_161; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_162 = proc_1_io_pipe_phv_out_data_162; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_163 = proc_1_io_pipe_phv_out_data_163; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_164 = proc_1_io_pipe_phv_out_data_164; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_165 = proc_1_io_pipe_phv_out_data_165; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_166 = proc_1_io_pipe_phv_out_data_166; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_167 = proc_1_io_pipe_phv_out_data_167; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_168 = proc_1_io_pipe_phv_out_data_168; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_169 = proc_1_io_pipe_phv_out_data_169; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_170 = proc_1_io_pipe_phv_out_data_170; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_171 = proc_1_io_pipe_phv_out_data_171; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_172 = proc_1_io_pipe_phv_out_data_172; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_173 = proc_1_io_pipe_phv_out_data_173; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_174 = proc_1_io_pipe_phv_out_data_174; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_175 = proc_1_io_pipe_phv_out_data_175; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_176 = proc_1_io_pipe_phv_out_data_176; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_177 = proc_1_io_pipe_phv_out_data_177; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_178 = proc_1_io_pipe_phv_out_data_178; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_179 = proc_1_io_pipe_phv_out_data_179; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_180 = proc_1_io_pipe_phv_out_data_180; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_181 = proc_1_io_pipe_phv_out_data_181; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_182 = proc_1_io_pipe_phv_out_data_182; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_183 = proc_1_io_pipe_phv_out_data_183; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_184 = proc_1_io_pipe_phv_out_data_184; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_185 = proc_1_io_pipe_phv_out_data_185; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_186 = proc_1_io_pipe_phv_out_data_186; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_187 = proc_1_io_pipe_phv_out_data_187; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_188 = proc_1_io_pipe_phv_out_data_188; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_189 = proc_1_io_pipe_phv_out_data_189; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_190 = proc_1_io_pipe_phv_out_data_190; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_191 = proc_1_io_pipe_phv_out_data_191; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_192 = proc_1_io_pipe_phv_out_data_192; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_193 = proc_1_io_pipe_phv_out_data_193; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_194 = proc_1_io_pipe_phv_out_data_194; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_195 = proc_1_io_pipe_phv_out_data_195; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_196 = proc_1_io_pipe_phv_out_data_196; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_197 = proc_1_io_pipe_phv_out_data_197; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_198 = proc_1_io_pipe_phv_out_data_198; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_199 = proc_1_io_pipe_phv_out_data_199; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_200 = proc_1_io_pipe_phv_out_data_200; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_201 = proc_1_io_pipe_phv_out_data_201; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_202 = proc_1_io_pipe_phv_out_data_202; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_203 = proc_1_io_pipe_phv_out_data_203; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_204 = proc_1_io_pipe_phv_out_data_204; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_205 = proc_1_io_pipe_phv_out_data_205; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_206 = proc_1_io_pipe_phv_out_data_206; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_207 = proc_1_io_pipe_phv_out_data_207; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_208 = proc_1_io_pipe_phv_out_data_208; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_209 = proc_1_io_pipe_phv_out_data_209; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_210 = proc_1_io_pipe_phv_out_data_210; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_211 = proc_1_io_pipe_phv_out_data_211; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_212 = proc_1_io_pipe_phv_out_data_212; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_213 = proc_1_io_pipe_phv_out_data_213; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_214 = proc_1_io_pipe_phv_out_data_214; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_215 = proc_1_io_pipe_phv_out_data_215; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_216 = proc_1_io_pipe_phv_out_data_216; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_217 = proc_1_io_pipe_phv_out_data_217; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_218 = proc_1_io_pipe_phv_out_data_218; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_219 = proc_1_io_pipe_phv_out_data_219; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_220 = proc_1_io_pipe_phv_out_data_220; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_221 = proc_1_io_pipe_phv_out_data_221; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_222 = proc_1_io_pipe_phv_out_data_222; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_223 = proc_1_io_pipe_phv_out_data_223; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_224 = proc_1_io_pipe_phv_out_data_224; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_225 = proc_1_io_pipe_phv_out_data_225; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_226 = proc_1_io_pipe_phv_out_data_226; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_227 = proc_1_io_pipe_phv_out_data_227; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_228 = proc_1_io_pipe_phv_out_data_228; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_229 = proc_1_io_pipe_phv_out_data_229; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_230 = proc_1_io_pipe_phv_out_data_230; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_231 = proc_1_io_pipe_phv_out_data_231; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_232 = proc_1_io_pipe_phv_out_data_232; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_233 = proc_1_io_pipe_phv_out_data_233; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_234 = proc_1_io_pipe_phv_out_data_234; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_235 = proc_1_io_pipe_phv_out_data_235; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_236 = proc_1_io_pipe_phv_out_data_236; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_237 = proc_1_io_pipe_phv_out_data_237; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_238 = proc_1_io_pipe_phv_out_data_238; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_239 = proc_1_io_pipe_phv_out_data_239; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_240 = proc_1_io_pipe_phv_out_data_240; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_241 = proc_1_io_pipe_phv_out_data_241; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_242 = proc_1_io_pipe_phv_out_data_242; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_243 = proc_1_io_pipe_phv_out_data_243; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_244 = proc_1_io_pipe_phv_out_data_244; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_245 = proc_1_io_pipe_phv_out_data_245; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_246 = proc_1_io_pipe_phv_out_data_246; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_247 = proc_1_io_pipe_phv_out_data_247; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_248 = proc_1_io_pipe_phv_out_data_248; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_249 = proc_1_io_pipe_phv_out_data_249; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_250 = proc_1_io_pipe_phv_out_data_250; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_251 = proc_1_io_pipe_phv_out_data_251; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_252 = proc_1_io_pipe_phv_out_data_252; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_253 = proc_1_io_pipe_phv_out_data_253; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_254 = proc_1_io_pipe_phv_out_data_254; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_data_255 = proc_1_io_pipe_phv_out_data_255; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_header_0 = proc_1_io_pipe_phv_out_header_0; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_header_1 = proc_1_io_pipe_phv_out_header_1; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_header_2 = proc_1_io_pipe_phv_out_header_2; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_header_3 = proc_1_io_pipe_phv_out_header_3; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_header_4 = proc_1_io_pipe_phv_out_header_4; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_header_5 = proc_1_io_pipe_phv_out_header_5; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_header_6 = proc_1_io_pipe_phv_out_header_6; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_header_7 = proc_1_io_pipe_phv_out_header_7; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_header_8 = proc_1_io_pipe_phv_out_header_8; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_header_9 = proc_1_io_pipe_phv_out_header_9; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_header_10 = proc_1_io_pipe_phv_out_header_10; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_header_11 = proc_1_io_pipe_phv_out_header_11; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_header_12 = proc_1_io_pipe_phv_out_header_12; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_header_13 = proc_1_io_pipe_phv_out_header_13; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_header_14 = proc_1_io_pipe_phv_out_header_14; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_header_15 = proc_1_io_pipe_phv_out_header_15; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_parse_current_state = proc_1_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_parse_current_offset = proc_1_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_parse_transition_field = proc_1_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_next_processor_id = proc_1_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 88:32]
  assign trans_1_io_pipe_phv_in_next_config_id = proc_1_io_pipe_phv_out_next_config_id; // @[ipsa.scala 88:32]
  assign trans_1_io_next_proc_exist = last_proc_id != 2'h1; // @[ipsa.scala 86:48]
  assign trans_1_io_next_proc_id_in = next_proc_id_1; // @[ipsa.scala 87:32]
  assign trans_2_clock = clock;
  assign trans_2_io_pipe_phv_in_data_0 = proc_2_io_pipe_phv_out_data_0; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_1 = proc_2_io_pipe_phv_out_data_1; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_2 = proc_2_io_pipe_phv_out_data_2; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_3 = proc_2_io_pipe_phv_out_data_3; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_4 = proc_2_io_pipe_phv_out_data_4; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_5 = proc_2_io_pipe_phv_out_data_5; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_6 = proc_2_io_pipe_phv_out_data_6; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_7 = proc_2_io_pipe_phv_out_data_7; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_8 = proc_2_io_pipe_phv_out_data_8; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_9 = proc_2_io_pipe_phv_out_data_9; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_10 = proc_2_io_pipe_phv_out_data_10; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_11 = proc_2_io_pipe_phv_out_data_11; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_12 = proc_2_io_pipe_phv_out_data_12; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_13 = proc_2_io_pipe_phv_out_data_13; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_14 = proc_2_io_pipe_phv_out_data_14; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_15 = proc_2_io_pipe_phv_out_data_15; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_16 = proc_2_io_pipe_phv_out_data_16; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_17 = proc_2_io_pipe_phv_out_data_17; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_18 = proc_2_io_pipe_phv_out_data_18; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_19 = proc_2_io_pipe_phv_out_data_19; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_20 = proc_2_io_pipe_phv_out_data_20; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_21 = proc_2_io_pipe_phv_out_data_21; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_22 = proc_2_io_pipe_phv_out_data_22; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_23 = proc_2_io_pipe_phv_out_data_23; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_24 = proc_2_io_pipe_phv_out_data_24; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_25 = proc_2_io_pipe_phv_out_data_25; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_26 = proc_2_io_pipe_phv_out_data_26; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_27 = proc_2_io_pipe_phv_out_data_27; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_28 = proc_2_io_pipe_phv_out_data_28; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_29 = proc_2_io_pipe_phv_out_data_29; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_30 = proc_2_io_pipe_phv_out_data_30; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_31 = proc_2_io_pipe_phv_out_data_31; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_32 = proc_2_io_pipe_phv_out_data_32; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_33 = proc_2_io_pipe_phv_out_data_33; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_34 = proc_2_io_pipe_phv_out_data_34; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_35 = proc_2_io_pipe_phv_out_data_35; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_36 = proc_2_io_pipe_phv_out_data_36; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_37 = proc_2_io_pipe_phv_out_data_37; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_38 = proc_2_io_pipe_phv_out_data_38; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_39 = proc_2_io_pipe_phv_out_data_39; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_40 = proc_2_io_pipe_phv_out_data_40; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_41 = proc_2_io_pipe_phv_out_data_41; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_42 = proc_2_io_pipe_phv_out_data_42; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_43 = proc_2_io_pipe_phv_out_data_43; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_44 = proc_2_io_pipe_phv_out_data_44; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_45 = proc_2_io_pipe_phv_out_data_45; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_46 = proc_2_io_pipe_phv_out_data_46; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_47 = proc_2_io_pipe_phv_out_data_47; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_48 = proc_2_io_pipe_phv_out_data_48; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_49 = proc_2_io_pipe_phv_out_data_49; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_50 = proc_2_io_pipe_phv_out_data_50; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_51 = proc_2_io_pipe_phv_out_data_51; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_52 = proc_2_io_pipe_phv_out_data_52; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_53 = proc_2_io_pipe_phv_out_data_53; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_54 = proc_2_io_pipe_phv_out_data_54; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_55 = proc_2_io_pipe_phv_out_data_55; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_56 = proc_2_io_pipe_phv_out_data_56; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_57 = proc_2_io_pipe_phv_out_data_57; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_58 = proc_2_io_pipe_phv_out_data_58; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_59 = proc_2_io_pipe_phv_out_data_59; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_60 = proc_2_io_pipe_phv_out_data_60; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_61 = proc_2_io_pipe_phv_out_data_61; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_62 = proc_2_io_pipe_phv_out_data_62; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_63 = proc_2_io_pipe_phv_out_data_63; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_64 = proc_2_io_pipe_phv_out_data_64; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_65 = proc_2_io_pipe_phv_out_data_65; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_66 = proc_2_io_pipe_phv_out_data_66; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_67 = proc_2_io_pipe_phv_out_data_67; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_68 = proc_2_io_pipe_phv_out_data_68; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_69 = proc_2_io_pipe_phv_out_data_69; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_70 = proc_2_io_pipe_phv_out_data_70; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_71 = proc_2_io_pipe_phv_out_data_71; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_72 = proc_2_io_pipe_phv_out_data_72; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_73 = proc_2_io_pipe_phv_out_data_73; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_74 = proc_2_io_pipe_phv_out_data_74; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_75 = proc_2_io_pipe_phv_out_data_75; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_76 = proc_2_io_pipe_phv_out_data_76; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_77 = proc_2_io_pipe_phv_out_data_77; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_78 = proc_2_io_pipe_phv_out_data_78; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_79 = proc_2_io_pipe_phv_out_data_79; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_80 = proc_2_io_pipe_phv_out_data_80; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_81 = proc_2_io_pipe_phv_out_data_81; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_82 = proc_2_io_pipe_phv_out_data_82; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_83 = proc_2_io_pipe_phv_out_data_83; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_84 = proc_2_io_pipe_phv_out_data_84; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_85 = proc_2_io_pipe_phv_out_data_85; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_86 = proc_2_io_pipe_phv_out_data_86; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_87 = proc_2_io_pipe_phv_out_data_87; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_88 = proc_2_io_pipe_phv_out_data_88; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_89 = proc_2_io_pipe_phv_out_data_89; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_90 = proc_2_io_pipe_phv_out_data_90; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_91 = proc_2_io_pipe_phv_out_data_91; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_92 = proc_2_io_pipe_phv_out_data_92; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_93 = proc_2_io_pipe_phv_out_data_93; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_94 = proc_2_io_pipe_phv_out_data_94; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_95 = proc_2_io_pipe_phv_out_data_95; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_96 = proc_2_io_pipe_phv_out_data_96; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_97 = proc_2_io_pipe_phv_out_data_97; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_98 = proc_2_io_pipe_phv_out_data_98; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_99 = proc_2_io_pipe_phv_out_data_99; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_100 = proc_2_io_pipe_phv_out_data_100; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_101 = proc_2_io_pipe_phv_out_data_101; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_102 = proc_2_io_pipe_phv_out_data_102; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_103 = proc_2_io_pipe_phv_out_data_103; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_104 = proc_2_io_pipe_phv_out_data_104; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_105 = proc_2_io_pipe_phv_out_data_105; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_106 = proc_2_io_pipe_phv_out_data_106; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_107 = proc_2_io_pipe_phv_out_data_107; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_108 = proc_2_io_pipe_phv_out_data_108; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_109 = proc_2_io_pipe_phv_out_data_109; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_110 = proc_2_io_pipe_phv_out_data_110; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_111 = proc_2_io_pipe_phv_out_data_111; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_112 = proc_2_io_pipe_phv_out_data_112; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_113 = proc_2_io_pipe_phv_out_data_113; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_114 = proc_2_io_pipe_phv_out_data_114; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_115 = proc_2_io_pipe_phv_out_data_115; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_116 = proc_2_io_pipe_phv_out_data_116; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_117 = proc_2_io_pipe_phv_out_data_117; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_118 = proc_2_io_pipe_phv_out_data_118; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_119 = proc_2_io_pipe_phv_out_data_119; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_120 = proc_2_io_pipe_phv_out_data_120; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_121 = proc_2_io_pipe_phv_out_data_121; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_122 = proc_2_io_pipe_phv_out_data_122; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_123 = proc_2_io_pipe_phv_out_data_123; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_124 = proc_2_io_pipe_phv_out_data_124; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_125 = proc_2_io_pipe_phv_out_data_125; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_126 = proc_2_io_pipe_phv_out_data_126; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_127 = proc_2_io_pipe_phv_out_data_127; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_128 = proc_2_io_pipe_phv_out_data_128; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_129 = proc_2_io_pipe_phv_out_data_129; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_130 = proc_2_io_pipe_phv_out_data_130; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_131 = proc_2_io_pipe_phv_out_data_131; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_132 = proc_2_io_pipe_phv_out_data_132; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_133 = proc_2_io_pipe_phv_out_data_133; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_134 = proc_2_io_pipe_phv_out_data_134; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_135 = proc_2_io_pipe_phv_out_data_135; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_136 = proc_2_io_pipe_phv_out_data_136; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_137 = proc_2_io_pipe_phv_out_data_137; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_138 = proc_2_io_pipe_phv_out_data_138; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_139 = proc_2_io_pipe_phv_out_data_139; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_140 = proc_2_io_pipe_phv_out_data_140; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_141 = proc_2_io_pipe_phv_out_data_141; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_142 = proc_2_io_pipe_phv_out_data_142; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_143 = proc_2_io_pipe_phv_out_data_143; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_144 = proc_2_io_pipe_phv_out_data_144; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_145 = proc_2_io_pipe_phv_out_data_145; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_146 = proc_2_io_pipe_phv_out_data_146; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_147 = proc_2_io_pipe_phv_out_data_147; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_148 = proc_2_io_pipe_phv_out_data_148; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_149 = proc_2_io_pipe_phv_out_data_149; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_150 = proc_2_io_pipe_phv_out_data_150; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_151 = proc_2_io_pipe_phv_out_data_151; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_152 = proc_2_io_pipe_phv_out_data_152; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_153 = proc_2_io_pipe_phv_out_data_153; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_154 = proc_2_io_pipe_phv_out_data_154; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_155 = proc_2_io_pipe_phv_out_data_155; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_156 = proc_2_io_pipe_phv_out_data_156; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_157 = proc_2_io_pipe_phv_out_data_157; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_158 = proc_2_io_pipe_phv_out_data_158; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_159 = proc_2_io_pipe_phv_out_data_159; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_160 = proc_2_io_pipe_phv_out_data_160; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_161 = proc_2_io_pipe_phv_out_data_161; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_162 = proc_2_io_pipe_phv_out_data_162; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_163 = proc_2_io_pipe_phv_out_data_163; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_164 = proc_2_io_pipe_phv_out_data_164; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_165 = proc_2_io_pipe_phv_out_data_165; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_166 = proc_2_io_pipe_phv_out_data_166; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_167 = proc_2_io_pipe_phv_out_data_167; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_168 = proc_2_io_pipe_phv_out_data_168; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_169 = proc_2_io_pipe_phv_out_data_169; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_170 = proc_2_io_pipe_phv_out_data_170; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_171 = proc_2_io_pipe_phv_out_data_171; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_172 = proc_2_io_pipe_phv_out_data_172; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_173 = proc_2_io_pipe_phv_out_data_173; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_174 = proc_2_io_pipe_phv_out_data_174; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_175 = proc_2_io_pipe_phv_out_data_175; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_176 = proc_2_io_pipe_phv_out_data_176; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_177 = proc_2_io_pipe_phv_out_data_177; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_178 = proc_2_io_pipe_phv_out_data_178; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_179 = proc_2_io_pipe_phv_out_data_179; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_180 = proc_2_io_pipe_phv_out_data_180; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_181 = proc_2_io_pipe_phv_out_data_181; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_182 = proc_2_io_pipe_phv_out_data_182; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_183 = proc_2_io_pipe_phv_out_data_183; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_184 = proc_2_io_pipe_phv_out_data_184; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_185 = proc_2_io_pipe_phv_out_data_185; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_186 = proc_2_io_pipe_phv_out_data_186; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_187 = proc_2_io_pipe_phv_out_data_187; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_188 = proc_2_io_pipe_phv_out_data_188; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_189 = proc_2_io_pipe_phv_out_data_189; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_190 = proc_2_io_pipe_phv_out_data_190; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_191 = proc_2_io_pipe_phv_out_data_191; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_192 = proc_2_io_pipe_phv_out_data_192; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_193 = proc_2_io_pipe_phv_out_data_193; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_194 = proc_2_io_pipe_phv_out_data_194; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_195 = proc_2_io_pipe_phv_out_data_195; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_196 = proc_2_io_pipe_phv_out_data_196; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_197 = proc_2_io_pipe_phv_out_data_197; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_198 = proc_2_io_pipe_phv_out_data_198; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_199 = proc_2_io_pipe_phv_out_data_199; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_200 = proc_2_io_pipe_phv_out_data_200; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_201 = proc_2_io_pipe_phv_out_data_201; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_202 = proc_2_io_pipe_phv_out_data_202; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_203 = proc_2_io_pipe_phv_out_data_203; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_204 = proc_2_io_pipe_phv_out_data_204; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_205 = proc_2_io_pipe_phv_out_data_205; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_206 = proc_2_io_pipe_phv_out_data_206; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_207 = proc_2_io_pipe_phv_out_data_207; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_208 = proc_2_io_pipe_phv_out_data_208; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_209 = proc_2_io_pipe_phv_out_data_209; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_210 = proc_2_io_pipe_phv_out_data_210; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_211 = proc_2_io_pipe_phv_out_data_211; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_212 = proc_2_io_pipe_phv_out_data_212; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_213 = proc_2_io_pipe_phv_out_data_213; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_214 = proc_2_io_pipe_phv_out_data_214; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_215 = proc_2_io_pipe_phv_out_data_215; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_216 = proc_2_io_pipe_phv_out_data_216; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_217 = proc_2_io_pipe_phv_out_data_217; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_218 = proc_2_io_pipe_phv_out_data_218; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_219 = proc_2_io_pipe_phv_out_data_219; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_220 = proc_2_io_pipe_phv_out_data_220; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_221 = proc_2_io_pipe_phv_out_data_221; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_222 = proc_2_io_pipe_phv_out_data_222; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_223 = proc_2_io_pipe_phv_out_data_223; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_224 = proc_2_io_pipe_phv_out_data_224; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_225 = proc_2_io_pipe_phv_out_data_225; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_226 = proc_2_io_pipe_phv_out_data_226; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_227 = proc_2_io_pipe_phv_out_data_227; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_228 = proc_2_io_pipe_phv_out_data_228; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_229 = proc_2_io_pipe_phv_out_data_229; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_230 = proc_2_io_pipe_phv_out_data_230; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_231 = proc_2_io_pipe_phv_out_data_231; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_232 = proc_2_io_pipe_phv_out_data_232; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_233 = proc_2_io_pipe_phv_out_data_233; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_234 = proc_2_io_pipe_phv_out_data_234; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_235 = proc_2_io_pipe_phv_out_data_235; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_236 = proc_2_io_pipe_phv_out_data_236; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_237 = proc_2_io_pipe_phv_out_data_237; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_238 = proc_2_io_pipe_phv_out_data_238; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_239 = proc_2_io_pipe_phv_out_data_239; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_240 = proc_2_io_pipe_phv_out_data_240; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_241 = proc_2_io_pipe_phv_out_data_241; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_242 = proc_2_io_pipe_phv_out_data_242; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_243 = proc_2_io_pipe_phv_out_data_243; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_244 = proc_2_io_pipe_phv_out_data_244; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_245 = proc_2_io_pipe_phv_out_data_245; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_246 = proc_2_io_pipe_phv_out_data_246; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_247 = proc_2_io_pipe_phv_out_data_247; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_248 = proc_2_io_pipe_phv_out_data_248; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_249 = proc_2_io_pipe_phv_out_data_249; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_250 = proc_2_io_pipe_phv_out_data_250; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_251 = proc_2_io_pipe_phv_out_data_251; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_252 = proc_2_io_pipe_phv_out_data_252; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_253 = proc_2_io_pipe_phv_out_data_253; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_254 = proc_2_io_pipe_phv_out_data_254; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_data_255 = proc_2_io_pipe_phv_out_data_255; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_header_0 = proc_2_io_pipe_phv_out_header_0; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_header_1 = proc_2_io_pipe_phv_out_header_1; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_header_2 = proc_2_io_pipe_phv_out_header_2; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_header_3 = proc_2_io_pipe_phv_out_header_3; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_header_4 = proc_2_io_pipe_phv_out_header_4; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_header_5 = proc_2_io_pipe_phv_out_header_5; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_header_6 = proc_2_io_pipe_phv_out_header_6; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_header_7 = proc_2_io_pipe_phv_out_header_7; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_header_8 = proc_2_io_pipe_phv_out_header_8; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_header_9 = proc_2_io_pipe_phv_out_header_9; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_header_10 = proc_2_io_pipe_phv_out_header_10; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_header_11 = proc_2_io_pipe_phv_out_header_11; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_header_12 = proc_2_io_pipe_phv_out_header_12; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_header_13 = proc_2_io_pipe_phv_out_header_13; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_header_14 = proc_2_io_pipe_phv_out_header_14; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_header_15 = proc_2_io_pipe_phv_out_header_15; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_parse_current_state = proc_2_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_parse_current_offset = proc_2_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_parse_transition_field = proc_2_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_next_processor_id = proc_2_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 88:32]
  assign trans_2_io_pipe_phv_in_next_config_id = proc_2_io_pipe_phv_out_next_config_id; // @[ipsa.scala 88:32]
  assign trans_2_io_next_proc_exist = last_proc_id != 2'h2; // @[ipsa.scala 86:48]
  assign trans_2_io_next_proc_id_in = next_proc_id_2; // @[ipsa.scala 87:32]
  assign trans_3_clock = clock;
  assign trans_3_io_pipe_phv_in_data_0 = proc_3_io_pipe_phv_out_data_0; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_1 = proc_3_io_pipe_phv_out_data_1; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_2 = proc_3_io_pipe_phv_out_data_2; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_3 = proc_3_io_pipe_phv_out_data_3; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_4 = proc_3_io_pipe_phv_out_data_4; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_5 = proc_3_io_pipe_phv_out_data_5; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_6 = proc_3_io_pipe_phv_out_data_6; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_7 = proc_3_io_pipe_phv_out_data_7; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_8 = proc_3_io_pipe_phv_out_data_8; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_9 = proc_3_io_pipe_phv_out_data_9; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_10 = proc_3_io_pipe_phv_out_data_10; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_11 = proc_3_io_pipe_phv_out_data_11; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_12 = proc_3_io_pipe_phv_out_data_12; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_13 = proc_3_io_pipe_phv_out_data_13; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_14 = proc_3_io_pipe_phv_out_data_14; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_15 = proc_3_io_pipe_phv_out_data_15; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_16 = proc_3_io_pipe_phv_out_data_16; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_17 = proc_3_io_pipe_phv_out_data_17; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_18 = proc_3_io_pipe_phv_out_data_18; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_19 = proc_3_io_pipe_phv_out_data_19; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_20 = proc_3_io_pipe_phv_out_data_20; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_21 = proc_3_io_pipe_phv_out_data_21; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_22 = proc_3_io_pipe_phv_out_data_22; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_23 = proc_3_io_pipe_phv_out_data_23; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_24 = proc_3_io_pipe_phv_out_data_24; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_25 = proc_3_io_pipe_phv_out_data_25; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_26 = proc_3_io_pipe_phv_out_data_26; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_27 = proc_3_io_pipe_phv_out_data_27; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_28 = proc_3_io_pipe_phv_out_data_28; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_29 = proc_3_io_pipe_phv_out_data_29; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_30 = proc_3_io_pipe_phv_out_data_30; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_31 = proc_3_io_pipe_phv_out_data_31; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_32 = proc_3_io_pipe_phv_out_data_32; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_33 = proc_3_io_pipe_phv_out_data_33; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_34 = proc_3_io_pipe_phv_out_data_34; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_35 = proc_3_io_pipe_phv_out_data_35; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_36 = proc_3_io_pipe_phv_out_data_36; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_37 = proc_3_io_pipe_phv_out_data_37; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_38 = proc_3_io_pipe_phv_out_data_38; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_39 = proc_3_io_pipe_phv_out_data_39; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_40 = proc_3_io_pipe_phv_out_data_40; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_41 = proc_3_io_pipe_phv_out_data_41; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_42 = proc_3_io_pipe_phv_out_data_42; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_43 = proc_3_io_pipe_phv_out_data_43; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_44 = proc_3_io_pipe_phv_out_data_44; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_45 = proc_3_io_pipe_phv_out_data_45; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_46 = proc_3_io_pipe_phv_out_data_46; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_47 = proc_3_io_pipe_phv_out_data_47; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_48 = proc_3_io_pipe_phv_out_data_48; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_49 = proc_3_io_pipe_phv_out_data_49; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_50 = proc_3_io_pipe_phv_out_data_50; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_51 = proc_3_io_pipe_phv_out_data_51; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_52 = proc_3_io_pipe_phv_out_data_52; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_53 = proc_3_io_pipe_phv_out_data_53; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_54 = proc_3_io_pipe_phv_out_data_54; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_55 = proc_3_io_pipe_phv_out_data_55; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_56 = proc_3_io_pipe_phv_out_data_56; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_57 = proc_3_io_pipe_phv_out_data_57; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_58 = proc_3_io_pipe_phv_out_data_58; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_59 = proc_3_io_pipe_phv_out_data_59; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_60 = proc_3_io_pipe_phv_out_data_60; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_61 = proc_3_io_pipe_phv_out_data_61; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_62 = proc_3_io_pipe_phv_out_data_62; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_63 = proc_3_io_pipe_phv_out_data_63; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_64 = proc_3_io_pipe_phv_out_data_64; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_65 = proc_3_io_pipe_phv_out_data_65; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_66 = proc_3_io_pipe_phv_out_data_66; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_67 = proc_3_io_pipe_phv_out_data_67; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_68 = proc_3_io_pipe_phv_out_data_68; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_69 = proc_3_io_pipe_phv_out_data_69; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_70 = proc_3_io_pipe_phv_out_data_70; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_71 = proc_3_io_pipe_phv_out_data_71; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_72 = proc_3_io_pipe_phv_out_data_72; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_73 = proc_3_io_pipe_phv_out_data_73; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_74 = proc_3_io_pipe_phv_out_data_74; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_75 = proc_3_io_pipe_phv_out_data_75; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_76 = proc_3_io_pipe_phv_out_data_76; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_77 = proc_3_io_pipe_phv_out_data_77; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_78 = proc_3_io_pipe_phv_out_data_78; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_79 = proc_3_io_pipe_phv_out_data_79; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_80 = proc_3_io_pipe_phv_out_data_80; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_81 = proc_3_io_pipe_phv_out_data_81; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_82 = proc_3_io_pipe_phv_out_data_82; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_83 = proc_3_io_pipe_phv_out_data_83; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_84 = proc_3_io_pipe_phv_out_data_84; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_85 = proc_3_io_pipe_phv_out_data_85; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_86 = proc_3_io_pipe_phv_out_data_86; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_87 = proc_3_io_pipe_phv_out_data_87; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_88 = proc_3_io_pipe_phv_out_data_88; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_89 = proc_3_io_pipe_phv_out_data_89; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_90 = proc_3_io_pipe_phv_out_data_90; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_91 = proc_3_io_pipe_phv_out_data_91; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_92 = proc_3_io_pipe_phv_out_data_92; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_93 = proc_3_io_pipe_phv_out_data_93; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_94 = proc_3_io_pipe_phv_out_data_94; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_95 = proc_3_io_pipe_phv_out_data_95; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_96 = proc_3_io_pipe_phv_out_data_96; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_97 = proc_3_io_pipe_phv_out_data_97; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_98 = proc_3_io_pipe_phv_out_data_98; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_99 = proc_3_io_pipe_phv_out_data_99; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_100 = proc_3_io_pipe_phv_out_data_100; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_101 = proc_3_io_pipe_phv_out_data_101; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_102 = proc_3_io_pipe_phv_out_data_102; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_103 = proc_3_io_pipe_phv_out_data_103; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_104 = proc_3_io_pipe_phv_out_data_104; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_105 = proc_3_io_pipe_phv_out_data_105; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_106 = proc_3_io_pipe_phv_out_data_106; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_107 = proc_3_io_pipe_phv_out_data_107; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_108 = proc_3_io_pipe_phv_out_data_108; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_109 = proc_3_io_pipe_phv_out_data_109; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_110 = proc_3_io_pipe_phv_out_data_110; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_111 = proc_3_io_pipe_phv_out_data_111; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_112 = proc_3_io_pipe_phv_out_data_112; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_113 = proc_3_io_pipe_phv_out_data_113; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_114 = proc_3_io_pipe_phv_out_data_114; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_115 = proc_3_io_pipe_phv_out_data_115; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_116 = proc_3_io_pipe_phv_out_data_116; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_117 = proc_3_io_pipe_phv_out_data_117; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_118 = proc_3_io_pipe_phv_out_data_118; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_119 = proc_3_io_pipe_phv_out_data_119; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_120 = proc_3_io_pipe_phv_out_data_120; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_121 = proc_3_io_pipe_phv_out_data_121; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_122 = proc_3_io_pipe_phv_out_data_122; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_123 = proc_3_io_pipe_phv_out_data_123; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_124 = proc_3_io_pipe_phv_out_data_124; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_125 = proc_3_io_pipe_phv_out_data_125; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_126 = proc_3_io_pipe_phv_out_data_126; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_127 = proc_3_io_pipe_phv_out_data_127; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_128 = proc_3_io_pipe_phv_out_data_128; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_129 = proc_3_io_pipe_phv_out_data_129; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_130 = proc_3_io_pipe_phv_out_data_130; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_131 = proc_3_io_pipe_phv_out_data_131; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_132 = proc_3_io_pipe_phv_out_data_132; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_133 = proc_3_io_pipe_phv_out_data_133; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_134 = proc_3_io_pipe_phv_out_data_134; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_135 = proc_3_io_pipe_phv_out_data_135; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_136 = proc_3_io_pipe_phv_out_data_136; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_137 = proc_3_io_pipe_phv_out_data_137; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_138 = proc_3_io_pipe_phv_out_data_138; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_139 = proc_3_io_pipe_phv_out_data_139; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_140 = proc_3_io_pipe_phv_out_data_140; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_141 = proc_3_io_pipe_phv_out_data_141; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_142 = proc_3_io_pipe_phv_out_data_142; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_143 = proc_3_io_pipe_phv_out_data_143; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_144 = proc_3_io_pipe_phv_out_data_144; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_145 = proc_3_io_pipe_phv_out_data_145; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_146 = proc_3_io_pipe_phv_out_data_146; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_147 = proc_3_io_pipe_phv_out_data_147; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_148 = proc_3_io_pipe_phv_out_data_148; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_149 = proc_3_io_pipe_phv_out_data_149; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_150 = proc_3_io_pipe_phv_out_data_150; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_151 = proc_3_io_pipe_phv_out_data_151; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_152 = proc_3_io_pipe_phv_out_data_152; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_153 = proc_3_io_pipe_phv_out_data_153; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_154 = proc_3_io_pipe_phv_out_data_154; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_155 = proc_3_io_pipe_phv_out_data_155; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_156 = proc_3_io_pipe_phv_out_data_156; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_157 = proc_3_io_pipe_phv_out_data_157; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_158 = proc_3_io_pipe_phv_out_data_158; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_159 = proc_3_io_pipe_phv_out_data_159; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_160 = proc_3_io_pipe_phv_out_data_160; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_161 = proc_3_io_pipe_phv_out_data_161; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_162 = proc_3_io_pipe_phv_out_data_162; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_163 = proc_3_io_pipe_phv_out_data_163; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_164 = proc_3_io_pipe_phv_out_data_164; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_165 = proc_3_io_pipe_phv_out_data_165; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_166 = proc_3_io_pipe_phv_out_data_166; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_167 = proc_3_io_pipe_phv_out_data_167; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_168 = proc_3_io_pipe_phv_out_data_168; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_169 = proc_3_io_pipe_phv_out_data_169; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_170 = proc_3_io_pipe_phv_out_data_170; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_171 = proc_3_io_pipe_phv_out_data_171; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_172 = proc_3_io_pipe_phv_out_data_172; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_173 = proc_3_io_pipe_phv_out_data_173; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_174 = proc_3_io_pipe_phv_out_data_174; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_175 = proc_3_io_pipe_phv_out_data_175; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_176 = proc_3_io_pipe_phv_out_data_176; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_177 = proc_3_io_pipe_phv_out_data_177; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_178 = proc_3_io_pipe_phv_out_data_178; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_179 = proc_3_io_pipe_phv_out_data_179; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_180 = proc_3_io_pipe_phv_out_data_180; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_181 = proc_3_io_pipe_phv_out_data_181; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_182 = proc_3_io_pipe_phv_out_data_182; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_183 = proc_3_io_pipe_phv_out_data_183; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_184 = proc_3_io_pipe_phv_out_data_184; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_185 = proc_3_io_pipe_phv_out_data_185; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_186 = proc_3_io_pipe_phv_out_data_186; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_187 = proc_3_io_pipe_phv_out_data_187; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_188 = proc_3_io_pipe_phv_out_data_188; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_189 = proc_3_io_pipe_phv_out_data_189; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_190 = proc_3_io_pipe_phv_out_data_190; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_191 = proc_3_io_pipe_phv_out_data_191; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_192 = proc_3_io_pipe_phv_out_data_192; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_193 = proc_3_io_pipe_phv_out_data_193; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_194 = proc_3_io_pipe_phv_out_data_194; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_195 = proc_3_io_pipe_phv_out_data_195; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_196 = proc_3_io_pipe_phv_out_data_196; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_197 = proc_3_io_pipe_phv_out_data_197; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_198 = proc_3_io_pipe_phv_out_data_198; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_199 = proc_3_io_pipe_phv_out_data_199; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_200 = proc_3_io_pipe_phv_out_data_200; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_201 = proc_3_io_pipe_phv_out_data_201; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_202 = proc_3_io_pipe_phv_out_data_202; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_203 = proc_3_io_pipe_phv_out_data_203; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_204 = proc_3_io_pipe_phv_out_data_204; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_205 = proc_3_io_pipe_phv_out_data_205; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_206 = proc_3_io_pipe_phv_out_data_206; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_207 = proc_3_io_pipe_phv_out_data_207; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_208 = proc_3_io_pipe_phv_out_data_208; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_209 = proc_3_io_pipe_phv_out_data_209; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_210 = proc_3_io_pipe_phv_out_data_210; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_211 = proc_3_io_pipe_phv_out_data_211; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_212 = proc_3_io_pipe_phv_out_data_212; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_213 = proc_3_io_pipe_phv_out_data_213; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_214 = proc_3_io_pipe_phv_out_data_214; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_215 = proc_3_io_pipe_phv_out_data_215; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_216 = proc_3_io_pipe_phv_out_data_216; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_217 = proc_3_io_pipe_phv_out_data_217; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_218 = proc_3_io_pipe_phv_out_data_218; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_219 = proc_3_io_pipe_phv_out_data_219; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_220 = proc_3_io_pipe_phv_out_data_220; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_221 = proc_3_io_pipe_phv_out_data_221; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_222 = proc_3_io_pipe_phv_out_data_222; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_223 = proc_3_io_pipe_phv_out_data_223; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_224 = proc_3_io_pipe_phv_out_data_224; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_225 = proc_3_io_pipe_phv_out_data_225; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_226 = proc_3_io_pipe_phv_out_data_226; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_227 = proc_3_io_pipe_phv_out_data_227; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_228 = proc_3_io_pipe_phv_out_data_228; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_229 = proc_3_io_pipe_phv_out_data_229; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_230 = proc_3_io_pipe_phv_out_data_230; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_231 = proc_3_io_pipe_phv_out_data_231; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_232 = proc_3_io_pipe_phv_out_data_232; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_233 = proc_3_io_pipe_phv_out_data_233; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_234 = proc_3_io_pipe_phv_out_data_234; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_235 = proc_3_io_pipe_phv_out_data_235; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_236 = proc_3_io_pipe_phv_out_data_236; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_237 = proc_3_io_pipe_phv_out_data_237; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_238 = proc_3_io_pipe_phv_out_data_238; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_239 = proc_3_io_pipe_phv_out_data_239; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_240 = proc_3_io_pipe_phv_out_data_240; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_241 = proc_3_io_pipe_phv_out_data_241; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_242 = proc_3_io_pipe_phv_out_data_242; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_243 = proc_3_io_pipe_phv_out_data_243; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_244 = proc_3_io_pipe_phv_out_data_244; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_245 = proc_3_io_pipe_phv_out_data_245; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_246 = proc_3_io_pipe_phv_out_data_246; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_247 = proc_3_io_pipe_phv_out_data_247; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_248 = proc_3_io_pipe_phv_out_data_248; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_249 = proc_3_io_pipe_phv_out_data_249; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_250 = proc_3_io_pipe_phv_out_data_250; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_251 = proc_3_io_pipe_phv_out_data_251; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_252 = proc_3_io_pipe_phv_out_data_252; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_253 = proc_3_io_pipe_phv_out_data_253; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_254 = proc_3_io_pipe_phv_out_data_254; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_data_255 = proc_3_io_pipe_phv_out_data_255; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_header_0 = proc_3_io_pipe_phv_out_header_0; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_header_1 = proc_3_io_pipe_phv_out_header_1; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_header_2 = proc_3_io_pipe_phv_out_header_2; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_header_3 = proc_3_io_pipe_phv_out_header_3; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_header_4 = proc_3_io_pipe_phv_out_header_4; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_header_5 = proc_3_io_pipe_phv_out_header_5; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_header_6 = proc_3_io_pipe_phv_out_header_6; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_header_7 = proc_3_io_pipe_phv_out_header_7; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_header_8 = proc_3_io_pipe_phv_out_header_8; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_header_9 = proc_3_io_pipe_phv_out_header_9; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_header_10 = proc_3_io_pipe_phv_out_header_10; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_header_11 = proc_3_io_pipe_phv_out_header_11; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_header_12 = proc_3_io_pipe_phv_out_header_12; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_header_13 = proc_3_io_pipe_phv_out_header_13; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_header_14 = proc_3_io_pipe_phv_out_header_14; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_header_15 = proc_3_io_pipe_phv_out_header_15; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_parse_current_state = proc_3_io_pipe_phv_out_parse_current_state; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_parse_current_offset = proc_3_io_pipe_phv_out_parse_current_offset; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_parse_transition_field = proc_3_io_pipe_phv_out_parse_transition_field; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_next_processor_id = proc_3_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 88:32]
  assign trans_3_io_pipe_phv_in_next_config_id = proc_3_io_pipe_phv_out_next_config_id; // @[ipsa.scala 88:32]
  assign trans_3_io_next_proc_exist = last_proc_id != 2'h3; // @[ipsa.scala 86:48]
  assign trans_3_io_next_proc_id_in = next_proc_id_3; // @[ipsa.scala 87:32]
  always @(posedge clock) begin
    if (io_mod_xbar_mod_en) begin // @[ipsa.scala 52:31]
      first_proc_id <= io_mod_xbar_mod_first_proc_id; // @[ipsa.scala 53:23]
    end
    if (io_mod_xbar_mod_en) begin // @[ipsa.scala 52:31]
      last_proc_id <= io_mod_xbar_mod_last_proc_id; // @[ipsa.scala 54:23]
    end
    if (io_mod_xbar_mod_en) begin // @[ipsa.scala 52:31]
      next_proc_id_0 <= io_mod_xbar_mod_next_proc_id_0; // @[ipsa.scala 56:29]
    end
    if (io_mod_xbar_mod_en) begin // @[ipsa.scala 52:31]
      next_proc_id_1 <= io_mod_xbar_mod_next_proc_id_1; // @[ipsa.scala 56:29]
    end
    if (io_mod_xbar_mod_en) begin // @[ipsa.scala 52:31]
      next_proc_id_2 <= io_mod_xbar_mod_next_proc_id_2; // @[ipsa.scala 56:29]
    end
    if (io_mod_xbar_mod_en) begin // @[ipsa.scala 52:31]
      next_proc_id_3 <= io_mod_xbar_mod_next_proc_id_3; // @[ipsa.scala 56:29]
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_0 <= amplifier_1_3_data_0;
    end else begin
      recv_0_data_0 <= amplifier_1_0_data_0;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_1 <= amplifier_1_3_data_1;
    end else begin
      recv_0_data_1 <= amplifier_1_0_data_1;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_2 <= amplifier_1_3_data_2;
    end else begin
      recv_0_data_2 <= amplifier_1_0_data_2;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_3 <= amplifier_1_3_data_3;
    end else begin
      recv_0_data_3 <= amplifier_1_0_data_3;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_4 <= amplifier_1_3_data_4;
    end else begin
      recv_0_data_4 <= amplifier_1_0_data_4;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_5 <= amplifier_1_3_data_5;
    end else begin
      recv_0_data_5 <= amplifier_1_0_data_5;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_6 <= amplifier_1_3_data_6;
    end else begin
      recv_0_data_6 <= amplifier_1_0_data_6;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_7 <= amplifier_1_3_data_7;
    end else begin
      recv_0_data_7 <= amplifier_1_0_data_7;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_8 <= amplifier_1_3_data_8;
    end else begin
      recv_0_data_8 <= amplifier_1_0_data_8;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_9 <= amplifier_1_3_data_9;
    end else begin
      recv_0_data_9 <= amplifier_1_0_data_9;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_10 <= amplifier_1_3_data_10;
    end else begin
      recv_0_data_10 <= amplifier_1_0_data_10;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_11 <= amplifier_1_3_data_11;
    end else begin
      recv_0_data_11 <= amplifier_1_0_data_11;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_12 <= amplifier_1_3_data_12;
    end else begin
      recv_0_data_12 <= amplifier_1_0_data_12;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_13 <= amplifier_1_3_data_13;
    end else begin
      recv_0_data_13 <= amplifier_1_0_data_13;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_14 <= amplifier_1_3_data_14;
    end else begin
      recv_0_data_14 <= amplifier_1_0_data_14;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_15 <= amplifier_1_3_data_15;
    end else begin
      recv_0_data_15 <= amplifier_1_0_data_15;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_16 <= amplifier_1_3_data_16;
    end else begin
      recv_0_data_16 <= amplifier_1_0_data_16;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_17 <= amplifier_1_3_data_17;
    end else begin
      recv_0_data_17 <= amplifier_1_0_data_17;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_18 <= amplifier_1_3_data_18;
    end else begin
      recv_0_data_18 <= amplifier_1_0_data_18;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_19 <= amplifier_1_3_data_19;
    end else begin
      recv_0_data_19 <= amplifier_1_0_data_19;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_20 <= amplifier_1_3_data_20;
    end else begin
      recv_0_data_20 <= amplifier_1_0_data_20;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_21 <= amplifier_1_3_data_21;
    end else begin
      recv_0_data_21 <= amplifier_1_0_data_21;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_22 <= amplifier_1_3_data_22;
    end else begin
      recv_0_data_22 <= amplifier_1_0_data_22;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_23 <= amplifier_1_3_data_23;
    end else begin
      recv_0_data_23 <= amplifier_1_0_data_23;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_24 <= amplifier_1_3_data_24;
    end else begin
      recv_0_data_24 <= amplifier_1_0_data_24;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_25 <= amplifier_1_3_data_25;
    end else begin
      recv_0_data_25 <= amplifier_1_0_data_25;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_26 <= amplifier_1_3_data_26;
    end else begin
      recv_0_data_26 <= amplifier_1_0_data_26;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_27 <= amplifier_1_3_data_27;
    end else begin
      recv_0_data_27 <= amplifier_1_0_data_27;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_28 <= amplifier_1_3_data_28;
    end else begin
      recv_0_data_28 <= amplifier_1_0_data_28;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_29 <= amplifier_1_3_data_29;
    end else begin
      recv_0_data_29 <= amplifier_1_0_data_29;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_30 <= amplifier_1_3_data_30;
    end else begin
      recv_0_data_30 <= amplifier_1_0_data_30;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_31 <= amplifier_1_3_data_31;
    end else begin
      recv_0_data_31 <= amplifier_1_0_data_31;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_32 <= amplifier_1_3_data_32;
    end else begin
      recv_0_data_32 <= amplifier_1_0_data_32;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_33 <= amplifier_1_3_data_33;
    end else begin
      recv_0_data_33 <= amplifier_1_0_data_33;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_34 <= amplifier_1_3_data_34;
    end else begin
      recv_0_data_34 <= amplifier_1_0_data_34;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_35 <= amplifier_1_3_data_35;
    end else begin
      recv_0_data_35 <= amplifier_1_0_data_35;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_36 <= amplifier_1_3_data_36;
    end else begin
      recv_0_data_36 <= amplifier_1_0_data_36;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_37 <= amplifier_1_3_data_37;
    end else begin
      recv_0_data_37 <= amplifier_1_0_data_37;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_38 <= amplifier_1_3_data_38;
    end else begin
      recv_0_data_38 <= amplifier_1_0_data_38;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_39 <= amplifier_1_3_data_39;
    end else begin
      recv_0_data_39 <= amplifier_1_0_data_39;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_40 <= amplifier_1_3_data_40;
    end else begin
      recv_0_data_40 <= amplifier_1_0_data_40;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_41 <= amplifier_1_3_data_41;
    end else begin
      recv_0_data_41 <= amplifier_1_0_data_41;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_42 <= amplifier_1_3_data_42;
    end else begin
      recv_0_data_42 <= amplifier_1_0_data_42;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_43 <= amplifier_1_3_data_43;
    end else begin
      recv_0_data_43 <= amplifier_1_0_data_43;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_44 <= amplifier_1_3_data_44;
    end else begin
      recv_0_data_44 <= amplifier_1_0_data_44;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_45 <= amplifier_1_3_data_45;
    end else begin
      recv_0_data_45 <= amplifier_1_0_data_45;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_46 <= amplifier_1_3_data_46;
    end else begin
      recv_0_data_46 <= amplifier_1_0_data_46;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_47 <= amplifier_1_3_data_47;
    end else begin
      recv_0_data_47 <= amplifier_1_0_data_47;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_48 <= amplifier_1_3_data_48;
    end else begin
      recv_0_data_48 <= amplifier_1_0_data_48;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_49 <= amplifier_1_3_data_49;
    end else begin
      recv_0_data_49 <= amplifier_1_0_data_49;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_50 <= amplifier_1_3_data_50;
    end else begin
      recv_0_data_50 <= amplifier_1_0_data_50;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_51 <= amplifier_1_3_data_51;
    end else begin
      recv_0_data_51 <= amplifier_1_0_data_51;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_52 <= amplifier_1_3_data_52;
    end else begin
      recv_0_data_52 <= amplifier_1_0_data_52;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_53 <= amplifier_1_3_data_53;
    end else begin
      recv_0_data_53 <= amplifier_1_0_data_53;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_54 <= amplifier_1_3_data_54;
    end else begin
      recv_0_data_54 <= amplifier_1_0_data_54;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_55 <= amplifier_1_3_data_55;
    end else begin
      recv_0_data_55 <= amplifier_1_0_data_55;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_56 <= amplifier_1_3_data_56;
    end else begin
      recv_0_data_56 <= amplifier_1_0_data_56;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_57 <= amplifier_1_3_data_57;
    end else begin
      recv_0_data_57 <= amplifier_1_0_data_57;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_58 <= amplifier_1_3_data_58;
    end else begin
      recv_0_data_58 <= amplifier_1_0_data_58;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_59 <= amplifier_1_3_data_59;
    end else begin
      recv_0_data_59 <= amplifier_1_0_data_59;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_60 <= amplifier_1_3_data_60;
    end else begin
      recv_0_data_60 <= amplifier_1_0_data_60;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_61 <= amplifier_1_3_data_61;
    end else begin
      recv_0_data_61 <= amplifier_1_0_data_61;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_62 <= amplifier_1_3_data_62;
    end else begin
      recv_0_data_62 <= amplifier_1_0_data_62;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_63 <= amplifier_1_3_data_63;
    end else begin
      recv_0_data_63 <= amplifier_1_0_data_63;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_64 <= amplifier_1_3_data_64;
    end else begin
      recv_0_data_64 <= amplifier_1_0_data_64;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_65 <= amplifier_1_3_data_65;
    end else begin
      recv_0_data_65 <= amplifier_1_0_data_65;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_66 <= amplifier_1_3_data_66;
    end else begin
      recv_0_data_66 <= amplifier_1_0_data_66;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_67 <= amplifier_1_3_data_67;
    end else begin
      recv_0_data_67 <= amplifier_1_0_data_67;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_68 <= amplifier_1_3_data_68;
    end else begin
      recv_0_data_68 <= amplifier_1_0_data_68;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_69 <= amplifier_1_3_data_69;
    end else begin
      recv_0_data_69 <= amplifier_1_0_data_69;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_70 <= amplifier_1_3_data_70;
    end else begin
      recv_0_data_70 <= amplifier_1_0_data_70;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_71 <= amplifier_1_3_data_71;
    end else begin
      recv_0_data_71 <= amplifier_1_0_data_71;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_72 <= amplifier_1_3_data_72;
    end else begin
      recv_0_data_72 <= amplifier_1_0_data_72;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_73 <= amplifier_1_3_data_73;
    end else begin
      recv_0_data_73 <= amplifier_1_0_data_73;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_74 <= amplifier_1_3_data_74;
    end else begin
      recv_0_data_74 <= amplifier_1_0_data_74;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_75 <= amplifier_1_3_data_75;
    end else begin
      recv_0_data_75 <= amplifier_1_0_data_75;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_76 <= amplifier_1_3_data_76;
    end else begin
      recv_0_data_76 <= amplifier_1_0_data_76;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_77 <= amplifier_1_3_data_77;
    end else begin
      recv_0_data_77 <= amplifier_1_0_data_77;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_78 <= amplifier_1_3_data_78;
    end else begin
      recv_0_data_78 <= amplifier_1_0_data_78;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_79 <= amplifier_1_3_data_79;
    end else begin
      recv_0_data_79 <= amplifier_1_0_data_79;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_80 <= amplifier_1_3_data_80;
    end else begin
      recv_0_data_80 <= amplifier_1_0_data_80;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_81 <= amplifier_1_3_data_81;
    end else begin
      recv_0_data_81 <= amplifier_1_0_data_81;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_82 <= amplifier_1_3_data_82;
    end else begin
      recv_0_data_82 <= amplifier_1_0_data_82;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_83 <= amplifier_1_3_data_83;
    end else begin
      recv_0_data_83 <= amplifier_1_0_data_83;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_84 <= amplifier_1_3_data_84;
    end else begin
      recv_0_data_84 <= amplifier_1_0_data_84;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_85 <= amplifier_1_3_data_85;
    end else begin
      recv_0_data_85 <= amplifier_1_0_data_85;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_86 <= amplifier_1_3_data_86;
    end else begin
      recv_0_data_86 <= amplifier_1_0_data_86;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_87 <= amplifier_1_3_data_87;
    end else begin
      recv_0_data_87 <= amplifier_1_0_data_87;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_88 <= amplifier_1_3_data_88;
    end else begin
      recv_0_data_88 <= amplifier_1_0_data_88;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_89 <= amplifier_1_3_data_89;
    end else begin
      recv_0_data_89 <= amplifier_1_0_data_89;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_90 <= amplifier_1_3_data_90;
    end else begin
      recv_0_data_90 <= amplifier_1_0_data_90;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_91 <= amplifier_1_3_data_91;
    end else begin
      recv_0_data_91 <= amplifier_1_0_data_91;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_92 <= amplifier_1_3_data_92;
    end else begin
      recv_0_data_92 <= amplifier_1_0_data_92;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_93 <= amplifier_1_3_data_93;
    end else begin
      recv_0_data_93 <= amplifier_1_0_data_93;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_94 <= amplifier_1_3_data_94;
    end else begin
      recv_0_data_94 <= amplifier_1_0_data_94;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_95 <= amplifier_1_3_data_95;
    end else begin
      recv_0_data_95 <= amplifier_1_0_data_95;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_96 <= amplifier_1_3_data_96;
    end else begin
      recv_0_data_96 <= amplifier_1_0_data_96;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_97 <= amplifier_1_3_data_97;
    end else begin
      recv_0_data_97 <= amplifier_1_0_data_97;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_98 <= amplifier_1_3_data_98;
    end else begin
      recv_0_data_98 <= amplifier_1_0_data_98;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_99 <= amplifier_1_3_data_99;
    end else begin
      recv_0_data_99 <= amplifier_1_0_data_99;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_100 <= amplifier_1_3_data_100;
    end else begin
      recv_0_data_100 <= amplifier_1_0_data_100;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_101 <= amplifier_1_3_data_101;
    end else begin
      recv_0_data_101 <= amplifier_1_0_data_101;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_102 <= amplifier_1_3_data_102;
    end else begin
      recv_0_data_102 <= amplifier_1_0_data_102;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_103 <= amplifier_1_3_data_103;
    end else begin
      recv_0_data_103 <= amplifier_1_0_data_103;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_104 <= amplifier_1_3_data_104;
    end else begin
      recv_0_data_104 <= amplifier_1_0_data_104;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_105 <= amplifier_1_3_data_105;
    end else begin
      recv_0_data_105 <= amplifier_1_0_data_105;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_106 <= amplifier_1_3_data_106;
    end else begin
      recv_0_data_106 <= amplifier_1_0_data_106;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_107 <= amplifier_1_3_data_107;
    end else begin
      recv_0_data_107 <= amplifier_1_0_data_107;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_108 <= amplifier_1_3_data_108;
    end else begin
      recv_0_data_108 <= amplifier_1_0_data_108;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_109 <= amplifier_1_3_data_109;
    end else begin
      recv_0_data_109 <= amplifier_1_0_data_109;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_110 <= amplifier_1_3_data_110;
    end else begin
      recv_0_data_110 <= amplifier_1_0_data_110;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_111 <= amplifier_1_3_data_111;
    end else begin
      recv_0_data_111 <= amplifier_1_0_data_111;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_112 <= amplifier_1_3_data_112;
    end else begin
      recv_0_data_112 <= amplifier_1_0_data_112;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_113 <= amplifier_1_3_data_113;
    end else begin
      recv_0_data_113 <= amplifier_1_0_data_113;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_114 <= amplifier_1_3_data_114;
    end else begin
      recv_0_data_114 <= amplifier_1_0_data_114;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_115 <= amplifier_1_3_data_115;
    end else begin
      recv_0_data_115 <= amplifier_1_0_data_115;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_116 <= amplifier_1_3_data_116;
    end else begin
      recv_0_data_116 <= amplifier_1_0_data_116;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_117 <= amplifier_1_3_data_117;
    end else begin
      recv_0_data_117 <= amplifier_1_0_data_117;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_118 <= amplifier_1_3_data_118;
    end else begin
      recv_0_data_118 <= amplifier_1_0_data_118;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_119 <= amplifier_1_3_data_119;
    end else begin
      recv_0_data_119 <= amplifier_1_0_data_119;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_120 <= amplifier_1_3_data_120;
    end else begin
      recv_0_data_120 <= amplifier_1_0_data_120;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_121 <= amplifier_1_3_data_121;
    end else begin
      recv_0_data_121 <= amplifier_1_0_data_121;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_122 <= amplifier_1_3_data_122;
    end else begin
      recv_0_data_122 <= amplifier_1_0_data_122;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_123 <= amplifier_1_3_data_123;
    end else begin
      recv_0_data_123 <= amplifier_1_0_data_123;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_124 <= amplifier_1_3_data_124;
    end else begin
      recv_0_data_124 <= amplifier_1_0_data_124;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_125 <= amplifier_1_3_data_125;
    end else begin
      recv_0_data_125 <= amplifier_1_0_data_125;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_126 <= amplifier_1_3_data_126;
    end else begin
      recv_0_data_126 <= amplifier_1_0_data_126;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_127 <= amplifier_1_3_data_127;
    end else begin
      recv_0_data_127 <= amplifier_1_0_data_127;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_128 <= amplifier_1_3_data_128;
    end else begin
      recv_0_data_128 <= amplifier_1_0_data_128;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_129 <= amplifier_1_3_data_129;
    end else begin
      recv_0_data_129 <= amplifier_1_0_data_129;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_130 <= amplifier_1_3_data_130;
    end else begin
      recv_0_data_130 <= amplifier_1_0_data_130;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_131 <= amplifier_1_3_data_131;
    end else begin
      recv_0_data_131 <= amplifier_1_0_data_131;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_132 <= amplifier_1_3_data_132;
    end else begin
      recv_0_data_132 <= amplifier_1_0_data_132;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_133 <= amplifier_1_3_data_133;
    end else begin
      recv_0_data_133 <= amplifier_1_0_data_133;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_134 <= amplifier_1_3_data_134;
    end else begin
      recv_0_data_134 <= amplifier_1_0_data_134;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_135 <= amplifier_1_3_data_135;
    end else begin
      recv_0_data_135 <= amplifier_1_0_data_135;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_136 <= amplifier_1_3_data_136;
    end else begin
      recv_0_data_136 <= amplifier_1_0_data_136;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_137 <= amplifier_1_3_data_137;
    end else begin
      recv_0_data_137 <= amplifier_1_0_data_137;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_138 <= amplifier_1_3_data_138;
    end else begin
      recv_0_data_138 <= amplifier_1_0_data_138;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_139 <= amplifier_1_3_data_139;
    end else begin
      recv_0_data_139 <= amplifier_1_0_data_139;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_140 <= amplifier_1_3_data_140;
    end else begin
      recv_0_data_140 <= amplifier_1_0_data_140;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_141 <= amplifier_1_3_data_141;
    end else begin
      recv_0_data_141 <= amplifier_1_0_data_141;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_142 <= amplifier_1_3_data_142;
    end else begin
      recv_0_data_142 <= amplifier_1_0_data_142;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_143 <= amplifier_1_3_data_143;
    end else begin
      recv_0_data_143 <= amplifier_1_0_data_143;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_144 <= amplifier_1_3_data_144;
    end else begin
      recv_0_data_144 <= amplifier_1_0_data_144;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_145 <= amplifier_1_3_data_145;
    end else begin
      recv_0_data_145 <= amplifier_1_0_data_145;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_146 <= amplifier_1_3_data_146;
    end else begin
      recv_0_data_146 <= amplifier_1_0_data_146;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_147 <= amplifier_1_3_data_147;
    end else begin
      recv_0_data_147 <= amplifier_1_0_data_147;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_148 <= amplifier_1_3_data_148;
    end else begin
      recv_0_data_148 <= amplifier_1_0_data_148;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_149 <= amplifier_1_3_data_149;
    end else begin
      recv_0_data_149 <= amplifier_1_0_data_149;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_150 <= amplifier_1_3_data_150;
    end else begin
      recv_0_data_150 <= amplifier_1_0_data_150;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_151 <= amplifier_1_3_data_151;
    end else begin
      recv_0_data_151 <= amplifier_1_0_data_151;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_152 <= amplifier_1_3_data_152;
    end else begin
      recv_0_data_152 <= amplifier_1_0_data_152;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_153 <= amplifier_1_3_data_153;
    end else begin
      recv_0_data_153 <= amplifier_1_0_data_153;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_154 <= amplifier_1_3_data_154;
    end else begin
      recv_0_data_154 <= amplifier_1_0_data_154;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_155 <= amplifier_1_3_data_155;
    end else begin
      recv_0_data_155 <= amplifier_1_0_data_155;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_156 <= amplifier_1_3_data_156;
    end else begin
      recv_0_data_156 <= amplifier_1_0_data_156;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_157 <= amplifier_1_3_data_157;
    end else begin
      recv_0_data_157 <= amplifier_1_0_data_157;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_158 <= amplifier_1_3_data_158;
    end else begin
      recv_0_data_158 <= amplifier_1_0_data_158;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_159 <= amplifier_1_3_data_159;
    end else begin
      recv_0_data_159 <= amplifier_1_0_data_159;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_160 <= amplifier_1_3_data_160;
    end else begin
      recv_0_data_160 <= amplifier_1_0_data_160;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_161 <= amplifier_1_3_data_161;
    end else begin
      recv_0_data_161 <= amplifier_1_0_data_161;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_162 <= amplifier_1_3_data_162;
    end else begin
      recv_0_data_162 <= amplifier_1_0_data_162;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_163 <= amplifier_1_3_data_163;
    end else begin
      recv_0_data_163 <= amplifier_1_0_data_163;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_164 <= amplifier_1_3_data_164;
    end else begin
      recv_0_data_164 <= amplifier_1_0_data_164;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_165 <= amplifier_1_3_data_165;
    end else begin
      recv_0_data_165 <= amplifier_1_0_data_165;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_166 <= amplifier_1_3_data_166;
    end else begin
      recv_0_data_166 <= amplifier_1_0_data_166;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_167 <= amplifier_1_3_data_167;
    end else begin
      recv_0_data_167 <= amplifier_1_0_data_167;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_168 <= amplifier_1_3_data_168;
    end else begin
      recv_0_data_168 <= amplifier_1_0_data_168;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_169 <= amplifier_1_3_data_169;
    end else begin
      recv_0_data_169 <= amplifier_1_0_data_169;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_170 <= amplifier_1_3_data_170;
    end else begin
      recv_0_data_170 <= amplifier_1_0_data_170;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_171 <= amplifier_1_3_data_171;
    end else begin
      recv_0_data_171 <= amplifier_1_0_data_171;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_172 <= amplifier_1_3_data_172;
    end else begin
      recv_0_data_172 <= amplifier_1_0_data_172;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_173 <= amplifier_1_3_data_173;
    end else begin
      recv_0_data_173 <= amplifier_1_0_data_173;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_174 <= amplifier_1_3_data_174;
    end else begin
      recv_0_data_174 <= amplifier_1_0_data_174;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_175 <= amplifier_1_3_data_175;
    end else begin
      recv_0_data_175 <= amplifier_1_0_data_175;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_176 <= amplifier_1_3_data_176;
    end else begin
      recv_0_data_176 <= amplifier_1_0_data_176;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_177 <= amplifier_1_3_data_177;
    end else begin
      recv_0_data_177 <= amplifier_1_0_data_177;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_178 <= amplifier_1_3_data_178;
    end else begin
      recv_0_data_178 <= amplifier_1_0_data_178;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_179 <= amplifier_1_3_data_179;
    end else begin
      recv_0_data_179 <= amplifier_1_0_data_179;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_180 <= amplifier_1_3_data_180;
    end else begin
      recv_0_data_180 <= amplifier_1_0_data_180;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_181 <= amplifier_1_3_data_181;
    end else begin
      recv_0_data_181 <= amplifier_1_0_data_181;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_182 <= amplifier_1_3_data_182;
    end else begin
      recv_0_data_182 <= amplifier_1_0_data_182;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_183 <= amplifier_1_3_data_183;
    end else begin
      recv_0_data_183 <= amplifier_1_0_data_183;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_184 <= amplifier_1_3_data_184;
    end else begin
      recv_0_data_184 <= amplifier_1_0_data_184;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_185 <= amplifier_1_3_data_185;
    end else begin
      recv_0_data_185 <= amplifier_1_0_data_185;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_186 <= amplifier_1_3_data_186;
    end else begin
      recv_0_data_186 <= amplifier_1_0_data_186;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_187 <= amplifier_1_3_data_187;
    end else begin
      recv_0_data_187 <= amplifier_1_0_data_187;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_188 <= amplifier_1_3_data_188;
    end else begin
      recv_0_data_188 <= amplifier_1_0_data_188;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_189 <= amplifier_1_3_data_189;
    end else begin
      recv_0_data_189 <= amplifier_1_0_data_189;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_190 <= amplifier_1_3_data_190;
    end else begin
      recv_0_data_190 <= amplifier_1_0_data_190;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_191 <= amplifier_1_3_data_191;
    end else begin
      recv_0_data_191 <= amplifier_1_0_data_191;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_192 <= amplifier_1_3_data_192;
    end else begin
      recv_0_data_192 <= amplifier_1_0_data_192;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_193 <= amplifier_1_3_data_193;
    end else begin
      recv_0_data_193 <= amplifier_1_0_data_193;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_194 <= amplifier_1_3_data_194;
    end else begin
      recv_0_data_194 <= amplifier_1_0_data_194;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_195 <= amplifier_1_3_data_195;
    end else begin
      recv_0_data_195 <= amplifier_1_0_data_195;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_196 <= amplifier_1_3_data_196;
    end else begin
      recv_0_data_196 <= amplifier_1_0_data_196;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_197 <= amplifier_1_3_data_197;
    end else begin
      recv_0_data_197 <= amplifier_1_0_data_197;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_198 <= amplifier_1_3_data_198;
    end else begin
      recv_0_data_198 <= amplifier_1_0_data_198;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_199 <= amplifier_1_3_data_199;
    end else begin
      recv_0_data_199 <= amplifier_1_0_data_199;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_200 <= amplifier_1_3_data_200;
    end else begin
      recv_0_data_200 <= amplifier_1_0_data_200;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_201 <= amplifier_1_3_data_201;
    end else begin
      recv_0_data_201 <= amplifier_1_0_data_201;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_202 <= amplifier_1_3_data_202;
    end else begin
      recv_0_data_202 <= amplifier_1_0_data_202;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_203 <= amplifier_1_3_data_203;
    end else begin
      recv_0_data_203 <= amplifier_1_0_data_203;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_204 <= amplifier_1_3_data_204;
    end else begin
      recv_0_data_204 <= amplifier_1_0_data_204;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_205 <= amplifier_1_3_data_205;
    end else begin
      recv_0_data_205 <= amplifier_1_0_data_205;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_206 <= amplifier_1_3_data_206;
    end else begin
      recv_0_data_206 <= amplifier_1_0_data_206;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_207 <= amplifier_1_3_data_207;
    end else begin
      recv_0_data_207 <= amplifier_1_0_data_207;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_208 <= amplifier_1_3_data_208;
    end else begin
      recv_0_data_208 <= amplifier_1_0_data_208;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_209 <= amplifier_1_3_data_209;
    end else begin
      recv_0_data_209 <= amplifier_1_0_data_209;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_210 <= amplifier_1_3_data_210;
    end else begin
      recv_0_data_210 <= amplifier_1_0_data_210;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_211 <= amplifier_1_3_data_211;
    end else begin
      recv_0_data_211 <= amplifier_1_0_data_211;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_212 <= amplifier_1_3_data_212;
    end else begin
      recv_0_data_212 <= amplifier_1_0_data_212;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_213 <= amplifier_1_3_data_213;
    end else begin
      recv_0_data_213 <= amplifier_1_0_data_213;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_214 <= amplifier_1_3_data_214;
    end else begin
      recv_0_data_214 <= amplifier_1_0_data_214;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_215 <= amplifier_1_3_data_215;
    end else begin
      recv_0_data_215 <= amplifier_1_0_data_215;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_216 <= amplifier_1_3_data_216;
    end else begin
      recv_0_data_216 <= amplifier_1_0_data_216;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_217 <= amplifier_1_3_data_217;
    end else begin
      recv_0_data_217 <= amplifier_1_0_data_217;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_218 <= amplifier_1_3_data_218;
    end else begin
      recv_0_data_218 <= amplifier_1_0_data_218;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_219 <= amplifier_1_3_data_219;
    end else begin
      recv_0_data_219 <= amplifier_1_0_data_219;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_220 <= amplifier_1_3_data_220;
    end else begin
      recv_0_data_220 <= amplifier_1_0_data_220;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_221 <= amplifier_1_3_data_221;
    end else begin
      recv_0_data_221 <= amplifier_1_0_data_221;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_222 <= amplifier_1_3_data_222;
    end else begin
      recv_0_data_222 <= amplifier_1_0_data_222;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_223 <= amplifier_1_3_data_223;
    end else begin
      recv_0_data_223 <= amplifier_1_0_data_223;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_224 <= amplifier_1_3_data_224;
    end else begin
      recv_0_data_224 <= amplifier_1_0_data_224;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_225 <= amplifier_1_3_data_225;
    end else begin
      recv_0_data_225 <= amplifier_1_0_data_225;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_226 <= amplifier_1_3_data_226;
    end else begin
      recv_0_data_226 <= amplifier_1_0_data_226;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_227 <= amplifier_1_3_data_227;
    end else begin
      recv_0_data_227 <= amplifier_1_0_data_227;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_228 <= amplifier_1_3_data_228;
    end else begin
      recv_0_data_228 <= amplifier_1_0_data_228;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_229 <= amplifier_1_3_data_229;
    end else begin
      recv_0_data_229 <= amplifier_1_0_data_229;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_230 <= amplifier_1_3_data_230;
    end else begin
      recv_0_data_230 <= amplifier_1_0_data_230;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_231 <= amplifier_1_3_data_231;
    end else begin
      recv_0_data_231 <= amplifier_1_0_data_231;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_232 <= amplifier_1_3_data_232;
    end else begin
      recv_0_data_232 <= amplifier_1_0_data_232;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_233 <= amplifier_1_3_data_233;
    end else begin
      recv_0_data_233 <= amplifier_1_0_data_233;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_234 <= amplifier_1_3_data_234;
    end else begin
      recv_0_data_234 <= amplifier_1_0_data_234;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_235 <= amplifier_1_3_data_235;
    end else begin
      recv_0_data_235 <= amplifier_1_0_data_235;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_236 <= amplifier_1_3_data_236;
    end else begin
      recv_0_data_236 <= amplifier_1_0_data_236;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_237 <= amplifier_1_3_data_237;
    end else begin
      recv_0_data_237 <= amplifier_1_0_data_237;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_238 <= amplifier_1_3_data_238;
    end else begin
      recv_0_data_238 <= amplifier_1_0_data_238;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_239 <= amplifier_1_3_data_239;
    end else begin
      recv_0_data_239 <= amplifier_1_0_data_239;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_240 <= amplifier_1_3_data_240;
    end else begin
      recv_0_data_240 <= amplifier_1_0_data_240;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_241 <= amplifier_1_3_data_241;
    end else begin
      recv_0_data_241 <= amplifier_1_0_data_241;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_242 <= amplifier_1_3_data_242;
    end else begin
      recv_0_data_242 <= amplifier_1_0_data_242;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_243 <= amplifier_1_3_data_243;
    end else begin
      recv_0_data_243 <= amplifier_1_0_data_243;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_244 <= amplifier_1_3_data_244;
    end else begin
      recv_0_data_244 <= amplifier_1_0_data_244;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_245 <= amplifier_1_3_data_245;
    end else begin
      recv_0_data_245 <= amplifier_1_0_data_245;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_246 <= amplifier_1_3_data_246;
    end else begin
      recv_0_data_246 <= amplifier_1_0_data_246;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_247 <= amplifier_1_3_data_247;
    end else begin
      recv_0_data_247 <= amplifier_1_0_data_247;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_248 <= amplifier_1_3_data_248;
    end else begin
      recv_0_data_248 <= amplifier_1_0_data_248;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_249 <= amplifier_1_3_data_249;
    end else begin
      recv_0_data_249 <= amplifier_1_0_data_249;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_250 <= amplifier_1_3_data_250;
    end else begin
      recv_0_data_250 <= amplifier_1_0_data_250;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_251 <= amplifier_1_3_data_251;
    end else begin
      recv_0_data_251 <= amplifier_1_0_data_251;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_252 <= amplifier_1_3_data_252;
    end else begin
      recv_0_data_252 <= amplifier_1_0_data_252;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_253 <= amplifier_1_3_data_253;
    end else begin
      recv_0_data_253 <= amplifier_1_0_data_253;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_254 <= amplifier_1_3_data_254;
    end else begin
      recv_0_data_254 <= amplifier_1_0_data_254;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_data_255 <= amplifier_1_3_data_255;
    end else begin
      recv_0_data_255 <= amplifier_1_0_data_255;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_header_0 <= amplifier_1_3_header_0;
    end else begin
      recv_0_header_0 <= amplifier_1_0_header_0;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_header_1 <= amplifier_1_3_header_1;
    end else begin
      recv_0_header_1 <= amplifier_1_0_header_1;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_header_2 <= amplifier_1_3_header_2;
    end else begin
      recv_0_header_2 <= amplifier_1_0_header_2;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_header_3 <= amplifier_1_3_header_3;
    end else begin
      recv_0_header_3 <= amplifier_1_0_header_3;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_header_4 <= amplifier_1_3_header_4;
    end else begin
      recv_0_header_4 <= amplifier_1_0_header_4;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_header_5 <= amplifier_1_3_header_5;
    end else begin
      recv_0_header_5 <= amplifier_1_0_header_5;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_header_6 <= amplifier_1_3_header_6;
    end else begin
      recv_0_header_6 <= amplifier_1_0_header_6;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_header_7 <= amplifier_1_3_header_7;
    end else begin
      recv_0_header_7 <= amplifier_1_0_header_7;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_header_8 <= amplifier_1_3_header_8;
    end else begin
      recv_0_header_8 <= amplifier_1_0_header_8;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_header_9 <= amplifier_1_3_header_9;
    end else begin
      recv_0_header_9 <= amplifier_1_0_header_9;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_header_10 <= amplifier_1_3_header_10;
    end else begin
      recv_0_header_10 <= amplifier_1_0_header_10;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_header_11 <= amplifier_1_3_header_11;
    end else begin
      recv_0_header_11 <= amplifier_1_0_header_11;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_header_12 <= amplifier_1_3_header_12;
    end else begin
      recv_0_header_12 <= amplifier_1_0_header_12;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_header_13 <= amplifier_1_3_header_13;
    end else begin
      recv_0_header_13 <= amplifier_1_0_header_13;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_header_14 <= amplifier_1_3_header_14;
    end else begin
      recv_0_header_14 <= amplifier_1_0_header_14;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_header_15 <= amplifier_1_3_header_15;
    end else begin
      recv_0_header_15 <= amplifier_1_0_header_15;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_parse_current_state <= amplifier_1_3_parse_current_state;
    end else begin
      recv_0_parse_current_state <= amplifier_1_0_parse_current_state;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_parse_current_offset <= amplifier_1_3_parse_current_offset;
    end else begin
      recv_0_parse_current_offset <= amplifier_1_0_parse_current_offset;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_parse_transition_field <= amplifier_1_3_parse_transition_field;
    end else begin
      recv_0_parse_transition_field <= amplifier_1_0_parse_transition_field;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_next_processor_id <= amplifier_1_3_next_processor_id;
    end else begin
      recv_0_next_processor_id <= amplifier_1_0_next_processor_id;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_next_config_id <= amplifier_1_3_next_config_id;
    end else begin
      recv_0_next_config_id <= amplifier_1_0_next_config_id;
    end
    if (_recv_0_T) begin // @[ipsa.scala 152:23]
      recv_0_is_valid_processor <= amplifier_1_3_is_valid_processor;
    end else begin
      recv_0_is_valid_processor <= amplifier_1_0_is_valid_processor;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_0 <= amplifier_1_2_data_0;
    end else begin
      recv_1_data_0 <= amplifier_1_1_data_0;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_1 <= amplifier_1_2_data_1;
    end else begin
      recv_1_data_1 <= amplifier_1_1_data_1;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_2 <= amplifier_1_2_data_2;
    end else begin
      recv_1_data_2 <= amplifier_1_1_data_2;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_3 <= amplifier_1_2_data_3;
    end else begin
      recv_1_data_3 <= amplifier_1_1_data_3;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_4 <= amplifier_1_2_data_4;
    end else begin
      recv_1_data_4 <= amplifier_1_1_data_4;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_5 <= amplifier_1_2_data_5;
    end else begin
      recv_1_data_5 <= amplifier_1_1_data_5;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_6 <= amplifier_1_2_data_6;
    end else begin
      recv_1_data_6 <= amplifier_1_1_data_6;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_7 <= amplifier_1_2_data_7;
    end else begin
      recv_1_data_7 <= amplifier_1_1_data_7;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_8 <= amplifier_1_2_data_8;
    end else begin
      recv_1_data_8 <= amplifier_1_1_data_8;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_9 <= amplifier_1_2_data_9;
    end else begin
      recv_1_data_9 <= amplifier_1_1_data_9;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_10 <= amplifier_1_2_data_10;
    end else begin
      recv_1_data_10 <= amplifier_1_1_data_10;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_11 <= amplifier_1_2_data_11;
    end else begin
      recv_1_data_11 <= amplifier_1_1_data_11;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_12 <= amplifier_1_2_data_12;
    end else begin
      recv_1_data_12 <= amplifier_1_1_data_12;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_13 <= amplifier_1_2_data_13;
    end else begin
      recv_1_data_13 <= amplifier_1_1_data_13;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_14 <= amplifier_1_2_data_14;
    end else begin
      recv_1_data_14 <= amplifier_1_1_data_14;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_15 <= amplifier_1_2_data_15;
    end else begin
      recv_1_data_15 <= amplifier_1_1_data_15;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_16 <= amplifier_1_2_data_16;
    end else begin
      recv_1_data_16 <= amplifier_1_1_data_16;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_17 <= amplifier_1_2_data_17;
    end else begin
      recv_1_data_17 <= amplifier_1_1_data_17;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_18 <= amplifier_1_2_data_18;
    end else begin
      recv_1_data_18 <= amplifier_1_1_data_18;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_19 <= amplifier_1_2_data_19;
    end else begin
      recv_1_data_19 <= amplifier_1_1_data_19;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_20 <= amplifier_1_2_data_20;
    end else begin
      recv_1_data_20 <= amplifier_1_1_data_20;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_21 <= amplifier_1_2_data_21;
    end else begin
      recv_1_data_21 <= amplifier_1_1_data_21;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_22 <= amplifier_1_2_data_22;
    end else begin
      recv_1_data_22 <= amplifier_1_1_data_22;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_23 <= amplifier_1_2_data_23;
    end else begin
      recv_1_data_23 <= amplifier_1_1_data_23;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_24 <= amplifier_1_2_data_24;
    end else begin
      recv_1_data_24 <= amplifier_1_1_data_24;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_25 <= amplifier_1_2_data_25;
    end else begin
      recv_1_data_25 <= amplifier_1_1_data_25;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_26 <= amplifier_1_2_data_26;
    end else begin
      recv_1_data_26 <= amplifier_1_1_data_26;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_27 <= amplifier_1_2_data_27;
    end else begin
      recv_1_data_27 <= amplifier_1_1_data_27;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_28 <= amplifier_1_2_data_28;
    end else begin
      recv_1_data_28 <= amplifier_1_1_data_28;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_29 <= amplifier_1_2_data_29;
    end else begin
      recv_1_data_29 <= amplifier_1_1_data_29;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_30 <= amplifier_1_2_data_30;
    end else begin
      recv_1_data_30 <= amplifier_1_1_data_30;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_31 <= amplifier_1_2_data_31;
    end else begin
      recv_1_data_31 <= amplifier_1_1_data_31;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_32 <= amplifier_1_2_data_32;
    end else begin
      recv_1_data_32 <= amplifier_1_1_data_32;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_33 <= amplifier_1_2_data_33;
    end else begin
      recv_1_data_33 <= amplifier_1_1_data_33;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_34 <= amplifier_1_2_data_34;
    end else begin
      recv_1_data_34 <= amplifier_1_1_data_34;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_35 <= amplifier_1_2_data_35;
    end else begin
      recv_1_data_35 <= amplifier_1_1_data_35;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_36 <= amplifier_1_2_data_36;
    end else begin
      recv_1_data_36 <= amplifier_1_1_data_36;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_37 <= amplifier_1_2_data_37;
    end else begin
      recv_1_data_37 <= amplifier_1_1_data_37;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_38 <= amplifier_1_2_data_38;
    end else begin
      recv_1_data_38 <= amplifier_1_1_data_38;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_39 <= amplifier_1_2_data_39;
    end else begin
      recv_1_data_39 <= amplifier_1_1_data_39;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_40 <= amplifier_1_2_data_40;
    end else begin
      recv_1_data_40 <= amplifier_1_1_data_40;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_41 <= amplifier_1_2_data_41;
    end else begin
      recv_1_data_41 <= amplifier_1_1_data_41;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_42 <= amplifier_1_2_data_42;
    end else begin
      recv_1_data_42 <= amplifier_1_1_data_42;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_43 <= amplifier_1_2_data_43;
    end else begin
      recv_1_data_43 <= amplifier_1_1_data_43;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_44 <= amplifier_1_2_data_44;
    end else begin
      recv_1_data_44 <= amplifier_1_1_data_44;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_45 <= amplifier_1_2_data_45;
    end else begin
      recv_1_data_45 <= amplifier_1_1_data_45;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_46 <= amplifier_1_2_data_46;
    end else begin
      recv_1_data_46 <= amplifier_1_1_data_46;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_47 <= amplifier_1_2_data_47;
    end else begin
      recv_1_data_47 <= amplifier_1_1_data_47;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_48 <= amplifier_1_2_data_48;
    end else begin
      recv_1_data_48 <= amplifier_1_1_data_48;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_49 <= amplifier_1_2_data_49;
    end else begin
      recv_1_data_49 <= amplifier_1_1_data_49;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_50 <= amplifier_1_2_data_50;
    end else begin
      recv_1_data_50 <= amplifier_1_1_data_50;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_51 <= amplifier_1_2_data_51;
    end else begin
      recv_1_data_51 <= amplifier_1_1_data_51;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_52 <= amplifier_1_2_data_52;
    end else begin
      recv_1_data_52 <= amplifier_1_1_data_52;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_53 <= amplifier_1_2_data_53;
    end else begin
      recv_1_data_53 <= amplifier_1_1_data_53;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_54 <= amplifier_1_2_data_54;
    end else begin
      recv_1_data_54 <= amplifier_1_1_data_54;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_55 <= amplifier_1_2_data_55;
    end else begin
      recv_1_data_55 <= amplifier_1_1_data_55;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_56 <= amplifier_1_2_data_56;
    end else begin
      recv_1_data_56 <= amplifier_1_1_data_56;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_57 <= amplifier_1_2_data_57;
    end else begin
      recv_1_data_57 <= amplifier_1_1_data_57;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_58 <= amplifier_1_2_data_58;
    end else begin
      recv_1_data_58 <= amplifier_1_1_data_58;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_59 <= amplifier_1_2_data_59;
    end else begin
      recv_1_data_59 <= amplifier_1_1_data_59;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_60 <= amplifier_1_2_data_60;
    end else begin
      recv_1_data_60 <= amplifier_1_1_data_60;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_61 <= amplifier_1_2_data_61;
    end else begin
      recv_1_data_61 <= amplifier_1_1_data_61;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_62 <= amplifier_1_2_data_62;
    end else begin
      recv_1_data_62 <= amplifier_1_1_data_62;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_63 <= amplifier_1_2_data_63;
    end else begin
      recv_1_data_63 <= amplifier_1_1_data_63;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_64 <= amplifier_1_2_data_64;
    end else begin
      recv_1_data_64 <= amplifier_1_1_data_64;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_65 <= amplifier_1_2_data_65;
    end else begin
      recv_1_data_65 <= amplifier_1_1_data_65;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_66 <= amplifier_1_2_data_66;
    end else begin
      recv_1_data_66 <= amplifier_1_1_data_66;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_67 <= amplifier_1_2_data_67;
    end else begin
      recv_1_data_67 <= amplifier_1_1_data_67;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_68 <= amplifier_1_2_data_68;
    end else begin
      recv_1_data_68 <= amplifier_1_1_data_68;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_69 <= amplifier_1_2_data_69;
    end else begin
      recv_1_data_69 <= amplifier_1_1_data_69;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_70 <= amplifier_1_2_data_70;
    end else begin
      recv_1_data_70 <= amplifier_1_1_data_70;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_71 <= amplifier_1_2_data_71;
    end else begin
      recv_1_data_71 <= amplifier_1_1_data_71;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_72 <= amplifier_1_2_data_72;
    end else begin
      recv_1_data_72 <= amplifier_1_1_data_72;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_73 <= amplifier_1_2_data_73;
    end else begin
      recv_1_data_73 <= amplifier_1_1_data_73;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_74 <= amplifier_1_2_data_74;
    end else begin
      recv_1_data_74 <= amplifier_1_1_data_74;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_75 <= amplifier_1_2_data_75;
    end else begin
      recv_1_data_75 <= amplifier_1_1_data_75;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_76 <= amplifier_1_2_data_76;
    end else begin
      recv_1_data_76 <= amplifier_1_1_data_76;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_77 <= amplifier_1_2_data_77;
    end else begin
      recv_1_data_77 <= amplifier_1_1_data_77;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_78 <= amplifier_1_2_data_78;
    end else begin
      recv_1_data_78 <= amplifier_1_1_data_78;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_79 <= amplifier_1_2_data_79;
    end else begin
      recv_1_data_79 <= amplifier_1_1_data_79;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_80 <= amplifier_1_2_data_80;
    end else begin
      recv_1_data_80 <= amplifier_1_1_data_80;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_81 <= amplifier_1_2_data_81;
    end else begin
      recv_1_data_81 <= amplifier_1_1_data_81;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_82 <= amplifier_1_2_data_82;
    end else begin
      recv_1_data_82 <= amplifier_1_1_data_82;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_83 <= amplifier_1_2_data_83;
    end else begin
      recv_1_data_83 <= amplifier_1_1_data_83;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_84 <= amplifier_1_2_data_84;
    end else begin
      recv_1_data_84 <= amplifier_1_1_data_84;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_85 <= amplifier_1_2_data_85;
    end else begin
      recv_1_data_85 <= amplifier_1_1_data_85;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_86 <= amplifier_1_2_data_86;
    end else begin
      recv_1_data_86 <= amplifier_1_1_data_86;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_87 <= amplifier_1_2_data_87;
    end else begin
      recv_1_data_87 <= amplifier_1_1_data_87;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_88 <= amplifier_1_2_data_88;
    end else begin
      recv_1_data_88 <= amplifier_1_1_data_88;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_89 <= amplifier_1_2_data_89;
    end else begin
      recv_1_data_89 <= amplifier_1_1_data_89;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_90 <= amplifier_1_2_data_90;
    end else begin
      recv_1_data_90 <= amplifier_1_1_data_90;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_91 <= amplifier_1_2_data_91;
    end else begin
      recv_1_data_91 <= amplifier_1_1_data_91;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_92 <= amplifier_1_2_data_92;
    end else begin
      recv_1_data_92 <= amplifier_1_1_data_92;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_93 <= amplifier_1_2_data_93;
    end else begin
      recv_1_data_93 <= amplifier_1_1_data_93;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_94 <= amplifier_1_2_data_94;
    end else begin
      recv_1_data_94 <= amplifier_1_1_data_94;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_95 <= amplifier_1_2_data_95;
    end else begin
      recv_1_data_95 <= amplifier_1_1_data_95;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_96 <= amplifier_1_2_data_96;
    end else begin
      recv_1_data_96 <= amplifier_1_1_data_96;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_97 <= amplifier_1_2_data_97;
    end else begin
      recv_1_data_97 <= amplifier_1_1_data_97;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_98 <= amplifier_1_2_data_98;
    end else begin
      recv_1_data_98 <= amplifier_1_1_data_98;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_99 <= amplifier_1_2_data_99;
    end else begin
      recv_1_data_99 <= amplifier_1_1_data_99;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_100 <= amplifier_1_2_data_100;
    end else begin
      recv_1_data_100 <= amplifier_1_1_data_100;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_101 <= amplifier_1_2_data_101;
    end else begin
      recv_1_data_101 <= amplifier_1_1_data_101;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_102 <= amplifier_1_2_data_102;
    end else begin
      recv_1_data_102 <= amplifier_1_1_data_102;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_103 <= amplifier_1_2_data_103;
    end else begin
      recv_1_data_103 <= amplifier_1_1_data_103;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_104 <= amplifier_1_2_data_104;
    end else begin
      recv_1_data_104 <= amplifier_1_1_data_104;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_105 <= amplifier_1_2_data_105;
    end else begin
      recv_1_data_105 <= amplifier_1_1_data_105;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_106 <= amplifier_1_2_data_106;
    end else begin
      recv_1_data_106 <= amplifier_1_1_data_106;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_107 <= amplifier_1_2_data_107;
    end else begin
      recv_1_data_107 <= amplifier_1_1_data_107;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_108 <= amplifier_1_2_data_108;
    end else begin
      recv_1_data_108 <= amplifier_1_1_data_108;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_109 <= amplifier_1_2_data_109;
    end else begin
      recv_1_data_109 <= amplifier_1_1_data_109;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_110 <= amplifier_1_2_data_110;
    end else begin
      recv_1_data_110 <= amplifier_1_1_data_110;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_111 <= amplifier_1_2_data_111;
    end else begin
      recv_1_data_111 <= amplifier_1_1_data_111;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_112 <= amplifier_1_2_data_112;
    end else begin
      recv_1_data_112 <= amplifier_1_1_data_112;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_113 <= amplifier_1_2_data_113;
    end else begin
      recv_1_data_113 <= amplifier_1_1_data_113;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_114 <= amplifier_1_2_data_114;
    end else begin
      recv_1_data_114 <= amplifier_1_1_data_114;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_115 <= amplifier_1_2_data_115;
    end else begin
      recv_1_data_115 <= amplifier_1_1_data_115;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_116 <= amplifier_1_2_data_116;
    end else begin
      recv_1_data_116 <= amplifier_1_1_data_116;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_117 <= amplifier_1_2_data_117;
    end else begin
      recv_1_data_117 <= amplifier_1_1_data_117;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_118 <= amplifier_1_2_data_118;
    end else begin
      recv_1_data_118 <= amplifier_1_1_data_118;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_119 <= amplifier_1_2_data_119;
    end else begin
      recv_1_data_119 <= amplifier_1_1_data_119;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_120 <= amplifier_1_2_data_120;
    end else begin
      recv_1_data_120 <= amplifier_1_1_data_120;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_121 <= amplifier_1_2_data_121;
    end else begin
      recv_1_data_121 <= amplifier_1_1_data_121;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_122 <= amplifier_1_2_data_122;
    end else begin
      recv_1_data_122 <= amplifier_1_1_data_122;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_123 <= amplifier_1_2_data_123;
    end else begin
      recv_1_data_123 <= amplifier_1_1_data_123;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_124 <= amplifier_1_2_data_124;
    end else begin
      recv_1_data_124 <= amplifier_1_1_data_124;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_125 <= amplifier_1_2_data_125;
    end else begin
      recv_1_data_125 <= amplifier_1_1_data_125;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_126 <= amplifier_1_2_data_126;
    end else begin
      recv_1_data_126 <= amplifier_1_1_data_126;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_127 <= amplifier_1_2_data_127;
    end else begin
      recv_1_data_127 <= amplifier_1_1_data_127;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_128 <= amplifier_1_2_data_128;
    end else begin
      recv_1_data_128 <= amplifier_1_1_data_128;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_129 <= amplifier_1_2_data_129;
    end else begin
      recv_1_data_129 <= amplifier_1_1_data_129;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_130 <= amplifier_1_2_data_130;
    end else begin
      recv_1_data_130 <= amplifier_1_1_data_130;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_131 <= amplifier_1_2_data_131;
    end else begin
      recv_1_data_131 <= amplifier_1_1_data_131;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_132 <= amplifier_1_2_data_132;
    end else begin
      recv_1_data_132 <= amplifier_1_1_data_132;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_133 <= amplifier_1_2_data_133;
    end else begin
      recv_1_data_133 <= amplifier_1_1_data_133;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_134 <= amplifier_1_2_data_134;
    end else begin
      recv_1_data_134 <= amplifier_1_1_data_134;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_135 <= amplifier_1_2_data_135;
    end else begin
      recv_1_data_135 <= amplifier_1_1_data_135;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_136 <= amplifier_1_2_data_136;
    end else begin
      recv_1_data_136 <= amplifier_1_1_data_136;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_137 <= amplifier_1_2_data_137;
    end else begin
      recv_1_data_137 <= amplifier_1_1_data_137;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_138 <= amplifier_1_2_data_138;
    end else begin
      recv_1_data_138 <= amplifier_1_1_data_138;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_139 <= amplifier_1_2_data_139;
    end else begin
      recv_1_data_139 <= amplifier_1_1_data_139;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_140 <= amplifier_1_2_data_140;
    end else begin
      recv_1_data_140 <= amplifier_1_1_data_140;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_141 <= amplifier_1_2_data_141;
    end else begin
      recv_1_data_141 <= amplifier_1_1_data_141;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_142 <= amplifier_1_2_data_142;
    end else begin
      recv_1_data_142 <= amplifier_1_1_data_142;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_143 <= amplifier_1_2_data_143;
    end else begin
      recv_1_data_143 <= amplifier_1_1_data_143;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_144 <= amplifier_1_2_data_144;
    end else begin
      recv_1_data_144 <= amplifier_1_1_data_144;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_145 <= amplifier_1_2_data_145;
    end else begin
      recv_1_data_145 <= amplifier_1_1_data_145;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_146 <= amplifier_1_2_data_146;
    end else begin
      recv_1_data_146 <= amplifier_1_1_data_146;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_147 <= amplifier_1_2_data_147;
    end else begin
      recv_1_data_147 <= amplifier_1_1_data_147;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_148 <= amplifier_1_2_data_148;
    end else begin
      recv_1_data_148 <= amplifier_1_1_data_148;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_149 <= amplifier_1_2_data_149;
    end else begin
      recv_1_data_149 <= amplifier_1_1_data_149;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_150 <= amplifier_1_2_data_150;
    end else begin
      recv_1_data_150 <= amplifier_1_1_data_150;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_151 <= amplifier_1_2_data_151;
    end else begin
      recv_1_data_151 <= amplifier_1_1_data_151;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_152 <= amplifier_1_2_data_152;
    end else begin
      recv_1_data_152 <= amplifier_1_1_data_152;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_153 <= amplifier_1_2_data_153;
    end else begin
      recv_1_data_153 <= amplifier_1_1_data_153;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_154 <= amplifier_1_2_data_154;
    end else begin
      recv_1_data_154 <= amplifier_1_1_data_154;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_155 <= amplifier_1_2_data_155;
    end else begin
      recv_1_data_155 <= amplifier_1_1_data_155;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_156 <= amplifier_1_2_data_156;
    end else begin
      recv_1_data_156 <= amplifier_1_1_data_156;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_157 <= amplifier_1_2_data_157;
    end else begin
      recv_1_data_157 <= amplifier_1_1_data_157;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_158 <= amplifier_1_2_data_158;
    end else begin
      recv_1_data_158 <= amplifier_1_1_data_158;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_159 <= amplifier_1_2_data_159;
    end else begin
      recv_1_data_159 <= amplifier_1_1_data_159;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_160 <= amplifier_1_2_data_160;
    end else begin
      recv_1_data_160 <= amplifier_1_1_data_160;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_161 <= amplifier_1_2_data_161;
    end else begin
      recv_1_data_161 <= amplifier_1_1_data_161;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_162 <= amplifier_1_2_data_162;
    end else begin
      recv_1_data_162 <= amplifier_1_1_data_162;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_163 <= amplifier_1_2_data_163;
    end else begin
      recv_1_data_163 <= amplifier_1_1_data_163;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_164 <= amplifier_1_2_data_164;
    end else begin
      recv_1_data_164 <= amplifier_1_1_data_164;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_165 <= amplifier_1_2_data_165;
    end else begin
      recv_1_data_165 <= amplifier_1_1_data_165;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_166 <= amplifier_1_2_data_166;
    end else begin
      recv_1_data_166 <= amplifier_1_1_data_166;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_167 <= amplifier_1_2_data_167;
    end else begin
      recv_1_data_167 <= amplifier_1_1_data_167;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_168 <= amplifier_1_2_data_168;
    end else begin
      recv_1_data_168 <= amplifier_1_1_data_168;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_169 <= amplifier_1_2_data_169;
    end else begin
      recv_1_data_169 <= amplifier_1_1_data_169;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_170 <= amplifier_1_2_data_170;
    end else begin
      recv_1_data_170 <= amplifier_1_1_data_170;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_171 <= amplifier_1_2_data_171;
    end else begin
      recv_1_data_171 <= amplifier_1_1_data_171;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_172 <= amplifier_1_2_data_172;
    end else begin
      recv_1_data_172 <= amplifier_1_1_data_172;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_173 <= amplifier_1_2_data_173;
    end else begin
      recv_1_data_173 <= amplifier_1_1_data_173;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_174 <= amplifier_1_2_data_174;
    end else begin
      recv_1_data_174 <= amplifier_1_1_data_174;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_175 <= amplifier_1_2_data_175;
    end else begin
      recv_1_data_175 <= amplifier_1_1_data_175;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_176 <= amplifier_1_2_data_176;
    end else begin
      recv_1_data_176 <= amplifier_1_1_data_176;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_177 <= amplifier_1_2_data_177;
    end else begin
      recv_1_data_177 <= amplifier_1_1_data_177;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_178 <= amplifier_1_2_data_178;
    end else begin
      recv_1_data_178 <= amplifier_1_1_data_178;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_179 <= amplifier_1_2_data_179;
    end else begin
      recv_1_data_179 <= amplifier_1_1_data_179;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_180 <= amplifier_1_2_data_180;
    end else begin
      recv_1_data_180 <= amplifier_1_1_data_180;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_181 <= amplifier_1_2_data_181;
    end else begin
      recv_1_data_181 <= amplifier_1_1_data_181;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_182 <= amplifier_1_2_data_182;
    end else begin
      recv_1_data_182 <= amplifier_1_1_data_182;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_183 <= amplifier_1_2_data_183;
    end else begin
      recv_1_data_183 <= amplifier_1_1_data_183;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_184 <= amplifier_1_2_data_184;
    end else begin
      recv_1_data_184 <= amplifier_1_1_data_184;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_185 <= amplifier_1_2_data_185;
    end else begin
      recv_1_data_185 <= amplifier_1_1_data_185;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_186 <= amplifier_1_2_data_186;
    end else begin
      recv_1_data_186 <= amplifier_1_1_data_186;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_187 <= amplifier_1_2_data_187;
    end else begin
      recv_1_data_187 <= amplifier_1_1_data_187;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_188 <= amplifier_1_2_data_188;
    end else begin
      recv_1_data_188 <= amplifier_1_1_data_188;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_189 <= amplifier_1_2_data_189;
    end else begin
      recv_1_data_189 <= amplifier_1_1_data_189;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_190 <= amplifier_1_2_data_190;
    end else begin
      recv_1_data_190 <= amplifier_1_1_data_190;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_191 <= amplifier_1_2_data_191;
    end else begin
      recv_1_data_191 <= amplifier_1_1_data_191;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_192 <= amplifier_1_2_data_192;
    end else begin
      recv_1_data_192 <= amplifier_1_1_data_192;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_193 <= amplifier_1_2_data_193;
    end else begin
      recv_1_data_193 <= amplifier_1_1_data_193;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_194 <= amplifier_1_2_data_194;
    end else begin
      recv_1_data_194 <= amplifier_1_1_data_194;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_195 <= amplifier_1_2_data_195;
    end else begin
      recv_1_data_195 <= amplifier_1_1_data_195;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_196 <= amplifier_1_2_data_196;
    end else begin
      recv_1_data_196 <= amplifier_1_1_data_196;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_197 <= amplifier_1_2_data_197;
    end else begin
      recv_1_data_197 <= amplifier_1_1_data_197;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_198 <= amplifier_1_2_data_198;
    end else begin
      recv_1_data_198 <= amplifier_1_1_data_198;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_199 <= amplifier_1_2_data_199;
    end else begin
      recv_1_data_199 <= amplifier_1_1_data_199;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_200 <= amplifier_1_2_data_200;
    end else begin
      recv_1_data_200 <= amplifier_1_1_data_200;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_201 <= amplifier_1_2_data_201;
    end else begin
      recv_1_data_201 <= amplifier_1_1_data_201;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_202 <= amplifier_1_2_data_202;
    end else begin
      recv_1_data_202 <= amplifier_1_1_data_202;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_203 <= amplifier_1_2_data_203;
    end else begin
      recv_1_data_203 <= amplifier_1_1_data_203;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_204 <= amplifier_1_2_data_204;
    end else begin
      recv_1_data_204 <= amplifier_1_1_data_204;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_205 <= amplifier_1_2_data_205;
    end else begin
      recv_1_data_205 <= amplifier_1_1_data_205;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_206 <= amplifier_1_2_data_206;
    end else begin
      recv_1_data_206 <= amplifier_1_1_data_206;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_207 <= amplifier_1_2_data_207;
    end else begin
      recv_1_data_207 <= amplifier_1_1_data_207;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_208 <= amplifier_1_2_data_208;
    end else begin
      recv_1_data_208 <= amplifier_1_1_data_208;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_209 <= amplifier_1_2_data_209;
    end else begin
      recv_1_data_209 <= amplifier_1_1_data_209;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_210 <= amplifier_1_2_data_210;
    end else begin
      recv_1_data_210 <= amplifier_1_1_data_210;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_211 <= amplifier_1_2_data_211;
    end else begin
      recv_1_data_211 <= amplifier_1_1_data_211;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_212 <= amplifier_1_2_data_212;
    end else begin
      recv_1_data_212 <= amplifier_1_1_data_212;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_213 <= amplifier_1_2_data_213;
    end else begin
      recv_1_data_213 <= amplifier_1_1_data_213;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_214 <= amplifier_1_2_data_214;
    end else begin
      recv_1_data_214 <= amplifier_1_1_data_214;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_215 <= amplifier_1_2_data_215;
    end else begin
      recv_1_data_215 <= amplifier_1_1_data_215;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_216 <= amplifier_1_2_data_216;
    end else begin
      recv_1_data_216 <= amplifier_1_1_data_216;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_217 <= amplifier_1_2_data_217;
    end else begin
      recv_1_data_217 <= amplifier_1_1_data_217;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_218 <= amplifier_1_2_data_218;
    end else begin
      recv_1_data_218 <= amplifier_1_1_data_218;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_219 <= amplifier_1_2_data_219;
    end else begin
      recv_1_data_219 <= amplifier_1_1_data_219;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_220 <= amplifier_1_2_data_220;
    end else begin
      recv_1_data_220 <= amplifier_1_1_data_220;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_221 <= amplifier_1_2_data_221;
    end else begin
      recv_1_data_221 <= amplifier_1_1_data_221;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_222 <= amplifier_1_2_data_222;
    end else begin
      recv_1_data_222 <= amplifier_1_1_data_222;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_223 <= amplifier_1_2_data_223;
    end else begin
      recv_1_data_223 <= amplifier_1_1_data_223;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_224 <= amplifier_1_2_data_224;
    end else begin
      recv_1_data_224 <= amplifier_1_1_data_224;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_225 <= amplifier_1_2_data_225;
    end else begin
      recv_1_data_225 <= amplifier_1_1_data_225;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_226 <= amplifier_1_2_data_226;
    end else begin
      recv_1_data_226 <= amplifier_1_1_data_226;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_227 <= amplifier_1_2_data_227;
    end else begin
      recv_1_data_227 <= amplifier_1_1_data_227;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_228 <= amplifier_1_2_data_228;
    end else begin
      recv_1_data_228 <= amplifier_1_1_data_228;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_229 <= amplifier_1_2_data_229;
    end else begin
      recv_1_data_229 <= amplifier_1_1_data_229;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_230 <= amplifier_1_2_data_230;
    end else begin
      recv_1_data_230 <= amplifier_1_1_data_230;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_231 <= amplifier_1_2_data_231;
    end else begin
      recv_1_data_231 <= amplifier_1_1_data_231;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_232 <= amplifier_1_2_data_232;
    end else begin
      recv_1_data_232 <= amplifier_1_1_data_232;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_233 <= amplifier_1_2_data_233;
    end else begin
      recv_1_data_233 <= amplifier_1_1_data_233;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_234 <= amplifier_1_2_data_234;
    end else begin
      recv_1_data_234 <= amplifier_1_1_data_234;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_235 <= amplifier_1_2_data_235;
    end else begin
      recv_1_data_235 <= amplifier_1_1_data_235;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_236 <= amplifier_1_2_data_236;
    end else begin
      recv_1_data_236 <= amplifier_1_1_data_236;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_237 <= amplifier_1_2_data_237;
    end else begin
      recv_1_data_237 <= amplifier_1_1_data_237;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_238 <= amplifier_1_2_data_238;
    end else begin
      recv_1_data_238 <= amplifier_1_1_data_238;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_239 <= amplifier_1_2_data_239;
    end else begin
      recv_1_data_239 <= amplifier_1_1_data_239;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_240 <= amplifier_1_2_data_240;
    end else begin
      recv_1_data_240 <= amplifier_1_1_data_240;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_241 <= amplifier_1_2_data_241;
    end else begin
      recv_1_data_241 <= amplifier_1_1_data_241;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_242 <= amplifier_1_2_data_242;
    end else begin
      recv_1_data_242 <= amplifier_1_1_data_242;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_243 <= amplifier_1_2_data_243;
    end else begin
      recv_1_data_243 <= amplifier_1_1_data_243;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_244 <= amplifier_1_2_data_244;
    end else begin
      recv_1_data_244 <= amplifier_1_1_data_244;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_245 <= amplifier_1_2_data_245;
    end else begin
      recv_1_data_245 <= amplifier_1_1_data_245;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_246 <= amplifier_1_2_data_246;
    end else begin
      recv_1_data_246 <= amplifier_1_1_data_246;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_247 <= amplifier_1_2_data_247;
    end else begin
      recv_1_data_247 <= amplifier_1_1_data_247;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_248 <= amplifier_1_2_data_248;
    end else begin
      recv_1_data_248 <= amplifier_1_1_data_248;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_249 <= amplifier_1_2_data_249;
    end else begin
      recv_1_data_249 <= amplifier_1_1_data_249;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_250 <= amplifier_1_2_data_250;
    end else begin
      recv_1_data_250 <= amplifier_1_1_data_250;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_251 <= amplifier_1_2_data_251;
    end else begin
      recv_1_data_251 <= amplifier_1_1_data_251;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_252 <= amplifier_1_2_data_252;
    end else begin
      recv_1_data_252 <= amplifier_1_1_data_252;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_253 <= amplifier_1_2_data_253;
    end else begin
      recv_1_data_253 <= amplifier_1_1_data_253;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_254 <= amplifier_1_2_data_254;
    end else begin
      recv_1_data_254 <= amplifier_1_1_data_254;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_data_255 <= amplifier_1_2_data_255;
    end else begin
      recv_1_data_255 <= amplifier_1_1_data_255;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_header_0 <= amplifier_1_2_header_0;
    end else begin
      recv_1_header_0 <= amplifier_1_1_header_0;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_header_1 <= amplifier_1_2_header_1;
    end else begin
      recv_1_header_1 <= amplifier_1_1_header_1;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_header_2 <= amplifier_1_2_header_2;
    end else begin
      recv_1_header_2 <= amplifier_1_1_header_2;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_header_3 <= amplifier_1_2_header_3;
    end else begin
      recv_1_header_3 <= amplifier_1_1_header_3;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_header_4 <= amplifier_1_2_header_4;
    end else begin
      recv_1_header_4 <= amplifier_1_1_header_4;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_header_5 <= amplifier_1_2_header_5;
    end else begin
      recv_1_header_5 <= amplifier_1_1_header_5;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_header_6 <= amplifier_1_2_header_6;
    end else begin
      recv_1_header_6 <= amplifier_1_1_header_6;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_header_7 <= amplifier_1_2_header_7;
    end else begin
      recv_1_header_7 <= amplifier_1_1_header_7;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_header_8 <= amplifier_1_2_header_8;
    end else begin
      recv_1_header_8 <= amplifier_1_1_header_8;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_header_9 <= amplifier_1_2_header_9;
    end else begin
      recv_1_header_9 <= amplifier_1_1_header_9;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_header_10 <= amplifier_1_2_header_10;
    end else begin
      recv_1_header_10 <= amplifier_1_1_header_10;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_header_11 <= amplifier_1_2_header_11;
    end else begin
      recv_1_header_11 <= amplifier_1_1_header_11;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_header_12 <= amplifier_1_2_header_12;
    end else begin
      recv_1_header_12 <= amplifier_1_1_header_12;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_header_13 <= amplifier_1_2_header_13;
    end else begin
      recv_1_header_13 <= amplifier_1_1_header_13;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_header_14 <= amplifier_1_2_header_14;
    end else begin
      recv_1_header_14 <= amplifier_1_1_header_14;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_header_15 <= amplifier_1_2_header_15;
    end else begin
      recv_1_header_15 <= amplifier_1_1_header_15;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_parse_current_state <= amplifier_1_2_parse_current_state;
    end else begin
      recv_1_parse_current_state <= amplifier_1_1_parse_current_state;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_parse_current_offset <= amplifier_1_2_parse_current_offset;
    end else begin
      recv_1_parse_current_offset <= amplifier_1_1_parse_current_offset;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_parse_transition_field <= amplifier_1_2_parse_transition_field;
    end else begin
      recv_1_parse_transition_field <= amplifier_1_1_parse_transition_field;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_next_processor_id <= amplifier_1_2_next_processor_id;
    end else begin
      recv_1_next_processor_id <= amplifier_1_1_next_processor_id;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_next_config_id <= amplifier_1_2_next_config_id;
    end else begin
      recv_1_next_config_id <= amplifier_1_1_next_config_id;
    end
    if (_recv_1_T) begin // @[ipsa.scala 152:23]
      recv_1_is_valid_processor <= amplifier_1_2_is_valid_processor;
    end else begin
      recv_1_is_valid_processor <= amplifier_1_1_is_valid_processor;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_0 <= amplifier_1_1_data_0;
    end else begin
      recv_2_data_0 <= amplifier_1_2_data_0;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_1 <= amplifier_1_1_data_1;
    end else begin
      recv_2_data_1 <= amplifier_1_2_data_1;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_2 <= amplifier_1_1_data_2;
    end else begin
      recv_2_data_2 <= amplifier_1_2_data_2;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_3 <= amplifier_1_1_data_3;
    end else begin
      recv_2_data_3 <= amplifier_1_2_data_3;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_4 <= amplifier_1_1_data_4;
    end else begin
      recv_2_data_4 <= amplifier_1_2_data_4;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_5 <= amplifier_1_1_data_5;
    end else begin
      recv_2_data_5 <= amplifier_1_2_data_5;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_6 <= amplifier_1_1_data_6;
    end else begin
      recv_2_data_6 <= amplifier_1_2_data_6;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_7 <= amplifier_1_1_data_7;
    end else begin
      recv_2_data_7 <= amplifier_1_2_data_7;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_8 <= amplifier_1_1_data_8;
    end else begin
      recv_2_data_8 <= amplifier_1_2_data_8;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_9 <= amplifier_1_1_data_9;
    end else begin
      recv_2_data_9 <= amplifier_1_2_data_9;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_10 <= amplifier_1_1_data_10;
    end else begin
      recv_2_data_10 <= amplifier_1_2_data_10;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_11 <= amplifier_1_1_data_11;
    end else begin
      recv_2_data_11 <= amplifier_1_2_data_11;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_12 <= amplifier_1_1_data_12;
    end else begin
      recv_2_data_12 <= amplifier_1_2_data_12;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_13 <= amplifier_1_1_data_13;
    end else begin
      recv_2_data_13 <= amplifier_1_2_data_13;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_14 <= amplifier_1_1_data_14;
    end else begin
      recv_2_data_14 <= amplifier_1_2_data_14;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_15 <= amplifier_1_1_data_15;
    end else begin
      recv_2_data_15 <= amplifier_1_2_data_15;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_16 <= amplifier_1_1_data_16;
    end else begin
      recv_2_data_16 <= amplifier_1_2_data_16;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_17 <= amplifier_1_1_data_17;
    end else begin
      recv_2_data_17 <= amplifier_1_2_data_17;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_18 <= amplifier_1_1_data_18;
    end else begin
      recv_2_data_18 <= amplifier_1_2_data_18;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_19 <= amplifier_1_1_data_19;
    end else begin
      recv_2_data_19 <= amplifier_1_2_data_19;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_20 <= amplifier_1_1_data_20;
    end else begin
      recv_2_data_20 <= amplifier_1_2_data_20;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_21 <= amplifier_1_1_data_21;
    end else begin
      recv_2_data_21 <= amplifier_1_2_data_21;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_22 <= amplifier_1_1_data_22;
    end else begin
      recv_2_data_22 <= amplifier_1_2_data_22;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_23 <= amplifier_1_1_data_23;
    end else begin
      recv_2_data_23 <= amplifier_1_2_data_23;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_24 <= amplifier_1_1_data_24;
    end else begin
      recv_2_data_24 <= amplifier_1_2_data_24;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_25 <= amplifier_1_1_data_25;
    end else begin
      recv_2_data_25 <= amplifier_1_2_data_25;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_26 <= amplifier_1_1_data_26;
    end else begin
      recv_2_data_26 <= amplifier_1_2_data_26;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_27 <= amplifier_1_1_data_27;
    end else begin
      recv_2_data_27 <= amplifier_1_2_data_27;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_28 <= amplifier_1_1_data_28;
    end else begin
      recv_2_data_28 <= amplifier_1_2_data_28;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_29 <= amplifier_1_1_data_29;
    end else begin
      recv_2_data_29 <= amplifier_1_2_data_29;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_30 <= amplifier_1_1_data_30;
    end else begin
      recv_2_data_30 <= amplifier_1_2_data_30;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_31 <= amplifier_1_1_data_31;
    end else begin
      recv_2_data_31 <= amplifier_1_2_data_31;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_32 <= amplifier_1_1_data_32;
    end else begin
      recv_2_data_32 <= amplifier_1_2_data_32;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_33 <= amplifier_1_1_data_33;
    end else begin
      recv_2_data_33 <= amplifier_1_2_data_33;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_34 <= amplifier_1_1_data_34;
    end else begin
      recv_2_data_34 <= amplifier_1_2_data_34;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_35 <= amplifier_1_1_data_35;
    end else begin
      recv_2_data_35 <= amplifier_1_2_data_35;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_36 <= amplifier_1_1_data_36;
    end else begin
      recv_2_data_36 <= amplifier_1_2_data_36;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_37 <= amplifier_1_1_data_37;
    end else begin
      recv_2_data_37 <= amplifier_1_2_data_37;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_38 <= amplifier_1_1_data_38;
    end else begin
      recv_2_data_38 <= amplifier_1_2_data_38;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_39 <= amplifier_1_1_data_39;
    end else begin
      recv_2_data_39 <= amplifier_1_2_data_39;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_40 <= amplifier_1_1_data_40;
    end else begin
      recv_2_data_40 <= amplifier_1_2_data_40;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_41 <= amplifier_1_1_data_41;
    end else begin
      recv_2_data_41 <= amplifier_1_2_data_41;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_42 <= amplifier_1_1_data_42;
    end else begin
      recv_2_data_42 <= amplifier_1_2_data_42;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_43 <= amplifier_1_1_data_43;
    end else begin
      recv_2_data_43 <= amplifier_1_2_data_43;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_44 <= amplifier_1_1_data_44;
    end else begin
      recv_2_data_44 <= amplifier_1_2_data_44;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_45 <= amplifier_1_1_data_45;
    end else begin
      recv_2_data_45 <= amplifier_1_2_data_45;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_46 <= amplifier_1_1_data_46;
    end else begin
      recv_2_data_46 <= amplifier_1_2_data_46;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_47 <= amplifier_1_1_data_47;
    end else begin
      recv_2_data_47 <= amplifier_1_2_data_47;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_48 <= amplifier_1_1_data_48;
    end else begin
      recv_2_data_48 <= amplifier_1_2_data_48;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_49 <= amplifier_1_1_data_49;
    end else begin
      recv_2_data_49 <= amplifier_1_2_data_49;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_50 <= amplifier_1_1_data_50;
    end else begin
      recv_2_data_50 <= amplifier_1_2_data_50;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_51 <= amplifier_1_1_data_51;
    end else begin
      recv_2_data_51 <= amplifier_1_2_data_51;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_52 <= amplifier_1_1_data_52;
    end else begin
      recv_2_data_52 <= amplifier_1_2_data_52;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_53 <= amplifier_1_1_data_53;
    end else begin
      recv_2_data_53 <= amplifier_1_2_data_53;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_54 <= amplifier_1_1_data_54;
    end else begin
      recv_2_data_54 <= amplifier_1_2_data_54;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_55 <= amplifier_1_1_data_55;
    end else begin
      recv_2_data_55 <= amplifier_1_2_data_55;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_56 <= amplifier_1_1_data_56;
    end else begin
      recv_2_data_56 <= amplifier_1_2_data_56;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_57 <= amplifier_1_1_data_57;
    end else begin
      recv_2_data_57 <= amplifier_1_2_data_57;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_58 <= amplifier_1_1_data_58;
    end else begin
      recv_2_data_58 <= amplifier_1_2_data_58;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_59 <= amplifier_1_1_data_59;
    end else begin
      recv_2_data_59 <= amplifier_1_2_data_59;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_60 <= amplifier_1_1_data_60;
    end else begin
      recv_2_data_60 <= amplifier_1_2_data_60;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_61 <= amplifier_1_1_data_61;
    end else begin
      recv_2_data_61 <= amplifier_1_2_data_61;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_62 <= amplifier_1_1_data_62;
    end else begin
      recv_2_data_62 <= amplifier_1_2_data_62;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_63 <= amplifier_1_1_data_63;
    end else begin
      recv_2_data_63 <= amplifier_1_2_data_63;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_64 <= amplifier_1_1_data_64;
    end else begin
      recv_2_data_64 <= amplifier_1_2_data_64;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_65 <= amplifier_1_1_data_65;
    end else begin
      recv_2_data_65 <= amplifier_1_2_data_65;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_66 <= amplifier_1_1_data_66;
    end else begin
      recv_2_data_66 <= amplifier_1_2_data_66;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_67 <= amplifier_1_1_data_67;
    end else begin
      recv_2_data_67 <= amplifier_1_2_data_67;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_68 <= amplifier_1_1_data_68;
    end else begin
      recv_2_data_68 <= amplifier_1_2_data_68;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_69 <= amplifier_1_1_data_69;
    end else begin
      recv_2_data_69 <= amplifier_1_2_data_69;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_70 <= amplifier_1_1_data_70;
    end else begin
      recv_2_data_70 <= amplifier_1_2_data_70;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_71 <= amplifier_1_1_data_71;
    end else begin
      recv_2_data_71 <= amplifier_1_2_data_71;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_72 <= amplifier_1_1_data_72;
    end else begin
      recv_2_data_72 <= amplifier_1_2_data_72;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_73 <= amplifier_1_1_data_73;
    end else begin
      recv_2_data_73 <= amplifier_1_2_data_73;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_74 <= amplifier_1_1_data_74;
    end else begin
      recv_2_data_74 <= amplifier_1_2_data_74;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_75 <= amplifier_1_1_data_75;
    end else begin
      recv_2_data_75 <= amplifier_1_2_data_75;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_76 <= amplifier_1_1_data_76;
    end else begin
      recv_2_data_76 <= amplifier_1_2_data_76;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_77 <= amplifier_1_1_data_77;
    end else begin
      recv_2_data_77 <= amplifier_1_2_data_77;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_78 <= amplifier_1_1_data_78;
    end else begin
      recv_2_data_78 <= amplifier_1_2_data_78;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_79 <= amplifier_1_1_data_79;
    end else begin
      recv_2_data_79 <= amplifier_1_2_data_79;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_80 <= amplifier_1_1_data_80;
    end else begin
      recv_2_data_80 <= amplifier_1_2_data_80;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_81 <= amplifier_1_1_data_81;
    end else begin
      recv_2_data_81 <= amplifier_1_2_data_81;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_82 <= amplifier_1_1_data_82;
    end else begin
      recv_2_data_82 <= amplifier_1_2_data_82;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_83 <= amplifier_1_1_data_83;
    end else begin
      recv_2_data_83 <= amplifier_1_2_data_83;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_84 <= amplifier_1_1_data_84;
    end else begin
      recv_2_data_84 <= amplifier_1_2_data_84;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_85 <= amplifier_1_1_data_85;
    end else begin
      recv_2_data_85 <= amplifier_1_2_data_85;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_86 <= amplifier_1_1_data_86;
    end else begin
      recv_2_data_86 <= amplifier_1_2_data_86;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_87 <= amplifier_1_1_data_87;
    end else begin
      recv_2_data_87 <= amplifier_1_2_data_87;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_88 <= amplifier_1_1_data_88;
    end else begin
      recv_2_data_88 <= amplifier_1_2_data_88;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_89 <= amplifier_1_1_data_89;
    end else begin
      recv_2_data_89 <= amplifier_1_2_data_89;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_90 <= amplifier_1_1_data_90;
    end else begin
      recv_2_data_90 <= amplifier_1_2_data_90;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_91 <= amplifier_1_1_data_91;
    end else begin
      recv_2_data_91 <= amplifier_1_2_data_91;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_92 <= amplifier_1_1_data_92;
    end else begin
      recv_2_data_92 <= amplifier_1_2_data_92;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_93 <= amplifier_1_1_data_93;
    end else begin
      recv_2_data_93 <= amplifier_1_2_data_93;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_94 <= amplifier_1_1_data_94;
    end else begin
      recv_2_data_94 <= amplifier_1_2_data_94;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_95 <= amplifier_1_1_data_95;
    end else begin
      recv_2_data_95 <= amplifier_1_2_data_95;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_96 <= amplifier_1_1_data_96;
    end else begin
      recv_2_data_96 <= amplifier_1_2_data_96;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_97 <= amplifier_1_1_data_97;
    end else begin
      recv_2_data_97 <= amplifier_1_2_data_97;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_98 <= amplifier_1_1_data_98;
    end else begin
      recv_2_data_98 <= amplifier_1_2_data_98;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_99 <= amplifier_1_1_data_99;
    end else begin
      recv_2_data_99 <= amplifier_1_2_data_99;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_100 <= amplifier_1_1_data_100;
    end else begin
      recv_2_data_100 <= amplifier_1_2_data_100;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_101 <= amplifier_1_1_data_101;
    end else begin
      recv_2_data_101 <= amplifier_1_2_data_101;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_102 <= amplifier_1_1_data_102;
    end else begin
      recv_2_data_102 <= amplifier_1_2_data_102;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_103 <= amplifier_1_1_data_103;
    end else begin
      recv_2_data_103 <= amplifier_1_2_data_103;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_104 <= amplifier_1_1_data_104;
    end else begin
      recv_2_data_104 <= amplifier_1_2_data_104;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_105 <= amplifier_1_1_data_105;
    end else begin
      recv_2_data_105 <= amplifier_1_2_data_105;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_106 <= amplifier_1_1_data_106;
    end else begin
      recv_2_data_106 <= amplifier_1_2_data_106;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_107 <= amplifier_1_1_data_107;
    end else begin
      recv_2_data_107 <= amplifier_1_2_data_107;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_108 <= amplifier_1_1_data_108;
    end else begin
      recv_2_data_108 <= amplifier_1_2_data_108;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_109 <= amplifier_1_1_data_109;
    end else begin
      recv_2_data_109 <= amplifier_1_2_data_109;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_110 <= amplifier_1_1_data_110;
    end else begin
      recv_2_data_110 <= amplifier_1_2_data_110;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_111 <= amplifier_1_1_data_111;
    end else begin
      recv_2_data_111 <= amplifier_1_2_data_111;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_112 <= amplifier_1_1_data_112;
    end else begin
      recv_2_data_112 <= amplifier_1_2_data_112;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_113 <= amplifier_1_1_data_113;
    end else begin
      recv_2_data_113 <= amplifier_1_2_data_113;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_114 <= amplifier_1_1_data_114;
    end else begin
      recv_2_data_114 <= amplifier_1_2_data_114;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_115 <= amplifier_1_1_data_115;
    end else begin
      recv_2_data_115 <= amplifier_1_2_data_115;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_116 <= amplifier_1_1_data_116;
    end else begin
      recv_2_data_116 <= amplifier_1_2_data_116;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_117 <= amplifier_1_1_data_117;
    end else begin
      recv_2_data_117 <= amplifier_1_2_data_117;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_118 <= amplifier_1_1_data_118;
    end else begin
      recv_2_data_118 <= amplifier_1_2_data_118;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_119 <= amplifier_1_1_data_119;
    end else begin
      recv_2_data_119 <= amplifier_1_2_data_119;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_120 <= amplifier_1_1_data_120;
    end else begin
      recv_2_data_120 <= amplifier_1_2_data_120;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_121 <= amplifier_1_1_data_121;
    end else begin
      recv_2_data_121 <= amplifier_1_2_data_121;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_122 <= amplifier_1_1_data_122;
    end else begin
      recv_2_data_122 <= amplifier_1_2_data_122;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_123 <= amplifier_1_1_data_123;
    end else begin
      recv_2_data_123 <= amplifier_1_2_data_123;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_124 <= amplifier_1_1_data_124;
    end else begin
      recv_2_data_124 <= amplifier_1_2_data_124;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_125 <= amplifier_1_1_data_125;
    end else begin
      recv_2_data_125 <= amplifier_1_2_data_125;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_126 <= amplifier_1_1_data_126;
    end else begin
      recv_2_data_126 <= amplifier_1_2_data_126;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_127 <= amplifier_1_1_data_127;
    end else begin
      recv_2_data_127 <= amplifier_1_2_data_127;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_128 <= amplifier_1_1_data_128;
    end else begin
      recv_2_data_128 <= amplifier_1_2_data_128;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_129 <= amplifier_1_1_data_129;
    end else begin
      recv_2_data_129 <= amplifier_1_2_data_129;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_130 <= amplifier_1_1_data_130;
    end else begin
      recv_2_data_130 <= amplifier_1_2_data_130;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_131 <= amplifier_1_1_data_131;
    end else begin
      recv_2_data_131 <= amplifier_1_2_data_131;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_132 <= amplifier_1_1_data_132;
    end else begin
      recv_2_data_132 <= amplifier_1_2_data_132;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_133 <= amplifier_1_1_data_133;
    end else begin
      recv_2_data_133 <= amplifier_1_2_data_133;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_134 <= amplifier_1_1_data_134;
    end else begin
      recv_2_data_134 <= amplifier_1_2_data_134;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_135 <= amplifier_1_1_data_135;
    end else begin
      recv_2_data_135 <= amplifier_1_2_data_135;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_136 <= amplifier_1_1_data_136;
    end else begin
      recv_2_data_136 <= amplifier_1_2_data_136;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_137 <= amplifier_1_1_data_137;
    end else begin
      recv_2_data_137 <= amplifier_1_2_data_137;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_138 <= amplifier_1_1_data_138;
    end else begin
      recv_2_data_138 <= amplifier_1_2_data_138;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_139 <= amplifier_1_1_data_139;
    end else begin
      recv_2_data_139 <= amplifier_1_2_data_139;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_140 <= amplifier_1_1_data_140;
    end else begin
      recv_2_data_140 <= amplifier_1_2_data_140;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_141 <= amplifier_1_1_data_141;
    end else begin
      recv_2_data_141 <= amplifier_1_2_data_141;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_142 <= amplifier_1_1_data_142;
    end else begin
      recv_2_data_142 <= amplifier_1_2_data_142;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_143 <= amplifier_1_1_data_143;
    end else begin
      recv_2_data_143 <= amplifier_1_2_data_143;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_144 <= amplifier_1_1_data_144;
    end else begin
      recv_2_data_144 <= amplifier_1_2_data_144;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_145 <= amplifier_1_1_data_145;
    end else begin
      recv_2_data_145 <= amplifier_1_2_data_145;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_146 <= amplifier_1_1_data_146;
    end else begin
      recv_2_data_146 <= amplifier_1_2_data_146;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_147 <= amplifier_1_1_data_147;
    end else begin
      recv_2_data_147 <= amplifier_1_2_data_147;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_148 <= amplifier_1_1_data_148;
    end else begin
      recv_2_data_148 <= amplifier_1_2_data_148;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_149 <= amplifier_1_1_data_149;
    end else begin
      recv_2_data_149 <= amplifier_1_2_data_149;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_150 <= amplifier_1_1_data_150;
    end else begin
      recv_2_data_150 <= amplifier_1_2_data_150;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_151 <= amplifier_1_1_data_151;
    end else begin
      recv_2_data_151 <= amplifier_1_2_data_151;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_152 <= amplifier_1_1_data_152;
    end else begin
      recv_2_data_152 <= amplifier_1_2_data_152;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_153 <= amplifier_1_1_data_153;
    end else begin
      recv_2_data_153 <= amplifier_1_2_data_153;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_154 <= amplifier_1_1_data_154;
    end else begin
      recv_2_data_154 <= amplifier_1_2_data_154;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_155 <= amplifier_1_1_data_155;
    end else begin
      recv_2_data_155 <= amplifier_1_2_data_155;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_156 <= amplifier_1_1_data_156;
    end else begin
      recv_2_data_156 <= amplifier_1_2_data_156;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_157 <= amplifier_1_1_data_157;
    end else begin
      recv_2_data_157 <= amplifier_1_2_data_157;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_158 <= amplifier_1_1_data_158;
    end else begin
      recv_2_data_158 <= amplifier_1_2_data_158;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_159 <= amplifier_1_1_data_159;
    end else begin
      recv_2_data_159 <= amplifier_1_2_data_159;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_160 <= amplifier_1_1_data_160;
    end else begin
      recv_2_data_160 <= amplifier_1_2_data_160;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_161 <= amplifier_1_1_data_161;
    end else begin
      recv_2_data_161 <= amplifier_1_2_data_161;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_162 <= amplifier_1_1_data_162;
    end else begin
      recv_2_data_162 <= amplifier_1_2_data_162;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_163 <= amplifier_1_1_data_163;
    end else begin
      recv_2_data_163 <= amplifier_1_2_data_163;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_164 <= amplifier_1_1_data_164;
    end else begin
      recv_2_data_164 <= amplifier_1_2_data_164;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_165 <= amplifier_1_1_data_165;
    end else begin
      recv_2_data_165 <= amplifier_1_2_data_165;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_166 <= amplifier_1_1_data_166;
    end else begin
      recv_2_data_166 <= amplifier_1_2_data_166;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_167 <= amplifier_1_1_data_167;
    end else begin
      recv_2_data_167 <= amplifier_1_2_data_167;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_168 <= amplifier_1_1_data_168;
    end else begin
      recv_2_data_168 <= amplifier_1_2_data_168;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_169 <= amplifier_1_1_data_169;
    end else begin
      recv_2_data_169 <= amplifier_1_2_data_169;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_170 <= amplifier_1_1_data_170;
    end else begin
      recv_2_data_170 <= amplifier_1_2_data_170;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_171 <= amplifier_1_1_data_171;
    end else begin
      recv_2_data_171 <= amplifier_1_2_data_171;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_172 <= amplifier_1_1_data_172;
    end else begin
      recv_2_data_172 <= amplifier_1_2_data_172;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_173 <= amplifier_1_1_data_173;
    end else begin
      recv_2_data_173 <= amplifier_1_2_data_173;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_174 <= amplifier_1_1_data_174;
    end else begin
      recv_2_data_174 <= amplifier_1_2_data_174;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_175 <= amplifier_1_1_data_175;
    end else begin
      recv_2_data_175 <= amplifier_1_2_data_175;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_176 <= amplifier_1_1_data_176;
    end else begin
      recv_2_data_176 <= amplifier_1_2_data_176;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_177 <= amplifier_1_1_data_177;
    end else begin
      recv_2_data_177 <= amplifier_1_2_data_177;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_178 <= amplifier_1_1_data_178;
    end else begin
      recv_2_data_178 <= amplifier_1_2_data_178;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_179 <= amplifier_1_1_data_179;
    end else begin
      recv_2_data_179 <= amplifier_1_2_data_179;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_180 <= amplifier_1_1_data_180;
    end else begin
      recv_2_data_180 <= amplifier_1_2_data_180;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_181 <= amplifier_1_1_data_181;
    end else begin
      recv_2_data_181 <= amplifier_1_2_data_181;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_182 <= amplifier_1_1_data_182;
    end else begin
      recv_2_data_182 <= amplifier_1_2_data_182;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_183 <= amplifier_1_1_data_183;
    end else begin
      recv_2_data_183 <= amplifier_1_2_data_183;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_184 <= amplifier_1_1_data_184;
    end else begin
      recv_2_data_184 <= amplifier_1_2_data_184;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_185 <= amplifier_1_1_data_185;
    end else begin
      recv_2_data_185 <= amplifier_1_2_data_185;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_186 <= amplifier_1_1_data_186;
    end else begin
      recv_2_data_186 <= amplifier_1_2_data_186;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_187 <= amplifier_1_1_data_187;
    end else begin
      recv_2_data_187 <= amplifier_1_2_data_187;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_188 <= amplifier_1_1_data_188;
    end else begin
      recv_2_data_188 <= amplifier_1_2_data_188;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_189 <= amplifier_1_1_data_189;
    end else begin
      recv_2_data_189 <= amplifier_1_2_data_189;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_190 <= amplifier_1_1_data_190;
    end else begin
      recv_2_data_190 <= amplifier_1_2_data_190;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_191 <= amplifier_1_1_data_191;
    end else begin
      recv_2_data_191 <= amplifier_1_2_data_191;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_192 <= amplifier_1_1_data_192;
    end else begin
      recv_2_data_192 <= amplifier_1_2_data_192;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_193 <= amplifier_1_1_data_193;
    end else begin
      recv_2_data_193 <= amplifier_1_2_data_193;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_194 <= amplifier_1_1_data_194;
    end else begin
      recv_2_data_194 <= amplifier_1_2_data_194;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_195 <= amplifier_1_1_data_195;
    end else begin
      recv_2_data_195 <= amplifier_1_2_data_195;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_196 <= amplifier_1_1_data_196;
    end else begin
      recv_2_data_196 <= amplifier_1_2_data_196;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_197 <= amplifier_1_1_data_197;
    end else begin
      recv_2_data_197 <= amplifier_1_2_data_197;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_198 <= amplifier_1_1_data_198;
    end else begin
      recv_2_data_198 <= amplifier_1_2_data_198;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_199 <= amplifier_1_1_data_199;
    end else begin
      recv_2_data_199 <= amplifier_1_2_data_199;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_200 <= amplifier_1_1_data_200;
    end else begin
      recv_2_data_200 <= amplifier_1_2_data_200;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_201 <= amplifier_1_1_data_201;
    end else begin
      recv_2_data_201 <= amplifier_1_2_data_201;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_202 <= amplifier_1_1_data_202;
    end else begin
      recv_2_data_202 <= amplifier_1_2_data_202;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_203 <= amplifier_1_1_data_203;
    end else begin
      recv_2_data_203 <= amplifier_1_2_data_203;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_204 <= amplifier_1_1_data_204;
    end else begin
      recv_2_data_204 <= amplifier_1_2_data_204;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_205 <= amplifier_1_1_data_205;
    end else begin
      recv_2_data_205 <= amplifier_1_2_data_205;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_206 <= amplifier_1_1_data_206;
    end else begin
      recv_2_data_206 <= amplifier_1_2_data_206;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_207 <= amplifier_1_1_data_207;
    end else begin
      recv_2_data_207 <= amplifier_1_2_data_207;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_208 <= amplifier_1_1_data_208;
    end else begin
      recv_2_data_208 <= amplifier_1_2_data_208;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_209 <= amplifier_1_1_data_209;
    end else begin
      recv_2_data_209 <= amplifier_1_2_data_209;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_210 <= amplifier_1_1_data_210;
    end else begin
      recv_2_data_210 <= amplifier_1_2_data_210;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_211 <= amplifier_1_1_data_211;
    end else begin
      recv_2_data_211 <= amplifier_1_2_data_211;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_212 <= amplifier_1_1_data_212;
    end else begin
      recv_2_data_212 <= amplifier_1_2_data_212;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_213 <= amplifier_1_1_data_213;
    end else begin
      recv_2_data_213 <= amplifier_1_2_data_213;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_214 <= amplifier_1_1_data_214;
    end else begin
      recv_2_data_214 <= amplifier_1_2_data_214;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_215 <= amplifier_1_1_data_215;
    end else begin
      recv_2_data_215 <= amplifier_1_2_data_215;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_216 <= amplifier_1_1_data_216;
    end else begin
      recv_2_data_216 <= amplifier_1_2_data_216;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_217 <= amplifier_1_1_data_217;
    end else begin
      recv_2_data_217 <= amplifier_1_2_data_217;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_218 <= amplifier_1_1_data_218;
    end else begin
      recv_2_data_218 <= amplifier_1_2_data_218;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_219 <= amplifier_1_1_data_219;
    end else begin
      recv_2_data_219 <= amplifier_1_2_data_219;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_220 <= amplifier_1_1_data_220;
    end else begin
      recv_2_data_220 <= amplifier_1_2_data_220;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_221 <= amplifier_1_1_data_221;
    end else begin
      recv_2_data_221 <= amplifier_1_2_data_221;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_222 <= amplifier_1_1_data_222;
    end else begin
      recv_2_data_222 <= amplifier_1_2_data_222;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_223 <= amplifier_1_1_data_223;
    end else begin
      recv_2_data_223 <= amplifier_1_2_data_223;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_224 <= amplifier_1_1_data_224;
    end else begin
      recv_2_data_224 <= amplifier_1_2_data_224;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_225 <= amplifier_1_1_data_225;
    end else begin
      recv_2_data_225 <= amplifier_1_2_data_225;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_226 <= amplifier_1_1_data_226;
    end else begin
      recv_2_data_226 <= amplifier_1_2_data_226;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_227 <= amplifier_1_1_data_227;
    end else begin
      recv_2_data_227 <= amplifier_1_2_data_227;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_228 <= amplifier_1_1_data_228;
    end else begin
      recv_2_data_228 <= amplifier_1_2_data_228;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_229 <= amplifier_1_1_data_229;
    end else begin
      recv_2_data_229 <= amplifier_1_2_data_229;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_230 <= amplifier_1_1_data_230;
    end else begin
      recv_2_data_230 <= amplifier_1_2_data_230;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_231 <= amplifier_1_1_data_231;
    end else begin
      recv_2_data_231 <= amplifier_1_2_data_231;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_232 <= amplifier_1_1_data_232;
    end else begin
      recv_2_data_232 <= amplifier_1_2_data_232;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_233 <= amplifier_1_1_data_233;
    end else begin
      recv_2_data_233 <= amplifier_1_2_data_233;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_234 <= amplifier_1_1_data_234;
    end else begin
      recv_2_data_234 <= amplifier_1_2_data_234;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_235 <= amplifier_1_1_data_235;
    end else begin
      recv_2_data_235 <= amplifier_1_2_data_235;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_236 <= amplifier_1_1_data_236;
    end else begin
      recv_2_data_236 <= amplifier_1_2_data_236;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_237 <= amplifier_1_1_data_237;
    end else begin
      recv_2_data_237 <= amplifier_1_2_data_237;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_238 <= amplifier_1_1_data_238;
    end else begin
      recv_2_data_238 <= amplifier_1_2_data_238;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_239 <= amplifier_1_1_data_239;
    end else begin
      recv_2_data_239 <= amplifier_1_2_data_239;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_240 <= amplifier_1_1_data_240;
    end else begin
      recv_2_data_240 <= amplifier_1_2_data_240;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_241 <= amplifier_1_1_data_241;
    end else begin
      recv_2_data_241 <= amplifier_1_2_data_241;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_242 <= amplifier_1_1_data_242;
    end else begin
      recv_2_data_242 <= amplifier_1_2_data_242;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_243 <= amplifier_1_1_data_243;
    end else begin
      recv_2_data_243 <= amplifier_1_2_data_243;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_244 <= amplifier_1_1_data_244;
    end else begin
      recv_2_data_244 <= amplifier_1_2_data_244;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_245 <= amplifier_1_1_data_245;
    end else begin
      recv_2_data_245 <= amplifier_1_2_data_245;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_246 <= amplifier_1_1_data_246;
    end else begin
      recv_2_data_246 <= amplifier_1_2_data_246;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_247 <= amplifier_1_1_data_247;
    end else begin
      recv_2_data_247 <= amplifier_1_2_data_247;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_248 <= amplifier_1_1_data_248;
    end else begin
      recv_2_data_248 <= amplifier_1_2_data_248;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_249 <= amplifier_1_1_data_249;
    end else begin
      recv_2_data_249 <= amplifier_1_2_data_249;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_250 <= amplifier_1_1_data_250;
    end else begin
      recv_2_data_250 <= amplifier_1_2_data_250;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_251 <= amplifier_1_1_data_251;
    end else begin
      recv_2_data_251 <= amplifier_1_2_data_251;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_252 <= amplifier_1_1_data_252;
    end else begin
      recv_2_data_252 <= amplifier_1_2_data_252;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_253 <= amplifier_1_1_data_253;
    end else begin
      recv_2_data_253 <= amplifier_1_2_data_253;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_254 <= amplifier_1_1_data_254;
    end else begin
      recv_2_data_254 <= amplifier_1_2_data_254;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_data_255 <= amplifier_1_1_data_255;
    end else begin
      recv_2_data_255 <= amplifier_1_2_data_255;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_header_0 <= amplifier_1_1_header_0;
    end else begin
      recv_2_header_0 <= amplifier_1_2_header_0;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_header_1 <= amplifier_1_1_header_1;
    end else begin
      recv_2_header_1 <= amplifier_1_2_header_1;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_header_2 <= amplifier_1_1_header_2;
    end else begin
      recv_2_header_2 <= amplifier_1_2_header_2;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_header_3 <= amplifier_1_1_header_3;
    end else begin
      recv_2_header_3 <= amplifier_1_2_header_3;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_header_4 <= amplifier_1_1_header_4;
    end else begin
      recv_2_header_4 <= amplifier_1_2_header_4;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_header_5 <= amplifier_1_1_header_5;
    end else begin
      recv_2_header_5 <= amplifier_1_2_header_5;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_header_6 <= amplifier_1_1_header_6;
    end else begin
      recv_2_header_6 <= amplifier_1_2_header_6;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_header_7 <= amplifier_1_1_header_7;
    end else begin
      recv_2_header_7 <= amplifier_1_2_header_7;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_header_8 <= amplifier_1_1_header_8;
    end else begin
      recv_2_header_8 <= amplifier_1_2_header_8;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_header_9 <= amplifier_1_1_header_9;
    end else begin
      recv_2_header_9 <= amplifier_1_2_header_9;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_header_10 <= amplifier_1_1_header_10;
    end else begin
      recv_2_header_10 <= amplifier_1_2_header_10;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_header_11 <= amplifier_1_1_header_11;
    end else begin
      recv_2_header_11 <= amplifier_1_2_header_11;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_header_12 <= amplifier_1_1_header_12;
    end else begin
      recv_2_header_12 <= amplifier_1_2_header_12;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_header_13 <= amplifier_1_1_header_13;
    end else begin
      recv_2_header_13 <= amplifier_1_2_header_13;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_header_14 <= amplifier_1_1_header_14;
    end else begin
      recv_2_header_14 <= amplifier_1_2_header_14;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_header_15 <= amplifier_1_1_header_15;
    end else begin
      recv_2_header_15 <= amplifier_1_2_header_15;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_parse_current_state <= amplifier_1_1_parse_current_state;
    end else begin
      recv_2_parse_current_state <= amplifier_1_2_parse_current_state;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_parse_current_offset <= amplifier_1_1_parse_current_offset;
    end else begin
      recv_2_parse_current_offset <= amplifier_1_2_parse_current_offset;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_parse_transition_field <= amplifier_1_1_parse_transition_field;
    end else begin
      recv_2_parse_transition_field <= amplifier_1_2_parse_transition_field;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_next_processor_id <= amplifier_1_1_next_processor_id;
    end else begin
      recv_2_next_processor_id <= amplifier_1_2_next_processor_id;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_next_config_id <= amplifier_1_1_next_config_id;
    end else begin
      recv_2_next_config_id <= amplifier_1_2_next_config_id;
    end
    if (_recv_2_T) begin // @[ipsa.scala 155:23]
      recv_2_is_valid_processor <= amplifier_1_1_is_valid_processor;
    end else begin
      recv_2_is_valid_processor <= amplifier_1_2_is_valid_processor;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_0 <= amplifier_1_0_data_0;
    end else begin
      recv_3_data_0 <= amplifier_1_3_data_0;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_1 <= amplifier_1_0_data_1;
    end else begin
      recv_3_data_1 <= amplifier_1_3_data_1;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_2 <= amplifier_1_0_data_2;
    end else begin
      recv_3_data_2 <= amplifier_1_3_data_2;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_3 <= amplifier_1_0_data_3;
    end else begin
      recv_3_data_3 <= amplifier_1_3_data_3;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_4 <= amplifier_1_0_data_4;
    end else begin
      recv_3_data_4 <= amplifier_1_3_data_4;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_5 <= amplifier_1_0_data_5;
    end else begin
      recv_3_data_5 <= amplifier_1_3_data_5;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_6 <= amplifier_1_0_data_6;
    end else begin
      recv_3_data_6 <= amplifier_1_3_data_6;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_7 <= amplifier_1_0_data_7;
    end else begin
      recv_3_data_7 <= amplifier_1_3_data_7;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_8 <= amplifier_1_0_data_8;
    end else begin
      recv_3_data_8 <= amplifier_1_3_data_8;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_9 <= amplifier_1_0_data_9;
    end else begin
      recv_3_data_9 <= amplifier_1_3_data_9;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_10 <= amplifier_1_0_data_10;
    end else begin
      recv_3_data_10 <= amplifier_1_3_data_10;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_11 <= amplifier_1_0_data_11;
    end else begin
      recv_3_data_11 <= amplifier_1_3_data_11;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_12 <= amplifier_1_0_data_12;
    end else begin
      recv_3_data_12 <= amplifier_1_3_data_12;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_13 <= amplifier_1_0_data_13;
    end else begin
      recv_3_data_13 <= amplifier_1_3_data_13;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_14 <= amplifier_1_0_data_14;
    end else begin
      recv_3_data_14 <= amplifier_1_3_data_14;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_15 <= amplifier_1_0_data_15;
    end else begin
      recv_3_data_15 <= amplifier_1_3_data_15;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_16 <= amplifier_1_0_data_16;
    end else begin
      recv_3_data_16 <= amplifier_1_3_data_16;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_17 <= amplifier_1_0_data_17;
    end else begin
      recv_3_data_17 <= amplifier_1_3_data_17;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_18 <= amplifier_1_0_data_18;
    end else begin
      recv_3_data_18 <= amplifier_1_3_data_18;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_19 <= amplifier_1_0_data_19;
    end else begin
      recv_3_data_19 <= amplifier_1_3_data_19;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_20 <= amplifier_1_0_data_20;
    end else begin
      recv_3_data_20 <= amplifier_1_3_data_20;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_21 <= amplifier_1_0_data_21;
    end else begin
      recv_3_data_21 <= amplifier_1_3_data_21;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_22 <= amplifier_1_0_data_22;
    end else begin
      recv_3_data_22 <= amplifier_1_3_data_22;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_23 <= amplifier_1_0_data_23;
    end else begin
      recv_3_data_23 <= amplifier_1_3_data_23;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_24 <= amplifier_1_0_data_24;
    end else begin
      recv_3_data_24 <= amplifier_1_3_data_24;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_25 <= amplifier_1_0_data_25;
    end else begin
      recv_3_data_25 <= amplifier_1_3_data_25;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_26 <= amplifier_1_0_data_26;
    end else begin
      recv_3_data_26 <= amplifier_1_3_data_26;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_27 <= amplifier_1_0_data_27;
    end else begin
      recv_3_data_27 <= amplifier_1_3_data_27;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_28 <= amplifier_1_0_data_28;
    end else begin
      recv_3_data_28 <= amplifier_1_3_data_28;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_29 <= amplifier_1_0_data_29;
    end else begin
      recv_3_data_29 <= amplifier_1_3_data_29;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_30 <= amplifier_1_0_data_30;
    end else begin
      recv_3_data_30 <= amplifier_1_3_data_30;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_31 <= amplifier_1_0_data_31;
    end else begin
      recv_3_data_31 <= amplifier_1_3_data_31;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_32 <= amplifier_1_0_data_32;
    end else begin
      recv_3_data_32 <= amplifier_1_3_data_32;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_33 <= amplifier_1_0_data_33;
    end else begin
      recv_3_data_33 <= amplifier_1_3_data_33;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_34 <= amplifier_1_0_data_34;
    end else begin
      recv_3_data_34 <= amplifier_1_3_data_34;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_35 <= amplifier_1_0_data_35;
    end else begin
      recv_3_data_35 <= amplifier_1_3_data_35;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_36 <= amplifier_1_0_data_36;
    end else begin
      recv_3_data_36 <= amplifier_1_3_data_36;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_37 <= amplifier_1_0_data_37;
    end else begin
      recv_3_data_37 <= amplifier_1_3_data_37;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_38 <= amplifier_1_0_data_38;
    end else begin
      recv_3_data_38 <= amplifier_1_3_data_38;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_39 <= amplifier_1_0_data_39;
    end else begin
      recv_3_data_39 <= amplifier_1_3_data_39;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_40 <= amplifier_1_0_data_40;
    end else begin
      recv_3_data_40 <= amplifier_1_3_data_40;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_41 <= amplifier_1_0_data_41;
    end else begin
      recv_3_data_41 <= amplifier_1_3_data_41;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_42 <= amplifier_1_0_data_42;
    end else begin
      recv_3_data_42 <= amplifier_1_3_data_42;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_43 <= amplifier_1_0_data_43;
    end else begin
      recv_3_data_43 <= amplifier_1_3_data_43;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_44 <= amplifier_1_0_data_44;
    end else begin
      recv_3_data_44 <= amplifier_1_3_data_44;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_45 <= amplifier_1_0_data_45;
    end else begin
      recv_3_data_45 <= amplifier_1_3_data_45;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_46 <= amplifier_1_0_data_46;
    end else begin
      recv_3_data_46 <= amplifier_1_3_data_46;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_47 <= amplifier_1_0_data_47;
    end else begin
      recv_3_data_47 <= amplifier_1_3_data_47;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_48 <= amplifier_1_0_data_48;
    end else begin
      recv_3_data_48 <= amplifier_1_3_data_48;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_49 <= amplifier_1_0_data_49;
    end else begin
      recv_3_data_49 <= amplifier_1_3_data_49;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_50 <= amplifier_1_0_data_50;
    end else begin
      recv_3_data_50 <= amplifier_1_3_data_50;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_51 <= amplifier_1_0_data_51;
    end else begin
      recv_3_data_51 <= amplifier_1_3_data_51;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_52 <= amplifier_1_0_data_52;
    end else begin
      recv_3_data_52 <= amplifier_1_3_data_52;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_53 <= amplifier_1_0_data_53;
    end else begin
      recv_3_data_53 <= amplifier_1_3_data_53;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_54 <= amplifier_1_0_data_54;
    end else begin
      recv_3_data_54 <= amplifier_1_3_data_54;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_55 <= amplifier_1_0_data_55;
    end else begin
      recv_3_data_55 <= amplifier_1_3_data_55;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_56 <= amplifier_1_0_data_56;
    end else begin
      recv_3_data_56 <= amplifier_1_3_data_56;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_57 <= amplifier_1_0_data_57;
    end else begin
      recv_3_data_57 <= amplifier_1_3_data_57;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_58 <= amplifier_1_0_data_58;
    end else begin
      recv_3_data_58 <= amplifier_1_3_data_58;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_59 <= amplifier_1_0_data_59;
    end else begin
      recv_3_data_59 <= amplifier_1_3_data_59;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_60 <= amplifier_1_0_data_60;
    end else begin
      recv_3_data_60 <= amplifier_1_3_data_60;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_61 <= amplifier_1_0_data_61;
    end else begin
      recv_3_data_61 <= amplifier_1_3_data_61;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_62 <= amplifier_1_0_data_62;
    end else begin
      recv_3_data_62 <= amplifier_1_3_data_62;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_63 <= amplifier_1_0_data_63;
    end else begin
      recv_3_data_63 <= amplifier_1_3_data_63;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_64 <= amplifier_1_0_data_64;
    end else begin
      recv_3_data_64 <= amplifier_1_3_data_64;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_65 <= amplifier_1_0_data_65;
    end else begin
      recv_3_data_65 <= amplifier_1_3_data_65;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_66 <= amplifier_1_0_data_66;
    end else begin
      recv_3_data_66 <= amplifier_1_3_data_66;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_67 <= amplifier_1_0_data_67;
    end else begin
      recv_3_data_67 <= amplifier_1_3_data_67;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_68 <= amplifier_1_0_data_68;
    end else begin
      recv_3_data_68 <= amplifier_1_3_data_68;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_69 <= amplifier_1_0_data_69;
    end else begin
      recv_3_data_69 <= amplifier_1_3_data_69;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_70 <= amplifier_1_0_data_70;
    end else begin
      recv_3_data_70 <= amplifier_1_3_data_70;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_71 <= amplifier_1_0_data_71;
    end else begin
      recv_3_data_71 <= amplifier_1_3_data_71;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_72 <= amplifier_1_0_data_72;
    end else begin
      recv_3_data_72 <= amplifier_1_3_data_72;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_73 <= amplifier_1_0_data_73;
    end else begin
      recv_3_data_73 <= amplifier_1_3_data_73;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_74 <= amplifier_1_0_data_74;
    end else begin
      recv_3_data_74 <= amplifier_1_3_data_74;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_75 <= amplifier_1_0_data_75;
    end else begin
      recv_3_data_75 <= amplifier_1_3_data_75;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_76 <= amplifier_1_0_data_76;
    end else begin
      recv_3_data_76 <= amplifier_1_3_data_76;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_77 <= amplifier_1_0_data_77;
    end else begin
      recv_3_data_77 <= amplifier_1_3_data_77;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_78 <= amplifier_1_0_data_78;
    end else begin
      recv_3_data_78 <= amplifier_1_3_data_78;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_79 <= amplifier_1_0_data_79;
    end else begin
      recv_3_data_79 <= amplifier_1_3_data_79;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_80 <= amplifier_1_0_data_80;
    end else begin
      recv_3_data_80 <= amplifier_1_3_data_80;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_81 <= amplifier_1_0_data_81;
    end else begin
      recv_3_data_81 <= amplifier_1_3_data_81;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_82 <= amplifier_1_0_data_82;
    end else begin
      recv_3_data_82 <= amplifier_1_3_data_82;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_83 <= amplifier_1_0_data_83;
    end else begin
      recv_3_data_83 <= amplifier_1_3_data_83;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_84 <= amplifier_1_0_data_84;
    end else begin
      recv_3_data_84 <= amplifier_1_3_data_84;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_85 <= amplifier_1_0_data_85;
    end else begin
      recv_3_data_85 <= amplifier_1_3_data_85;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_86 <= amplifier_1_0_data_86;
    end else begin
      recv_3_data_86 <= amplifier_1_3_data_86;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_87 <= amplifier_1_0_data_87;
    end else begin
      recv_3_data_87 <= amplifier_1_3_data_87;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_88 <= amplifier_1_0_data_88;
    end else begin
      recv_3_data_88 <= amplifier_1_3_data_88;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_89 <= amplifier_1_0_data_89;
    end else begin
      recv_3_data_89 <= amplifier_1_3_data_89;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_90 <= amplifier_1_0_data_90;
    end else begin
      recv_3_data_90 <= amplifier_1_3_data_90;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_91 <= amplifier_1_0_data_91;
    end else begin
      recv_3_data_91 <= amplifier_1_3_data_91;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_92 <= amplifier_1_0_data_92;
    end else begin
      recv_3_data_92 <= amplifier_1_3_data_92;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_93 <= amplifier_1_0_data_93;
    end else begin
      recv_3_data_93 <= amplifier_1_3_data_93;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_94 <= amplifier_1_0_data_94;
    end else begin
      recv_3_data_94 <= amplifier_1_3_data_94;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_95 <= amplifier_1_0_data_95;
    end else begin
      recv_3_data_95 <= amplifier_1_3_data_95;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_96 <= amplifier_1_0_data_96;
    end else begin
      recv_3_data_96 <= amplifier_1_3_data_96;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_97 <= amplifier_1_0_data_97;
    end else begin
      recv_3_data_97 <= amplifier_1_3_data_97;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_98 <= amplifier_1_0_data_98;
    end else begin
      recv_3_data_98 <= amplifier_1_3_data_98;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_99 <= amplifier_1_0_data_99;
    end else begin
      recv_3_data_99 <= amplifier_1_3_data_99;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_100 <= amplifier_1_0_data_100;
    end else begin
      recv_3_data_100 <= amplifier_1_3_data_100;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_101 <= amplifier_1_0_data_101;
    end else begin
      recv_3_data_101 <= amplifier_1_3_data_101;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_102 <= amplifier_1_0_data_102;
    end else begin
      recv_3_data_102 <= amplifier_1_3_data_102;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_103 <= amplifier_1_0_data_103;
    end else begin
      recv_3_data_103 <= amplifier_1_3_data_103;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_104 <= amplifier_1_0_data_104;
    end else begin
      recv_3_data_104 <= amplifier_1_3_data_104;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_105 <= amplifier_1_0_data_105;
    end else begin
      recv_3_data_105 <= amplifier_1_3_data_105;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_106 <= amplifier_1_0_data_106;
    end else begin
      recv_3_data_106 <= amplifier_1_3_data_106;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_107 <= amplifier_1_0_data_107;
    end else begin
      recv_3_data_107 <= amplifier_1_3_data_107;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_108 <= amplifier_1_0_data_108;
    end else begin
      recv_3_data_108 <= amplifier_1_3_data_108;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_109 <= amplifier_1_0_data_109;
    end else begin
      recv_3_data_109 <= amplifier_1_3_data_109;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_110 <= amplifier_1_0_data_110;
    end else begin
      recv_3_data_110 <= amplifier_1_3_data_110;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_111 <= amplifier_1_0_data_111;
    end else begin
      recv_3_data_111 <= amplifier_1_3_data_111;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_112 <= amplifier_1_0_data_112;
    end else begin
      recv_3_data_112 <= amplifier_1_3_data_112;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_113 <= amplifier_1_0_data_113;
    end else begin
      recv_3_data_113 <= amplifier_1_3_data_113;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_114 <= amplifier_1_0_data_114;
    end else begin
      recv_3_data_114 <= amplifier_1_3_data_114;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_115 <= amplifier_1_0_data_115;
    end else begin
      recv_3_data_115 <= amplifier_1_3_data_115;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_116 <= amplifier_1_0_data_116;
    end else begin
      recv_3_data_116 <= amplifier_1_3_data_116;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_117 <= amplifier_1_0_data_117;
    end else begin
      recv_3_data_117 <= amplifier_1_3_data_117;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_118 <= amplifier_1_0_data_118;
    end else begin
      recv_3_data_118 <= amplifier_1_3_data_118;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_119 <= amplifier_1_0_data_119;
    end else begin
      recv_3_data_119 <= amplifier_1_3_data_119;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_120 <= amplifier_1_0_data_120;
    end else begin
      recv_3_data_120 <= amplifier_1_3_data_120;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_121 <= amplifier_1_0_data_121;
    end else begin
      recv_3_data_121 <= amplifier_1_3_data_121;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_122 <= amplifier_1_0_data_122;
    end else begin
      recv_3_data_122 <= amplifier_1_3_data_122;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_123 <= amplifier_1_0_data_123;
    end else begin
      recv_3_data_123 <= amplifier_1_3_data_123;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_124 <= amplifier_1_0_data_124;
    end else begin
      recv_3_data_124 <= amplifier_1_3_data_124;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_125 <= amplifier_1_0_data_125;
    end else begin
      recv_3_data_125 <= amplifier_1_3_data_125;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_126 <= amplifier_1_0_data_126;
    end else begin
      recv_3_data_126 <= amplifier_1_3_data_126;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_127 <= amplifier_1_0_data_127;
    end else begin
      recv_3_data_127 <= amplifier_1_3_data_127;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_128 <= amplifier_1_0_data_128;
    end else begin
      recv_3_data_128 <= amplifier_1_3_data_128;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_129 <= amplifier_1_0_data_129;
    end else begin
      recv_3_data_129 <= amplifier_1_3_data_129;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_130 <= amplifier_1_0_data_130;
    end else begin
      recv_3_data_130 <= amplifier_1_3_data_130;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_131 <= amplifier_1_0_data_131;
    end else begin
      recv_3_data_131 <= amplifier_1_3_data_131;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_132 <= amplifier_1_0_data_132;
    end else begin
      recv_3_data_132 <= amplifier_1_3_data_132;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_133 <= amplifier_1_0_data_133;
    end else begin
      recv_3_data_133 <= amplifier_1_3_data_133;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_134 <= amplifier_1_0_data_134;
    end else begin
      recv_3_data_134 <= amplifier_1_3_data_134;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_135 <= amplifier_1_0_data_135;
    end else begin
      recv_3_data_135 <= amplifier_1_3_data_135;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_136 <= amplifier_1_0_data_136;
    end else begin
      recv_3_data_136 <= amplifier_1_3_data_136;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_137 <= amplifier_1_0_data_137;
    end else begin
      recv_3_data_137 <= amplifier_1_3_data_137;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_138 <= amplifier_1_0_data_138;
    end else begin
      recv_3_data_138 <= amplifier_1_3_data_138;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_139 <= amplifier_1_0_data_139;
    end else begin
      recv_3_data_139 <= amplifier_1_3_data_139;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_140 <= amplifier_1_0_data_140;
    end else begin
      recv_3_data_140 <= amplifier_1_3_data_140;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_141 <= amplifier_1_0_data_141;
    end else begin
      recv_3_data_141 <= amplifier_1_3_data_141;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_142 <= amplifier_1_0_data_142;
    end else begin
      recv_3_data_142 <= amplifier_1_3_data_142;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_143 <= amplifier_1_0_data_143;
    end else begin
      recv_3_data_143 <= amplifier_1_3_data_143;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_144 <= amplifier_1_0_data_144;
    end else begin
      recv_3_data_144 <= amplifier_1_3_data_144;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_145 <= amplifier_1_0_data_145;
    end else begin
      recv_3_data_145 <= amplifier_1_3_data_145;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_146 <= amplifier_1_0_data_146;
    end else begin
      recv_3_data_146 <= amplifier_1_3_data_146;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_147 <= amplifier_1_0_data_147;
    end else begin
      recv_3_data_147 <= amplifier_1_3_data_147;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_148 <= amplifier_1_0_data_148;
    end else begin
      recv_3_data_148 <= amplifier_1_3_data_148;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_149 <= amplifier_1_0_data_149;
    end else begin
      recv_3_data_149 <= amplifier_1_3_data_149;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_150 <= amplifier_1_0_data_150;
    end else begin
      recv_3_data_150 <= amplifier_1_3_data_150;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_151 <= amplifier_1_0_data_151;
    end else begin
      recv_3_data_151 <= amplifier_1_3_data_151;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_152 <= amplifier_1_0_data_152;
    end else begin
      recv_3_data_152 <= amplifier_1_3_data_152;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_153 <= amplifier_1_0_data_153;
    end else begin
      recv_3_data_153 <= amplifier_1_3_data_153;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_154 <= amplifier_1_0_data_154;
    end else begin
      recv_3_data_154 <= amplifier_1_3_data_154;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_155 <= amplifier_1_0_data_155;
    end else begin
      recv_3_data_155 <= amplifier_1_3_data_155;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_156 <= amplifier_1_0_data_156;
    end else begin
      recv_3_data_156 <= amplifier_1_3_data_156;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_157 <= amplifier_1_0_data_157;
    end else begin
      recv_3_data_157 <= amplifier_1_3_data_157;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_158 <= amplifier_1_0_data_158;
    end else begin
      recv_3_data_158 <= amplifier_1_3_data_158;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_159 <= amplifier_1_0_data_159;
    end else begin
      recv_3_data_159 <= amplifier_1_3_data_159;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_160 <= amplifier_1_0_data_160;
    end else begin
      recv_3_data_160 <= amplifier_1_3_data_160;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_161 <= amplifier_1_0_data_161;
    end else begin
      recv_3_data_161 <= amplifier_1_3_data_161;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_162 <= amplifier_1_0_data_162;
    end else begin
      recv_3_data_162 <= amplifier_1_3_data_162;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_163 <= amplifier_1_0_data_163;
    end else begin
      recv_3_data_163 <= amplifier_1_3_data_163;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_164 <= amplifier_1_0_data_164;
    end else begin
      recv_3_data_164 <= amplifier_1_3_data_164;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_165 <= amplifier_1_0_data_165;
    end else begin
      recv_3_data_165 <= amplifier_1_3_data_165;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_166 <= amplifier_1_0_data_166;
    end else begin
      recv_3_data_166 <= amplifier_1_3_data_166;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_167 <= amplifier_1_0_data_167;
    end else begin
      recv_3_data_167 <= amplifier_1_3_data_167;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_168 <= amplifier_1_0_data_168;
    end else begin
      recv_3_data_168 <= amplifier_1_3_data_168;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_169 <= amplifier_1_0_data_169;
    end else begin
      recv_3_data_169 <= amplifier_1_3_data_169;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_170 <= amplifier_1_0_data_170;
    end else begin
      recv_3_data_170 <= amplifier_1_3_data_170;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_171 <= amplifier_1_0_data_171;
    end else begin
      recv_3_data_171 <= amplifier_1_3_data_171;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_172 <= amplifier_1_0_data_172;
    end else begin
      recv_3_data_172 <= amplifier_1_3_data_172;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_173 <= amplifier_1_0_data_173;
    end else begin
      recv_3_data_173 <= amplifier_1_3_data_173;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_174 <= amplifier_1_0_data_174;
    end else begin
      recv_3_data_174 <= amplifier_1_3_data_174;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_175 <= amplifier_1_0_data_175;
    end else begin
      recv_3_data_175 <= amplifier_1_3_data_175;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_176 <= amplifier_1_0_data_176;
    end else begin
      recv_3_data_176 <= amplifier_1_3_data_176;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_177 <= amplifier_1_0_data_177;
    end else begin
      recv_3_data_177 <= amplifier_1_3_data_177;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_178 <= amplifier_1_0_data_178;
    end else begin
      recv_3_data_178 <= amplifier_1_3_data_178;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_179 <= amplifier_1_0_data_179;
    end else begin
      recv_3_data_179 <= amplifier_1_3_data_179;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_180 <= amplifier_1_0_data_180;
    end else begin
      recv_3_data_180 <= amplifier_1_3_data_180;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_181 <= amplifier_1_0_data_181;
    end else begin
      recv_3_data_181 <= amplifier_1_3_data_181;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_182 <= amplifier_1_0_data_182;
    end else begin
      recv_3_data_182 <= amplifier_1_3_data_182;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_183 <= amplifier_1_0_data_183;
    end else begin
      recv_3_data_183 <= amplifier_1_3_data_183;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_184 <= amplifier_1_0_data_184;
    end else begin
      recv_3_data_184 <= amplifier_1_3_data_184;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_185 <= amplifier_1_0_data_185;
    end else begin
      recv_3_data_185 <= amplifier_1_3_data_185;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_186 <= amplifier_1_0_data_186;
    end else begin
      recv_3_data_186 <= amplifier_1_3_data_186;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_187 <= amplifier_1_0_data_187;
    end else begin
      recv_3_data_187 <= amplifier_1_3_data_187;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_188 <= amplifier_1_0_data_188;
    end else begin
      recv_3_data_188 <= amplifier_1_3_data_188;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_189 <= amplifier_1_0_data_189;
    end else begin
      recv_3_data_189 <= amplifier_1_3_data_189;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_190 <= amplifier_1_0_data_190;
    end else begin
      recv_3_data_190 <= amplifier_1_3_data_190;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_191 <= amplifier_1_0_data_191;
    end else begin
      recv_3_data_191 <= amplifier_1_3_data_191;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_192 <= amplifier_1_0_data_192;
    end else begin
      recv_3_data_192 <= amplifier_1_3_data_192;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_193 <= amplifier_1_0_data_193;
    end else begin
      recv_3_data_193 <= amplifier_1_3_data_193;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_194 <= amplifier_1_0_data_194;
    end else begin
      recv_3_data_194 <= amplifier_1_3_data_194;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_195 <= amplifier_1_0_data_195;
    end else begin
      recv_3_data_195 <= amplifier_1_3_data_195;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_196 <= amplifier_1_0_data_196;
    end else begin
      recv_3_data_196 <= amplifier_1_3_data_196;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_197 <= amplifier_1_0_data_197;
    end else begin
      recv_3_data_197 <= amplifier_1_3_data_197;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_198 <= amplifier_1_0_data_198;
    end else begin
      recv_3_data_198 <= amplifier_1_3_data_198;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_199 <= amplifier_1_0_data_199;
    end else begin
      recv_3_data_199 <= amplifier_1_3_data_199;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_200 <= amplifier_1_0_data_200;
    end else begin
      recv_3_data_200 <= amplifier_1_3_data_200;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_201 <= amplifier_1_0_data_201;
    end else begin
      recv_3_data_201 <= amplifier_1_3_data_201;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_202 <= amplifier_1_0_data_202;
    end else begin
      recv_3_data_202 <= amplifier_1_3_data_202;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_203 <= amplifier_1_0_data_203;
    end else begin
      recv_3_data_203 <= amplifier_1_3_data_203;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_204 <= amplifier_1_0_data_204;
    end else begin
      recv_3_data_204 <= amplifier_1_3_data_204;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_205 <= amplifier_1_0_data_205;
    end else begin
      recv_3_data_205 <= amplifier_1_3_data_205;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_206 <= amplifier_1_0_data_206;
    end else begin
      recv_3_data_206 <= amplifier_1_3_data_206;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_207 <= amplifier_1_0_data_207;
    end else begin
      recv_3_data_207 <= amplifier_1_3_data_207;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_208 <= amplifier_1_0_data_208;
    end else begin
      recv_3_data_208 <= amplifier_1_3_data_208;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_209 <= amplifier_1_0_data_209;
    end else begin
      recv_3_data_209 <= amplifier_1_3_data_209;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_210 <= amplifier_1_0_data_210;
    end else begin
      recv_3_data_210 <= amplifier_1_3_data_210;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_211 <= amplifier_1_0_data_211;
    end else begin
      recv_3_data_211 <= amplifier_1_3_data_211;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_212 <= amplifier_1_0_data_212;
    end else begin
      recv_3_data_212 <= amplifier_1_3_data_212;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_213 <= amplifier_1_0_data_213;
    end else begin
      recv_3_data_213 <= amplifier_1_3_data_213;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_214 <= amplifier_1_0_data_214;
    end else begin
      recv_3_data_214 <= amplifier_1_3_data_214;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_215 <= amplifier_1_0_data_215;
    end else begin
      recv_3_data_215 <= amplifier_1_3_data_215;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_216 <= amplifier_1_0_data_216;
    end else begin
      recv_3_data_216 <= amplifier_1_3_data_216;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_217 <= amplifier_1_0_data_217;
    end else begin
      recv_3_data_217 <= amplifier_1_3_data_217;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_218 <= amplifier_1_0_data_218;
    end else begin
      recv_3_data_218 <= amplifier_1_3_data_218;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_219 <= amplifier_1_0_data_219;
    end else begin
      recv_3_data_219 <= amplifier_1_3_data_219;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_220 <= amplifier_1_0_data_220;
    end else begin
      recv_3_data_220 <= amplifier_1_3_data_220;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_221 <= amplifier_1_0_data_221;
    end else begin
      recv_3_data_221 <= amplifier_1_3_data_221;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_222 <= amplifier_1_0_data_222;
    end else begin
      recv_3_data_222 <= amplifier_1_3_data_222;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_223 <= amplifier_1_0_data_223;
    end else begin
      recv_3_data_223 <= amplifier_1_3_data_223;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_224 <= amplifier_1_0_data_224;
    end else begin
      recv_3_data_224 <= amplifier_1_3_data_224;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_225 <= amplifier_1_0_data_225;
    end else begin
      recv_3_data_225 <= amplifier_1_3_data_225;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_226 <= amplifier_1_0_data_226;
    end else begin
      recv_3_data_226 <= amplifier_1_3_data_226;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_227 <= amplifier_1_0_data_227;
    end else begin
      recv_3_data_227 <= amplifier_1_3_data_227;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_228 <= amplifier_1_0_data_228;
    end else begin
      recv_3_data_228 <= amplifier_1_3_data_228;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_229 <= amplifier_1_0_data_229;
    end else begin
      recv_3_data_229 <= amplifier_1_3_data_229;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_230 <= amplifier_1_0_data_230;
    end else begin
      recv_3_data_230 <= amplifier_1_3_data_230;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_231 <= amplifier_1_0_data_231;
    end else begin
      recv_3_data_231 <= amplifier_1_3_data_231;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_232 <= amplifier_1_0_data_232;
    end else begin
      recv_3_data_232 <= amplifier_1_3_data_232;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_233 <= amplifier_1_0_data_233;
    end else begin
      recv_3_data_233 <= amplifier_1_3_data_233;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_234 <= amplifier_1_0_data_234;
    end else begin
      recv_3_data_234 <= amplifier_1_3_data_234;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_235 <= amplifier_1_0_data_235;
    end else begin
      recv_3_data_235 <= amplifier_1_3_data_235;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_236 <= amplifier_1_0_data_236;
    end else begin
      recv_3_data_236 <= amplifier_1_3_data_236;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_237 <= amplifier_1_0_data_237;
    end else begin
      recv_3_data_237 <= amplifier_1_3_data_237;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_238 <= amplifier_1_0_data_238;
    end else begin
      recv_3_data_238 <= amplifier_1_3_data_238;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_239 <= amplifier_1_0_data_239;
    end else begin
      recv_3_data_239 <= amplifier_1_3_data_239;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_240 <= amplifier_1_0_data_240;
    end else begin
      recv_3_data_240 <= amplifier_1_3_data_240;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_241 <= amplifier_1_0_data_241;
    end else begin
      recv_3_data_241 <= amplifier_1_3_data_241;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_242 <= amplifier_1_0_data_242;
    end else begin
      recv_3_data_242 <= amplifier_1_3_data_242;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_243 <= amplifier_1_0_data_243;
    end else begin
      recv_3_data_243 <= amplifier_1_3_data_243;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_244 <= amplifier_1_0_data_244;
    end else begin
      recv_3_data_244 <= amplifier_1_3_data_244;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_245 <= amplifier_1_0_data_245;
    end else begin
      recv_3_data_245 <= amplifier_1_3_data_245;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_246 <= amplifier_1_0_data_246;
    end else begin
      recv_3_data_246 <= amplifier_1_3_data_246;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_247 <= amplifier_1_0_data_247;
    end else begin
      recv_3_data_247 <= amplifier_1_3_data_247;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_248 <= amplifier_1_0_data_248;
    end else begin
      recv_3_data_248 <= amplifier_1_3_data_248;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_249 <= amplifier_1_0_data_249;
    end else begin
      recv_3_data_249 <= amplifier_1_3_data_249;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_250 <= amplifier_1_0_data_250;
    end else begin
      recv_3_data_250 <= amplifier_1_3_data_250;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_251 <= amplifier_1_0_data_251;
    end else begin
      recv_3_data_251 <= amplifier_1_3_data_251;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_252 <= amplifier_1_0_data_252;
    end else begin
      recv_3_data_252 <= amplifier_1_3_data_252;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_253 <= amplifier_1_0_data_253;
    end else begin
      recv_3_data_253 <= amplifier_1_3_data_253;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_254 <= amplifier_1_0_data_254;
    end else begin
      recv_3_data_254 <= amplifier_1_3_data_254;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_data_255 <= amplifier_1_0_data_255;
    end else begin
      recv_3_data_255 <= amplifier_1_3_data_255;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_header_0 <= amplifier_1_0_header_0;
    end else begin
      recv_3_header_0 <= amplifier_1_3_header_0;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_header_1 <= amplifier_1_0_header_1;
    end else begin
      recv_3_header_1 <= amplifier_1_3_header_1;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_header_2 <= amplifier_1_0_header_2;
    end else begin
      recv_3_header_2 <= amplifier_1_3_header_2;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_header_3 <= amplifier_1_0_header_3;
    end else begin
      recv_3_header_3 <= amplifier_1_3_header_3;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_header_4 <= amplifier_1_0_header_4;
    end else begin
      recv_3_header_4 <= amplifier_1_3_header_4;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_header_5 <= amplifier_1_0_header_5;
    end else begin
      recv_3_header_5 <= amplifier_1_3_header_5;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_header_6 <= amplifier_1_0_header_6;
    end else begin
      recv_3_header_6 <= amplifier_1_3_header_6;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_header_7 <= amplifier_1_0_header_7;
    end else begin
      recv_3_header_7 <= amplifier_1_3_header_7;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_header_8 <= amplifier_1_0_header_8;
    end else begin
      recv_3_header_8 <= amplifier_1_3_header_8;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_header_9 <= amplifier_1_0_header_9;
    end else begin
      recv_3_header_9 <= amplifier_1_3_header_9;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_header_10 <= amplifier_1_0_header_10;
    end else begin
      recv_3_header_10 <= amplifier_1_3_header_10;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_header_11 <= amplifier_1_0_header_11;
    end else begin
      recv_3_header_11 <= amplifier_1_3_header_11;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_header_12 <= amplifier_1_0_header_12;
    end else begin
      recv_3_header_12 <= amplifier_1_3_header_12;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_header_13 <= amplifier_1_0_header_13;
    end else begin
      recv_3_header_13 <= amplifier_1_3_header_13;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_header_14 <= amplifier_1_0_header_14;
    end else begin
      recv_3_header_14 <= amplifier_1_3_header_14;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_header_15 <= amplifier_1_0_header_15;
    end else begin
      recv_3_header_15 <= amplifier_1_3_header_15;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_parse_current_state <= amplifier_1_0_parse_current_state;
    end else begin
      recv_3_parse_current_state <= amplifier_1_3_parse_current_state;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_parse_current_offset <= amplifier_1_0_parse_current_offset;
    end else begin
      recv_3_parse_current_offset <= amplifier_1_3_parse_current_offset;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_parse_transition_field <= amplifier_1_0_parse_transition_field;
    end else begin
      recv_3_parse_transition_field <= amplifier_1_3_parse_transition_field;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_next_processor_id <= amplifier_1_0_next_processor_id;
    end else begin
      recv_3_next_processor_id <= amplifier_1_3_next_processor_id;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_next_config_id <= amplifier_1_0_next_config_id;
    end else begin
      recv_3_next_config_id <= amplifier_1_3_next_config_id;
    end
    if (_recv_3_T) begin // @[ipsa.scala 155:23]
      recv_3_is_valid_processor <= amplifier_1_0_is_valid_processor;
    end else begin
      recv_3_is_valid_processor <= amplifier_1_3_is_valid_processor;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_0 <= init_io_pipe_phv_out_data_0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_0 <= trans_1_io_pipe_phv_out_data_0;
    end else begin
      amplifier_0_0_data_0 <= trans_0_io_pipe_phv_out_data_0;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_1 <= init_io_pipe_phv_out_data_1; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_1 <= trans_1_io_pipe_phv_out_data_1;
    end else begin
      amplifier_0_0_data_1 <= trans_0_io_pipe_phv_out_data_1;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_2 <= init_io_pipe_phv_out_data_2; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_2 <= trans_1_io_pipe_phv_out_data_2;
    end else begin
      amplifier_0_0_data_2 <= trans_0_io_pipe_phv_out_data_2;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_3 <= init_io_pipe_phv_out_data_3; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_3 <= trans_1_io_pipe_phv_out_data_3;
    end else begin
      amplifier_0_0_data_3 <= trans_0_io_pipe_phv_out_data_3;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_4 <= init_io_pipe_phv_out_data_4; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_4 <= trans_1_io_pipe_phv_out_data_4;
    end else begin
      amplifier_0_0_data_4 <= trans_0_io_pipe_phv_out_data_4;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_5 <= init_io_pipe_phv_out_data_5; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_5 <= trans_1_io_pipe_phv_out_data_5;
    end else begin
      amplifier_0_0_data_5 <= trans_0_io_pipe_phv_out_data_5;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_6 <= init_io_pipe_phv_out_data_6; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_6 <= trans_1_io_pipe_phv_out_data_6;
    end else begin
      amplifier_0_0_data_6 <= trans_0_io_pipe_phv_out_data_6;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_7 <= init_io_pipe_phv_out_data_7; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_7 <= trans_1_io_pipe_phv_out_data_7;
    end else begin
      amplifier_0_0_data_7 <= trans_0_io_pipe_phv_out_data_7;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_8 <= init_io_pipe_phv_out_data_8; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_8 <= trans_1_io_pipe_phv_out_data_8;
    end else begin
      amplifier_0_0_data_8 <= trans_0_io_pipe_phv_out_data_8;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_9 <= init_io_pipe_phv_out_data_9; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_9 <= trans_1_io_pipe_phv_out_data_9;
    end else begin
      amplifier_0_0_data_9 <= trans_0_io_pipe_phv_out_data_9;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_10 <= init_io_pipe_phv_out_data_10; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_10 <= trans_1_io_pipe_phv_out_data_10;
    end else begin
      amplifier_0_0_data_10 <= trans_0_io_pipe_phv_out_data_10;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_11 <= init_io_pipe_phv_out_data_11; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_11 <= trans_1_io_pipe_phv_out_data_11;
    end else begin
      amplifier_0_0_data_11 <= trans_0_io_pipe_phv_out_data_11;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_12 <= init_io_pipe_phv_out_data_12; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_12 <= trans_1_io_pipe_phv_out_data_12;
    end else begin
      amplifier_0_0_data_12 <= trans_0_io_pipe_phv_out_data_12;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_13 <= init_io_pipe_phv_out_data_13; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_13 <= trans_1_io_pipe_phv_out_data_13;
    end else begin
      amplifier_0_0_data_13 <= trans_0_io_pipe_phv_out_data_13;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_14 <= init_io_pipe_phv_out_data_14; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_14 <= trans_1_io_pipe_phv_out_data_14;
    end else begin
      amplifier_0_0_data_14 <= trans_0_io_pipe_phv_out_data_14;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_15 <= init_io_pipe_phv_out_data_15; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_15 <= trans_1_io_pipe_phv_out_data_15;
    end else begin
      amplifier_0_0_data_15 <= trans_0_io_pipe_phv_out_data_15;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_16 <= init_io_pipe_phv_out_data_16; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_16 <= trans_1_io_pipe_phv_out_data_16;
    end else begin
      amplifier_0_0_data_16 <= trans_0_io_pipe_phv_out_data_16;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_17 <= init_io_pipe_phv_out_data_17; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_17 <= trans_1_io_pipe_phv_out_data_17;
    end else begin
      amplifier_0_0_data_17 <= trans_0_io_pipe_phv_out_data_17;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_18 <= init_io_pipe_phv_out_data_18; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_18 <= trans_1_io_pipe_phv_out_data_18;
    end else begin
      amplifier_0_0_data_18 <= trans_0_io_pipe_phv_out_data_18;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_19 <= init_io_pipe_phv_out_data_19; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_19 <= trans_1_io_pipe_phv_out_data_19;
    end else begin
      amplifier_0_0_data_19 <= trans_0_io_pipe_phv_out_data_19;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_20 <= init_io_pipe_phv_out_data_20; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_20 <= trans_1_io_pipe_phv_out_data_20;
    end else begin
      amplifier_0_0_data_20 <= trans_0_io_pipe_phv_out_data_20;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_21 <= init_io_pipe_phv_out_data_21; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_21 <= trans_1_io_pipe_phv_out_data_21;
    end else begin
      amplifier_0_0_data_21 <= trans_0_io_pipe_phv_out_data_21;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_22 <= init_io_pipe_phv_out_data_22; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_22 <= trans_1_io_pipe_phv_out_data_22;
    end else begin
      amplifier_0_0_data_22 <= trans_0_io_pipe_phv_out_data_22;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_23 <= init_io_pipe_phv_out_data_23; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_23 <= trans_1_io_pipe_phv_out_data_23;
    end else begin
      amplifier_0_0_data_23 <= trans_0_io_pipe_phv_out_data_23;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_24 <= init_io_pipe_phv_out_data_24; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_24 <= trans_1_io_pipe_phv_out_data_24;
    end else begin
      amplifier_0_0_data_24 <= trans_0_io_pipe_phv_out_data_24;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_25 <= init_io_pipe_phv_out_data_25; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_25 <= trans_1_io_pipe_phv_out_data_25;
    end else begin
      amplifier_0_0_data_25 <= trans_0_io_pipe_phv_out_data_25;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_26 <= init_io_pipe_phv_out_data_26; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_26 <= trans_1_io_pipe_phv_out_data_26;
    end else begin
      amplifier_0_0_data_26 <= trans_0_io_pipe_phv_out_data_26;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_27 <= init_io_pipe_phv_out_data_27; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_27 <= trans_1_io_pipe_phv_out_data_27;
    end else begin
      amplifier_0_0_data_27 <= trans_0_io_pipe_phv_out_data_27;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_28 <= init_io_pipe_phv_out_data_28; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_28 <= trans_1_io_pipe_phv_out_data_28;
    end else begin
      amplifier_0_0_data_28 <= trans_0_io_pipe_phv_out_data_28;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_29 <= init_io_pipe_phv_out_data_29; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_29 <= trans_1_io_pipe_phv_out_data_29;
    end else begin
      amplifier_0_0_data_29 <= trans_0_io_pipe_phv_out_data_29;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_30 <= init_io_pipe_phv_out_data_30; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_30 <= trans_1_io_pipe_phv_out_data_30;
    end else begin
      amplifier_0_0_data_30 <= trans_0_io_pipe_phv_out_data_30;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_31 <= init_io_pipe_phv_out_data_31; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_31 <= trans_1_io_pipe_phv_out_data_31;
    end else begin
      amplifier_0_0_data_31 <= trans_0_io_pipe_phv_out_data_31;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_32 <= init_io_pipe_phv_out_data_32; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_32 <= trans_1_io_pipe_phv_out_data_32;
    end else begin
      amplifier_0_0_data_32 <= trans_0_io_pipe_phv_out_data_32;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_33 <= init_io_pipe_phv_out_data_33; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_33 <= trans_1_io_pipe_phv_out_data_33;
    end else begin
      amplifier_0_0_data_33 <= trans_0_io_pipe_phv_out_data_33;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_34 <= init_io_pipe_phv_out_data_34; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_34 <= trans_1_io_pipe_phv_out_data_34;
    end else begin
      amplifier_0_0_data_34 <= trans_0_io_pipe_phv_out_data_34;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_35 <= init_io_pipe_phv_out_data_35; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_35 <= trans_1_io_pipe_phv_out_data_35;
    end else begin
      amplifier_0_0_data_35 <= trans_0_io_pipe_phv_out_data_35;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_36 <= init_io_pipe_phv_out_data_36; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_36 <= trans_1_io_pipe_phv_out_data_36;
    end else begin
      amplifier_0_0_data_36 <= trans_0_io_pipe_phv_out_data_36;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_37 <= init_io_pipe_phv_out_data_37; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_37 <= trans_1_io_pipe_phv_out_data_37;
    end else begin
      amplifier_0_0_data_37 <= trans_0_io_pipe_phv_out_data_37;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_38 <= init_io_pipe_phv_out_data_38; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_38 <= trans_1_io_pipe_phv_out_data_38;
    end else begin
      amplifier_0_0_data_38 <= trans_0_io_pipe_phv_out_data_38;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_39 <= init_io_pipe_phv_out_data_39; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_39 <= trans_1_io_pipe_phv_out_data_39;
    end else begin
      amplifier_0_0_data_39 <= trans_0_io_pipe_phv_out_data_39;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_40 <= init_io_pipe_phv_out_data_40; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_40 <= trans_1_io_pipe_phv_out_data_40;
    end else begin
      amplifier_0_0_data_40 <= trans_0_io_pipe_phv_out_data_40;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_41 <= init_io_pipe_phv_out_data_41; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_41 <= trans_1_io_pipe_phv_out_data_41;
    end else begin
      amplifier_0_0_data_41 <= trans_0_io_pipe_phv_out_data_41;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_42 <= init_io_pipe_phv_out_data_42; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_42 <= trans_1_io_pipe_phv_out_data_42;
    end else begin
      amplifier_0_0_data_42 <= trans_0_io_pipe_phv_out_data_42;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_43 <= init_io_pipe_phv_out_data_43; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_43 <= trans_1_io_pipe_phv_out_data_43;
    end else begin
      amplifier_0_0_data_43 <= trans_0_io_pipe_phv_out_data_43;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_44 <= init_io_pipe_phv_out_data_44; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_44 <= trans_1_io_pipe_phv_out_data_44;
    end else begin
      amplifier_0_0_data_44 <= trans_0_io_pipe_phv_out_data_44;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_45 <= init_io_pipe_phv_out_data_45; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_45 <= trans_1_io_pipe_phv_out_data_45;
    end else begin
      amplifier_0_0_data_45 <= trans_0_io_pipe_phv_out_data_45;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_46 <= init_io_pipe_phv_out_data_46; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_46 <= trans_1_io_pipe_phv_out_data_46;
    end else begin
      amplifier_0_0_data_46 <= trans_0_io_pipe_phv_out_data_46;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_47 <= init_io_pipe_phv_out_data_47; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_47 <= trans_1_io_pipe_phv_out_data_47;
    end else begin
      amplifier_0_0_data_47 <= trans_0_io_pipe_phv_out_data_47;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_48 <= init_io_pipe_phv_out_data_48; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_48 <= trans_1_io_pipe_phv_out_data_48;
    end else begin
      amplifier_0_0_data_48 <= trans_0_io_pipe_phv_out_data_48;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_49 <= init_io_pipe_phv_out_data_49; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_49 <= trans_1_io_pipe_phv_out_data_49;
    end else begin
      amplifier_0_0_data_49 <= trans_0_io_pipe_phv_out_data_49;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_50 <= init_io_pipe_phv_out_data_50; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_50 <= trans_1_io_pipe_phv_out_data_50;
    end else begin
      amplifier_0_0_data_50 <= trans_0_io_pipe_phv_out_data_50;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_51 <= init_io_pipe_phv_out_data_51; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_51 <= trans_1_io_pipe_phv_out_data_51;
    end else begin
      amplifier_0_0_data_51 <= trans_0_io_pipe_phv_out_data_51;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_52 <= init_io_pipe_phv_out_data_52; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_52 <= trans_1_io_pipe_phv_out_data_52;
    end else begin
      amplifier_0_0_data_52 <= trans_0_io_pipe_phv_out_data_52;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_53 <= init_io_pipe_phv_out_data_53; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_53 <= trans_1_io_pipe_phv_out_data_53;
    end else begin
      amplifier_0_0_data_53 <= trans_0_io_pipe_phv_out_data_53;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_54 <= init_io_pipe_phv_out_data_54; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_54 <= trans_1_io_pipe_phv_out_data_54;
    end else begin
      amplifier_0_0_data_54 <= trans_0_io_pipe_phv_out_data_54;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_55 <= init_io_pipe_phv_out_data_55; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_55 <= trans_1_io_pipe_phv_out_data_55;
    end else begin
      amplifier_0_0_data_55 <= trans_0_io_pipe_phv_out_data_55;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_56 <= init_io_pipe_phv_out_data_56; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_56 <= trans_1_io_pipe_phv_out_data_56;
    end else begin
      amplifier_0_0_data_56 <= trans_0_io_pipe_phv_out_data_56;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_57 <= init_io_pipe_phv_out_data_57; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_57 <= trans_1_io_pipe_phv_out_data_57;
    end else begin
      amplifier_0_0_data_57 <= trans_0_io_pipe_phv_out_data_57;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_58 <= init_io_pipe_phv_out_data_58; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_58 <= trans_1_io_pipe_phv_out_data_58;
    end else begin
      amplifier_0_0_data_58 <= trans_0_io_pipe_phv_out_data_58;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_59 <= init_io_pipe_phv_out_data_59; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_59 <= trans_1_io_pipe_phv_out_data_59;
    end else begin
      amplifier_0_0_data_59 <= trans_0_io_pipe_phv_out_data_59;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_60 <= init_io_pipe_phv_out_data_60; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_60 <= trans_1_io_pipe_phv_out_data_60;
    end else begin
      amplifier_0_0_data_60 <= trans_0_io_pipe_phv_out_data_60;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_61 <= init_io_pipe_phv_out_data_61; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_61 <= trans_1_io_pipe_phv_out_data_61;
    end else begin
      amplifier_0_0_data_61 <= trans_0_io_pipe_phv_out_data_61;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_62 <= init_io_pipe_phv_out_data_62; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_62 <= trans_1_io_pipe_phv_out_data_62;
    end else begin
      amplifier_0_0_data_62 <= trans_0_io_pipe_phv_out_data_62;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_63 <= init_io_pipe_phv_out_data_63; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_63 <= trans_1_io_pipe_phv_out_data_63;
    end else begin
      amplifier_0_0_data_63 <= trans_0_io_pipe_phv_out_data_63;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_64 <= init_io_pipe_phv_out_data_64; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_64 <= trans_1_io_pipe_phv_out_data_64;
    end else begin
      amplifier_0_0_data_64 <= trans_0_io_pipe_phv_out_data_64;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_65 <= init_io_pipe_phv_out_data_65; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_65 <= trans_1_io_pipe_phv_out_data_65;
    end else begin
      amplifier_0_0_data_65 <= trans_0_io_pipe_phv_out_data_65;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_66 <= init_io_pipe_phv_out_data_66; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_66 <= trans_1_io_pipe_phv_out_data_66;
    end else begin
      amplifier_0_0_data_66 <= trans_0_io_pipe_phv_out_data_66;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_67 <= init_io_pipe_phv_out_data_67; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_67 <= trans_1_io_pipe_phv_out_data_67;
    end else begin
      amplifier_0_0_data_67 <= trans_0_io_pipe_phv_out_data_67;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_68 <= init_io_pipe_phv_out_data_68; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_68 <= trans_1_io_pipe_phv_out_data_68;
    end else begin
      amplifier_0_0_data_68 <= trans_0_io_pipe_phv_out_data_68;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_69 <= init_io_pipe_phv_out_data_69; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_69 <= trans_1_io_pipe_phv_out_data_69;
    end else begin
      amplifier_0_0_data_69 <= trans_0_io_pipe_phv_out_data_69;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_70 <= init_io_pipe_phv_out_data_70; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_70 <= trans_1_io_pipe_phv_out_data_70;
    end else begin
      amplifier_0_0_data_70 <= trans_0_io_pipe_phv_out_data_70;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_71 <= init_io_pipe_phv_out_data_71; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_71 <= trans_1_io_pipe_phv_out_data_71;
    end else begin
      amplifier_0_0_data_71 <= trans_0_io_pipe_phv_out_data_71;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_72 <= init_io_pipe_phv_out_data_72; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_72 <= trans_1_io_pipe_phv_out_data_72;
    end else begin
      amplifier_0_0_data_72 <= trans_0_io_pipe_phv_out_data_72;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_73 <= init_io_pipe_phv_out_data_73; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_73 <= trans_1_io_pipe_phv_out_data_73;
    end else begin
      amplifier_0_0_data_73 <= trans_0_io_pipe_phv_out_data_73;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_74 <= init_io_pipe_phv_out_data_74; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_74 <= trans_1_io_pipe_phv_out_data_74;
    end else begin
      amplifier_0_0_data_74 <= trans_0_io_pipe_phv_out_data_74;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_75 <= init_io_pipe_phv_out_data_75; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_75 <= trans_1_io_pipe_phv_out_data_75;
    end else begin
      amplifier_0_0_data_75 <= trans_0_io_pipe_phv_out_data_75;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_76 <= init_io_pipe_phv_out_data_76; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_76 <= trans_1_io_pipe_phv_out_data_76;
    end else begin
      amplifier_0_0_data_76 <= trans_0_io_pipe_phv_out_data_76;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_77 <= init_io_pipe_phv_out_data_77; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_77 <= trans_1_io_pipe_phv_out_data_77;
    end else begin
      amplifier_0_0_data_77 <= trans_0_io_pipe_phv_out_data_77;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_78 <= init_io_pipe_phv_out_data_78; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_78 <= trans_1_io_pipe_phv_out_data_78;
    end else begin
      amplifier_0_0_data_78 <= trans_0_io_pipe_phv_out_data_78;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_79 <= init_io_pipe_phv_out_data_79; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_79 <= trans_1_io_pipe_phv_out_data_79;
    end else begin
      amplifier_0_0_data_79 <= trans_0_io_pipe_phv_out_data_79;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_80 <= init_io_pipe_phv_out_data_80; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_80 <= trans_1_io_pipe_phv_out_data_80;
    end else begin
      amplifier_0_0_data_80 <= trans_0_io_pipe_phv_out_data_80;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_81 <= init_io_pipe_phv_out_data_81; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_81 <= trans_1_io_pipe_phv_out_data_81;
    end else begin
      amplifier_0_0_data_81 <= trans_0_io_pipe_phv_out_data_81;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_82 <= init_io_pipe_phv_out_data_82; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_82 <= trans_1_io_pipe_phv_out_data_82;
    end else begin
      amplifier_0_0_data_82 <= trans_0_io_pipe_phv_out_data_82;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_83 <= init_io_pipe_phv_out_data_83; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_83 <= trans_1_io_pipe_phv_out_data_83;
    end else begin
      amplifier_0_0_data_83 <= trans_0_io_pipe_phv_out_data_83;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_84 <= init_io_pipe_phv_out_data_84; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_84 <= trans_1_io_pipe_phv_out_data_84;
    end else begin
      amplifier_0_0_data_84 <= trans_0_io_pipe_phv_out_data_84;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_85 <= init_io_pipe_phv_out_data_85; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_85 <= trans_1_io_pipe_phv_out_data_85;
    end else begin
      amplifier_0_0_data_85 <= trans_0_io_pipe_phv_out_data_85;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_86 <= init_io_pipe_phv_out_data_86; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_86 <= trans_1_io_pipe_phv_out_data_86;
    end else begin
      amplifier_0_0_data_86 <= trans_0_io_pipe_phv_out_data_86;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_87 <= init_io_pipe_phv_out_data_87; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_87 <= trans_1_io_pipe_phv_out_data_87;
    end else begin
      amplifier_0_0_data_87 <= trans_0_io_pipe_phv_out_data_87;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_88 <= init_io_pipe_phv_out_data_88; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_88 <= trans_1_io_pipe_phv_out_data_88;
    end else begin
      amplifier_0_0_data_88 <= trans_0_io_pipe_phv_out_data_88;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_89 <= init_io_pipe_phv_out_data_89; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_89 <= trans_1_io_pipe_phv_out_data_89;
    end else begin
      amplifier_0_0_data_89 <= trans_0_io_pipe_phv_out_data_89;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_90 <= init_io_pipe_phv_out_data_90; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_90 <= trans_1_io_pipe_phv_out_data_90;
    end else begin
      amplifier_0_0_data_90 <= trans_0_io_pipe_phv_out_data_90;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_91 <= init_io_pipe_phv_out_data_91; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_91 <= trans_1_io_pipe_phv_out_data_91;
    end else begin
      amplifier_0_0_data_91 <= trans_0_io_pipe_phv_out_data_91;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_92 <= init_io_pipe_phv_out_data_92; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_92 <= trans_1_io_pipe_phv_out_data_92;
    end else begin
      amplifier_0_0_data_92 <= trans_0_io_pipe_phv_out_data_92;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_93 <= init_io_pipe_phv_out_data_93; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_93 <= trans_1_io_pipe_phv_out_data_93;
    end else begin
      amplifier_0_0_data_93 <= trans_0_io_pipe_phv_out_data_93;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_94 <= init_io_pipe_phv_out_data_94; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_94 <= trans_1_io_pipe_phv_out_data_94;
    end else begin
      amplifier_0_0_data_94 <= trans_0_io_pipe_phv_out_data_94;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_95 <= init_io_pipe_phv_out_data_95; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_95 <= trans_1_io_pipe_phv_out_data_95;
    end else begin
      amplifier_0_0_data_95 <= trans_0_io_pipe_phv_out_data_95;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_96 <= init_io_pipe_phv_out_data_96; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_96 <= trans_1_io_pipe_phv_out_data_96;
    end else begin
      amplifier_0_0_data_96 <= trans_0_io_pipe_phv_out_data_96;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_97 <= init_io_pipe_phv_out_data_97; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_97 <= trans_1_io_pipe_phv_out_data_97;
    end else begin
      amplifier_0_0_data_97 <= trans_0_io_pipe_phv_out_data_97;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_98 <= init_io_pipe_phv_out_data_98; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_98 <= trans_1_io_pipe_phv_out_data_98;
    end else begin
      amplifier_0_0_data_98 <= trans_0_io_pipe_phv_out_data_98;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_99 <= init_io_pipe_phv_out_data_99; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_99 <= trans_1_io_pipe_phv_out_data_99;
    end else begin
      amplifier_0_0_data_99 <= trans_0_io_pipe_phv_out_data_99;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_100 <= init_io_pipe_phv_out_data_100; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_100 <= trans_1_io_pipe_phv_out_data_100;
    end else begin
      amplifier_0_0_data_100 <= trans_0_io_pipe_phv_out_data_100;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_101 <= init_io_pipe_phv_out_data_101; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_101 <= trans_1_io_pipe_phv_out_data_101;
    end else begin
      amplifier_0_0_data_101 <= trans_0_io_pipe_phv_out_data_101;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_102 <= init_io_pipe_phv_out_data_102; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_102 <= trans_1_io_pipe_phv_out_data_102;
    end else begin
      amplifier_0_0_data_102 <= trans_0_io_pipe_phv_out_data_102;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_103 <= init_io_pipe_phv_out_data_103; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_103 <= trans_1_io_pipe_phv_out_data_103;
    end else begin
      amplifier_0_0_data_103 <= trans_0_io_pipe_phv_out_data_103;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_104 <= init_io_pipe_phv_out_data_104; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_104 <= trans_1_io_pipe_phv_out_data_104;
    end else begin
      amplifier_0_0_data_104 <= trans_0_io_pipe_phv_out_data_104;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_105 <= init_io_pipe_phv_out_data_105; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_105 <= trans_1_io_pipe_phv_out_data_105;
    end else begin
      amplifier_0_0_data_105 <= trans_0_io_pipe_phv_out_data_105;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_106 <= init_io_pipe_phv_out_data_106; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_106 <= trans_1_io_pipe_phv_out_data_106;
    end else begin
      amplifier_0_0_data_106 <= trans_0_io_pipe_phv_out_data_106;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_107 <= init_io_pipe_phv_out_data_107; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_107 <= trans_1_io_pipe_phv_out_data_107;
    end else begin
      amplifier_0_0_data_107 <= trans_0_io_pipe_phv_out_data_107;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_108 <= init_io_pipe_phv_out_data_108; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_108 <= trans_1_io_pipe_phv_out_data_108;
    end else begin
      amplifier_0_0_data_108 <= trans_0_io_pipe_phv_out_data_108;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_109 <= init_io_pipe_phv_out_data_109; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_109 <= trans_1_io_pipe_phv_out_data_109;
    end else begin
      amplifier_0_0_data_109 <= trans_0_io_pipe_phv_out_data_109;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_110 <= init_io_pipe_phv_out_data_110; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_110 <= trans_1_io_pipe_phv_out_data_110;
    end else begin
      amplifier_0_0_data_110 <= trans_0_io_pipe_phv_out_data_110;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_111 <= init_io_pipe_phv_out_data_111; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_111 <= trans_1_io_pipe_phv_out_data_111;
    end else begin
      amplifier_0_0_data_111 <= trans_0_io_pipe_phv_out_data_111;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_112 <= init_io_pipe_phv_out_data_112; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_112 <= trans_1_io_pipe_phv_out_data_112;
    end else begin
      amplifier_0_0_data_112 <= trans_0_io_pipe_phv_out_data_112;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_113 <= init_io_pipe_phv_out_data_113; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_113 <= trans_1_io_pipe_phv_out_data_113;
    end else begin
      amplifier_0_0_data_113 <= trans_0_io_pipe_phv_out_data_113;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_114 <= init_io_pipe_phv_out_data_114; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_114 <= trans_1_io_pipe_phv_out_data_114;
    end else begin
      amplifier_0_0_data_114 <= trans_0_io_pipe_phv_out_data_114;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_115 <= init_io_pipe_phv_out_data_115; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_115 <= trans_1_io_pipe_phv_out_data_115;
    end else begin
      amplifier_0_0_data_115 <= trans_0_io_pipe_phv_out_data_115;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_116 <= init_io_pipe_phv_out_data_116; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_116 <= trans_1_io_pipe_phv_out_data_116;
    end else begin
      amplifier_0_0_data_116 <= trans_0_io_pipe_phv_out_data_116;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_117 <= init_io_pipe_phv_out_data_117; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_117 <= trans_1_io_pipe_phv_out_data_117;
    end else begin
      amplifier_0_0_data_117 <= trans_0_io_pipe_phv_out_data_117;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_118 <= init_io_pipe_phv_out_data_118; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_118 <= trans_1_io_pipe_phv_out_data_118;
    end else begin
      amplifier_0_0_data_118 <= trans_0_io_pipe_phv_out_data_118;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_119 <= init_io_pipe_phv_out_data_119; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_119 <= trans_1_io_pipe_phv_out_data_119;
    end else begin
      amplifier_0_0_data_119 <= trans_0_io_pipe_phv_out_data_119;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_120 <= init_io_pipe_phv_out_data_120; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_120 <= trans_1_io_pipe_phv_out_data_120;
    end else begin
      amplifier_0_0_data_120 <= trans_0_io_pipe_phv_out_data_120;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_121 <= init_io_pipe_phv_out_data_121; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_121 <= trans_1_io_pipe_phv_out_data_121;
    end else begin
      amplifier_0_0_data_121 <= trans_0_io_pipe_phv_out_data_121;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_122 <= init_io_pipe_phv_out_data_122; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_122 <= trans_1_io_pipe_phv_out_data_122;
    end else begin
      amplifier_0_0_data_122 <= trans_0_io_pipe_phv_out_data_122;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_123 <= init_io_pipe_phv_out_data_123; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_123 <= trans_1_io_pipe_phv_out_data_123;
    end else begin
      amplifier_0_0_data_123 <= trans_0_io_pipe_phv_out_data_123;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_124 <= init_io_pipe_phv_out_data_124; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_124 <= trans_1_io_pipe_phv_out_data_124;
    end else begin
      amplifier_0_0_data_124 <= trans_0_io_pipe_phv_out_data_124;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_125 <= init_io_pipe_phv_out_data_125; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_125 <= trans_1_io_pipe_phv_out_data_125;
    end else begin
      amplifier_0_0_data_125 <= trans_0_io_pipe_phv_out_data_125;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_126 <= init_io_pipe_phv_out_data_126; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_126 <= trans_1_io_pipe_phv_out_data_126;
    end else begin
      amplifier_0_0_data_126 <= trans_0_io_pipe_phv_out_data_126;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_127 <= init_io_pipe_phv_out_data_127; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_127 <= trans_1_io_pipe_phv_out_data_127;
    end else begin
      amplifier_0_0_data_127 <= trans_0_io_pipe_phv_out_data_127;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_128 <= init_io_pipe_phv_out_data_128; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_128 <= trans_1_io_pipe_phv_out_data_128;
    end else begin
      amplifier_0_0_data_128 <= trans_0_io_pipe_phv_out_data_128;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_129 <= init_io_pipe_phv_out_data_129; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_129 <= trans_1_io_pipe_phv_out_data_129;
    end else begin
      amplifier_0_0_data_129 <= trans_0_io_pipe_phv_out_data_129;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_130 <= init_io_pipe_phv_out_data_130; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_130 <= trans_1_io_pipe_phv_out_data_130;
    end else begin
      amplifier_0_0_data_130 <= trans_0_io_pipe_phv_out_data_130;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_131 <= init_io_pipe_phv_out_data_131; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_131 <= trans_1_io_pipe_phv_out_data_131;
    end else begin
      amplifier_0_0_data_131 <= trans_0_io_pipe_phv_out_data_131;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_132 <= init_io_pipe_phv_out_data_132; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_132 <= trans_1_io_pipe_phv_out_data_132;
    end else begin
      amplifier_0_0_data_132 <= trans_0_io_pipe_phv_out_data_132;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_133 <= init_io_pipe_phv_out_data_133; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_133 <= trans_1_io_pipe_phv_out_data_133;
    end else begin
      amplifier_0_0_data_133 <= trans_0_io_pipe_phv_out_data_133;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_134 <= init_io_pipe_phv_out_data_134; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_134 <= trans_1_io_pipe_phv_out_data_134;
    end else begin
      amplifier_0_0_data_134 <= trans_0_io_pipe_phv_out_data_134;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_135 <= init_io_pipe_phv_out_data_135; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_135 <= trans_1_io_pipe_phv_out_data_135;
    end else begin
      amplifier_0_0_data_135 <= trans_0_io_pipe_phv_out_data_135;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_136 <= init_io_pipe_phv_out_data_136; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_136 <= trans_1_io_pipe_phv_out_data_136;
    end else begin
      amplifier_0_0_data_136 <= trans_0_io_pipe_phv_out_data_136;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_137 <= init_io_pipe_phv_out_data_137; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_137 <= trans_1_io_pipe_phv_out_data_137;
    end else begin
      amplifier_0_0_data_137 <= trans_0_io_pipe_phv_out_data_137;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_138 <= init_io_pipe_phv_out_data_138; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_138 <= trans_1_io_pipe_phv_out_data_138;
    end else begin
      amplifier_0_0_data_138 <= trans_0_io_pipe_phv_out_data_138;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_139 <= init_io_pipe_phv_out_data_139; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_139 <= trans_1_io_pipe_phv_out_data_139;
    end else begin
      amplifier_0_0_data_139 <= trans_0_io_pipe_phv_out_data_139;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_140 <= init_io_pipe_phv_out_data_140; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_140 <= trans_1_io_pipe_phv_out_data_140;
    end else begin
      amplifier_0_0_data_140 <= trans_0_io_pipe_phv_out_data_140;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_141 <= init_io_pipe_phv_out_data_141; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_141 <= trans_1_io_pipe_phv_out_data_141;
    end else begin
      amplifier_0_0_data_141 <= trans_0_io_pipe_phv_out_data_141;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_142 <= init_io_pipe_phv_out_data_142; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_142 <= trans_1_io_pipe_phv_out_data_142;
    end else begin
      amplifier_0_0_data_142 <= trans_0_io_pipe_phv_out_data_142;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_143 <= init_io_pipe_phv_out_data_143; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_143 <= trans_1_io_pipe_phv_out_data_143;
    end else begin
      amplifier_0_0_data_143 <= trans_0_io_pipe_phv_out_data_143;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_144 <= init_io_pipe_phv_out_data_144; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_144 <= trans_1_io_pipe_phv_out_data_144;
    end else begin
      amplifier_0_0_data_144 <= trans_0_io_pipe_phv_out_data_144;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_145 <= init_io_pipe_phv_out_data_145; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_145 <= trans_1_io_pipe_phv_out_data_145;
    end else begin
      amplifier_0_0_data_145 <= trans_0_io_pipe_phv_out_data_145;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_146 <= init_io_pipe_phv_out_data_146; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_146 <= trans_1_io_pipe_phv_out_data_146;
    end else begin
      amplifier_0_0_data_146 <= trans_0_io_pipe_phv_out_data_146;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_147 <= init_io_pipe_phv_out_data_147; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_147 <= trans_1_io_pipe_phv_out_data_147;
    end else begin
      amplifier_0_0_data_147 <= trans_0_io_pipe_phv_out_data_147;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_148 <= init_io_pipe_phv_out_data_148; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_148 <= trans_1_io_pipe_phv_out_data_148;
    end else begin
      amplifier_0_0_data_148 <= trans_0_io_pipe_phv_out_data_148;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_149 <= init_io_pipe_phv_out_data_149; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_149 <= trans_1_io_pipe_phv_out_data_149;
    end else begin
      amplifier_0_0_data_149 <= trans_0_io_pipe_phv_out_data_149;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_150 <= init_io_pipe_phv_out_data_150; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_150 <= trans_1_io_pipe_phv_out_data_150;
    end else begin
      amplifier_0_0_data_150 <= trans_0_io_pipe_phv_out_data_150;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_151 <= init_io_pipe_phv_out_data_151; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_151 <= trans_1_io_pipe_phv_out_data_151;
    end else begin
      amplifier_0_0_data_151 <= trans_0_io_pipe_phv_out_data_151;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_152 <= init_io_pipe_phv_out_data_152; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_152 <= trans_1_io_pipe_phv_out_data_152;
    end else begin
      amplifier_0_0_data_152 <= trans_0_io_pipe_phv_out_data_152;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_153 <= init_io_pipe_phv_out_data_153; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_153 <= trans_1_io_pipe_phv_out_data_153;
    end else begin
      amplifier_0_0_data_153 <= trans_0_io_pipe_phv_out_data_153;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_154 <= init_io_pipe_phv_out_data_154; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_154 <= trans_1_io_pipe_phv_out_data_154;
    end else begin
      amplifier_0_0_data_154 <= trans_0_io_pipe_phv_out_data_154;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_155 <= init_io_pipe_phv_out_data_155; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_155 <= trans_1_io_pipe_phv_out_data_155;
    end else begin
      amplifier_0_0_data_155 <= trans_0_io_pipe_phv_out_data_155;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_156 <= init_io_pipe_phv_out_data_156; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_156 <= trans_1_io_pipe_phv_out_data_156;
    end else begin
      amplifier_0_0_data_156 <= trans_0_io_pipe_phv_out_data_156;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_157 <= init_io_pipe_phv_out_data_157; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_157 <= trans_1_io_pipe_phv_out_data_157;
    end else begin
      amplifier_0_0_data_157 <= trans_0_io_pipe_phv_out_data_157;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_158 <= init_io_pipe_phv_out_data_158; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_158 <= trans_1_io_pipe_phv_out_data_158;
    end else begin
      amplifier_0_0_data_158 <= trans_0_io_pipe_phv_out_data_158;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_159 <= init_io_pipe_phv_out_data_159; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_159 <= trans_1_io_pipe_phv_out_data_159;
    end else begin
      amplifier_0_0_data_159 <= trans_0_io_pipe_phv_out_data_159;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_160 <= init_io_pipe_phv_out_data_160; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_160 <= trans_1_io_pipe_phv_out_data_160;
    end else begin
      amplifier_0_0_data_160 <= trans_0_io_pipe_phv_out_data_160;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_161 <= init_io_pipe_phv_out_data_161; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_161 <= trans_1_io_pipe_phv_out_data_161;
    end else begin
      amplifier_0_0_data_161 <= trans_0_io_pipe_phv_out_data_161;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_162 <= init_io_pipe_phv_out_data_162; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_162 <= trans_1_io_pipe_phv_out_data_162;
    end else begin
      amplifier_0_0_data_162 <= trans_0_io_pipe_phv_out_data_162;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_163 <= init_io_pipe_phv_out_data_163; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_163 <= trans_1_io_pipe_phv_out_data_163;
    end else begin
      amplifier_0_0_data_163 <= trans_0_io_pipe_phv_out_data_163;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_164 <= init_io_pipe_phv_out_data_164; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_164 <= trans_1_io_pipe_phv_out_data_164;
    end else begin
      amplifier_0_0_data_164 <= trans_0_io_pipe_phv_out_data_164;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_165 <= init_io_pipe_phv_out_data_165; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_165 <= trans_1_io_pipe_phv_out_data_165;
    end else begin
      amplifier_0_0_data_165 <= trans_0_io_pipe_phv_out_data_165;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_166 <= init_io_pipe_phv_out_data_166; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_166 <= trans_1_io_pipe_phv_out_data_166;
    end else begin
      amplifier_0_0_data_166 <= trans_0_io_pipe_phv_out_data_166;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_167 <= init_io_pipe_phv_out_data_167; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_167 <= trans_1_io_pipe_phv_out_data_167;
    end else begin
      amplifier_0_0_data_167 <= trans_0_io_pipe_phv_out_data_167;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_168 <= init_io_pipe_phv_out_data_168; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_168 <= trans_1_io_pipe_phv_out_data_168;
    end else begin
      amplifier_0_0_data_168 <= trans_0_io_pipe_phv_out_data_168;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_169 <= init_io_pipe_phv_out_data_169; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_169 <= trans_1_io_pipe_phv_out_data_169;
    end else begin
      amplifier_0_0_data_169 <= trans_0_io_pipe_phv_out_data_169;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_170 <= init_io_pipe_phv_out_data_170; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_170 <= trans_1_io_pipe_phv_out_data_170;
    end else begin
      amplifier_0_0_data_170 <= trans_0_io_pipe_phv_out_data_170;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_171 <= init_io_pipe_phv_out_data_171; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_171 <= trans_1_io_pipe_phv_out_data_171;
    end else begin
      amplifier_0_0_data_171 <= trans_0_io_pipe_phv_out_data_171;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_172 <= init_io_pipe_phv_out_data_172; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_172 <= trans_1_io_pipe_phv_out_data_172;
    end else begin
      amplifier_0_0_data_172 <= trans_0_io_pipe_phv_out_data_172;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_173 <= init_io_pipe_phv_out_data_173; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_173 <= trans_1_io_pipe_phv_out_data_173;
    end else begin
      amplifier_0_0_data_173 <= trans_0_io_pipe_phv_out_data_173;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_174 <= init_io_pipe_phv_out_data_174; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_174 <= trans_1_io_pipe_phv_out_data_174;
    end else begin
      amplifier_0_0_data_174 <= trans_0_io_pipe_phv_out_data_174;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_175 <= init_io_pipe_phv_out_data_175; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_175 <= trans_1_io_pipe_phv_out_data_175;
    end else begin
      amplifier_0_0_data_175 <= trans_0_io_pipe_phv_out_data_175;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_176 <= init_io_pipe_phv_out_data_176; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_176 <= trans_1_io_pipe_phv_out_data_176;
    end else begin
      amplifier_0_0_data_176 <= trans_0_io_pipe_phv_out_data_176;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_177 <= init_io_pipe_phv_out_data_177; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_177 <= trans_1_io_pipe_phv_out_data_177;
    end else begin
      amplifier_0_0_data_177 <= trans_0_io_pipe_phv_out_data_177;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_178 <= init_io_pipe_phv_out_data_178; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_178 <= trans_1_io_pipe_phv_out_data_178;
    end else begin
      amplifier_0_0_data_178 <= trans_0_io_pipe_phv_out_data_178;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_179 <= init_io_pipe_phv_out_data_179; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_179 <= trans_1_io_pipe_phv_out_data_179;
    end else begin
      amplifier_0_0_data_179 <= trans_0_io_pipe_phv_out_data_179;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_180 <= init_io_pipe_phv_out_data_180; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_180 <= trans_1_io_pipe_phv_out_data_180;
    end else begin
      amplifier_0_0_data_180 <= trans_0_io_pipe_phv_out_data_180;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_181 <= init_io_pipe_phv_out_data_181; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_181 <= trans_1_io_pipe_phv_out_data_181;
    end else begin
      amplifier_0_0_data_181 <= trans_0_io_pipe_phv_out_data_181;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_182 <= init_io_pipe_phv_out_data_182; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_182 <= trans_1_io_pipe_phv_out_data_182;
    end else begin
      amplifier_0_0_data_182 <= trans_0_io_pipe_phv_out_data_182;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_183 <= init_io_pipe_phv_out_data_183; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_183 <= trans_1_io_pipe_phv_out_data_183;
    end else begin
      amplifier_0_0_data_183 <= trans_0_io_pipe_phv_out_data_183;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_184 <= init_io_pipe_phv_out_data_184; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_184 <= trans_1_io_pipe_phv_out_data_184;
    end else begin
      amplifier_0_0_data_184 <= trans_0_io_pipe_phv_out_data_184;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_185 <= init_io_pipe_phv_out_data_185; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_185 <= trans_1_io_pipe_phv_out_data_185;
    end else begin
      amplifier_0_0_data_185 <= trans_0_io_pipe_phv_out_data_185;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_186 <= init_io_pipe_phv_out_data_186; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_186 <= trans_1_io_pipe_phv_out_data_186;
    end else begin
      amplifier_0_0_data_186 <= trans_0_io_pipe_phv_out_data_186;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_187 <= init_io_pipe_phv_out_data_187; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_187 <= trans_1_io_pipe_phv_out_data_187;
    end else begin
      amplifier_0_0_data_187 <= trans_0_io_pipe_phv_out_data_187;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_188 <= init_io_pipe_phv_out_data_188; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_188 <= trans_1_io_pipe_phv_out_data_188;
    end else begin
      amplifier_0_0_data_188 <= trans_0_io_pipe_phv_out_data_188;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_189 <= init_io_pipe_phv_out_data_189; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_189 <= trans_1_io_pipe_phv_out_data_189;
    end else begin
      amplifier_0_0_data_189 <= trans_0_io_pipe_phv_out_data_189;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_190 <= init_io_pipe_phv_out_data_190; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_190 <= trans_1_io_pipe_phv_out_data_190;
    end else begin
      amplifier_0_0_data_190 <= trans_0_io_pipe_phv_out_data_190;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_191 <= init_io_pipe_phv_out_data_191; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_191 <= trans_1_io_pipe_phv_out_data_191;
    end else begin
      amplifier_0_0_data_191 <= trans_0_io_pipe_phv_out_data_191;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_192 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_192 <= trans_1_io_pipe_phv_out_data_192;
    end else begin
      amplifier_0_0_data_192 <= trans_0_io_pipe_phv_out_data_192;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_193 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_193 <= trans_1_io_pipe_phv_out_data_193;
    end else begin
      amplifier_0_0_data_193 <= trans_0_io_pipe_phv_out_data_193;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_194 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_194 <= trans_1_io_pipe_phv_out_data_194;
    end else begin
      amplifier_0_0_data_194 <= trans_0_io_pipe_phv_out_data_194;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_195 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_195 <= trans_1_io_pipe_phv_out_data_195;
    end else begin
      amplifier_0_0_data_195 <= trans_0_io_pipe_phv_out_data_195;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_196 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_196 <= trans_1_io_pipe_phv_out_data_196;
    end else begin
      amplifier_0_0_data_196 <= trans_0_io_pipe_phv_out_data_196;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_197 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_197 <= trans_1_io_pipe_phv_out_data_197;
    end else begin
      amplifier_0_0_data_197 <= trans_0_io_pipe_phv_out_data_197;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_198 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_198 <= trans_1_io_pipe_phv_out_data_198;
    end else begin
      amplifier_0_0_data_198 <= trans_0_io_pipe_phv_out_data_198;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_199 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_199 <= trans_1_io_pipe_phv_out_data_199;
    end else begin
      amplifier_0_0_data_199 <= trans_0_io_pipe_phv_out_data_199;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_200 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_200 <= trans_1_io_pipe_phv_out_data_200;
    end else begin
      amplifier_0_0_data_200 <= trans_0_io_pipe_phv_out_data_200;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_201 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_201 <= trans_1_io_pipe_phv_out_data_201;
    end else begin
      amplifier_0_0_data_201 <= trans_0_io_pipe_phv_out_data_201;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_202 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_202 <= trans_1_io_pipe_phv_out_data_202;
    end else begin
      amplifier_0_0_data_202 <= trans_0_io_pipe_phv_out_data_202;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_203 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_203 <= trans_1_io_pipe_phv_out_data_203;
    end else begin
      amplifier_0_0_data_203 <= trans_0_io_pipe_phv_out_data_203;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_204 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_204 <= trans_1_io_pipe_phv_out_data_204;
    end else begin
      amplifier_0_0_data_204 <= trans_0_io_pipe_phv_out_data_204;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_205 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_205 <= trans_1_io_pipe_phv_out_data_205;
    end else begin
      amplifier_0_0_data_205 <= trans_0_io_pipe_phv_out_data_205;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_206 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_206 <= trans_1_io_pipe_phv_out_data_206;
    end else begin
      amplifier_0_0_data_206 <= trans_0_io_pipe_phv_out_data_206;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_207 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_207 <= trans_1_io_pipe_phv_out_data_207;
    end else begin
      amplifier_0_0_data_207 <= trans_0_io_pipe_phv_out_data_207;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_208 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_208 <= trans_1_io_pipe_phv_out_data_208;
    end else begin
      amplifier_0_0_data_208 <= trans_0_io_pipe_phv_out_data_208;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_209 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_209 <= trans_1_io_pipe_phv_out_data_209;
    end else begin
      amplifier_0_0_data_209 <= trans_0_io_pipe_phv_out_data_209;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_210 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_210 <= trans_1_io_pipe_phv_out_data_210;
    end else begin
      amplifier_0_0_data_210 <= trans_0_io_pipe_phv_out_data_210;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_211 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_211 <= trans_1_io_pipe_phv_out_data_211;
    end else begin
      amplifier_0_0_data_211 <= trans_0_io_pipe_phv_out_data_211;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_212 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_212 <= trans_1_io_pipe_phv_out_data_212;
    end else begin
      amplifier_0_0_data_212 <= trans_0_io_pipe_phv_out_data_212;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_213 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_213 <= trans_1_io_pipe_phv_out_data_213;
    end else begin
      amplifier_0_0_data_213 <= trans_0_io_pipe_phv_out_data_213;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_214 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_214 <= trans_1_io_pipe_phv_out_data_214;
    end else begin
      amplifier_0_0_data_214 <= trans_0_io_pipe_phv_out_data_214;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_215 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_215 <= trans_1_io_pipe_phv_out_data_215;
    end else begin
      amplifier_0_0_data_215 <= trans_0_io_pipe_phv_out_data_215;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_216 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_216 <= trans_1_io_pipe_phv_out_data_216;
    end else begin
      amplifier_0_0_data_216 <= trans_0_io_pipe_phv_out_data_216;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_217 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_217 <= trans_1_io_pipe_phv_out_data_217;
    end else begin
      amplifier_0_0_data_217 <= trans_0_io_pipe_phv_out_data_217;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_218 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_218 <= trans_1_io_pipe_phv_out_data_218;
    end else begin
      amplifier_0_0_data_218 <= trans_0_io_pipe_phv_out_data_218;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_219 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_219 <= trans_1_io_pipe_phv_out_data_219;
    end else begin
      amplifier_0_0_data_219 <= trans_0_io_pipe_phv_out_data_219;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_220 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_220 <= trans_1_io_pipe_phv_out_data_220;
    end else begin
      amplifier_0_0_data_220 <= trans_0_io_pipe_phv_out_data_220;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_221 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_221 <= trans_1_io_pipe_phv_out_data_221;
    end else begin
      amplifier_0_0_data_221 <= trans_0_io_pipe_phv_out_data_221;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_222 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_222 <= trans_1_io_pipe_phv_out_data_222;
    end else begin
      amplifier_0_0_data_222 <= trans_0_io_pipe_phv_out_data_222;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_223 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_223 <= trans_1_io_pipe_phv_out_data_223;
    end else begin
      amplifier_0_0_data_223 <= trans_0_io_pipe_phv_out_data_223;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_224 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_224 <= trans_1_io_pipe_phv_out_data_224;
    end else begin
      amplifier_0_0_data_224 <= trans_0_io_pipe_phv_out_data_224;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_225 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_225 <= trans_1_io_pipe_phv_out_data_225;
    end else begin
      amplifier_0_0_data_225 <= trans_0_io_pipe_phv_out_data_225;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_226 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_226 <= trans_1_io_pipe_phv_out_data_226;
    end else begin
      amplifier_0_0_data_226 <= trans_0_io_pipe_phv_out_data_226;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_227 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_227 <= trans_1_io_pipe_phv_out_data_227;
    end else begin
      amplifier_0_0_data_227 <= trans_0_io_pipe_phv_out_data_227;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_228 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_228 <= trans_1_io_pipe_phv_out_data_228;
    end else begin
      amplifier_0_0_data_228 <= trans_0_io_pipe_phv_out_data_228;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_229 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_229 <= trans_1_io_pipe_phv_out_data_229;
    end else begin
      amplifier_0_0_data_229 <= trans_0_io_pipe_phv_out_data_229;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_230 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_230 <= trans_1_io_pipe_phv_out_data_230;
    end else begin
      amplifier_0_0_data_230 <= trans_0_io_pipe_phv_out_data_230;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_231 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_231 <= trans_1_io_pipe_phv_out_data_231;
    end else begin
      amplifier_0_0_data_231 <= trans_0_io_pipe_phv_out_data_231;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_232 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_232 <= trans_1_io_pipe_phv_out_data_232;
    end else begin
      amplifier_0_0_data_232 <= trans_0_io_pipe_phv_out_data_232;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_233 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_233 <= trans_1_io_pipe_phv_out_data_233;
    end else begin
      amplifier_0_0_data_233 <= trans_0_io_pipe_phv_out_data_233;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_234 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_234 <= trans_1_io_pipe_phv_out_data_234;
    end else begin
      amplifier_0_0_data_234 <= trans_0_io_pipe_phv_out_data_234;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_235 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_235 <= trans_1_io_pipe_phv_out_data_235;
    end else begin
      amplifier_0_0_data_235 <= trans_0_io_pipe_phv_out_data_235;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_236 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_236 <= trans_1_io_pipe_phv_out_data_236;
    end else begin
      amplifier_0_0_data_236 <= trans_0_io_pipe_phv_out_data_236;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_237 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_237 <= trans_1_io_pipe_phv_out_data_237;
    end else begin
      amplifier_0_0_data_237 <= trans_0_io_pipe_phv_out_data_237;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_238 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_238 <= trans_1_io_pipe_phv_out_data_238;
    end else begin
      amplifier_0_0_data_238 <= trans_0_io_pipe_phv_out_data_238;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_239 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_239 <= trans_1_io_pipe_phv_out_data_239;
    end else begin
      amplifier_0_0_data_239 <= trans_0_io_pipe_phv_out_data_239;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_240 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_240 <= trans_1_io_pipe_phv_out_data_240;
    end else begin
      amplifier_0_0_data_240 <= trans_0_io_pipe_phv_out_data_240;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_241 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_241 <= trans_1_io_pipe_phv_out_data_241;
    end else begin
      amplifier_0_0_data_241 <= trans_0_io_pipe_phv_out_data_241;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_242 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_242 <= trans_1_io_pipe_phv_out_data_242;
    end else begin
      amplifier_0_0_data_242 <= trans_0_io_pipe_phv_out_data_242;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_243 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_243 <= trans_1_io_pipe_phv_out_data_243;
    end else begin
      amplifier_0_0_data_243 <= trans_0_io_pipe_phv_out_data_243;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_244 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_244 <= trans_1_io_pipe_phv_out_data_244;
    end else begin
      amplifier_0_0_data_244 <= trans_0_io_pipe_phv_out_data_244;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_245 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_245 <= trans_1_io_pipe_phv_out_data_245;
    end else begin
      amplifier_0_0_data_245 <= trans_0_io_pipe_phv_out_data_245;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_246 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_246 <= trans_1_io_pipe_phv_out_data_246;
    end else begin
      amplifier_0_0_data_246 <= trans_0_io_pipe_phv_out_data_246;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_247 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_247 <= trans_1_io_pipe_phv_out_data_247;
    end else begin
      amplifier_0_0_data_247 <= trans_0_io_pipe_phv_out_data_247;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_248 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_248 <= trans_1_io_pipe_phv_out_data_248;
    end else begin
      amplifier_0_0_data_248 <= trans_0_io_pipe_phv_out_data_248;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_249 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_249 <= trans_1_io_pipe_phv_out_data_249;
    end else begin
      amplifier_0_0_data_249 <= trans_0_io_pipe_phv_out_data_249;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_250 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_250 <= trans_1_io_pipe_phv_out_data_250;
    end else begin
      amplifier_0_0_data_250 <= trans_0_io_pipe_phv_out_data_250;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_251 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_251 <= trans_1_io_pipe_phv_out_data_251;
    end else begin
      amplifier_0_0_data_251 <= trans_0_io_pipe_phv_out_data_251;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_252 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_252 <= trans_1_io_pipe_phv_out_data_252;
    end else begin
      amplifier_0_0_data_252 <= trans_0_io_pipe_phv_out_data_252;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_253 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_253 <= trans_1_io_pipe_phv_out_data_253;
    end else begin
      amplifier_0_0_data_253 <= trans_0_io_pipe_phv_out_data_253;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_254 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_254 <= trans_1_io_pipe_phv_out_data_254;
    end else begin
      amplifier_0_0_data_254 <= trans_0_io_pipe_phv_out_data_254;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_data_255 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_data_255 <= trans_1_io_pipe_phv_out_data_255;
    end else begin
      amplifier_0_0_data_255 <= trans_0_io_pipe_phv_out_data_255;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_header_0 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_header_0 <= trans_1_io_pipe_phv_out_header_0;
    end else begin
      amplifier_0_0_header_0 <= trans_0_io_pipe_phv_out_header_0;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_header_1 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_header_1 <= trans_1_io_pipe_phv_out_header_1;
    end else begin
      amplifier_0_0_header_1 <= trans_0_io_pipe_phv_out_header_1;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_header_2 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_header_2 <= trans_1_io_pipe_phv_out_header_2;
    end else begin
      amplifier_0_0_header_2 <= trans_0_io_pipe_phv_out_header_2;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_header_3 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_header_3 <= trans_1_io_pipe_phv_out_header_3;
    end else begin
      amplifier_0_0_header_3 <= trans_0_io_pipe_phv_out_header_3;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_header_4 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_header_4 <= trans_1_io_pipe_phv_out_header_4;
    end else begin
      amplifier_0_0_header_4 <= trans_0_io_pipe_phv_out_header_4;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_header_5 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_header_5 <= trans_1_io_pipe_phv_out_header_5;
    end else begin
      amplifier_0_0_header_5 <= trans_0_io_pipe_phv_out_header_5;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_header_6 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_header_6 <= trans_1_io_pipe_phv_out_header_6;
    end else begin
      amplifier_0_0_header_6 <= trans_0_io_pipe_phv_out_header_6;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_header_7 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_header_7 <= trans_1_io_pipe_phv_out_header_7;
    end else begin
      amplifier_0_0_header_7 <= trans_0_io_pipe_phv_out_header_7;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_header_8 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_header_8 <= trans_1_io_pipe_phv_out_header_8;
    end else begin
      amplifier_0_0_header_8 <= trans_0_io_pipe_phv_out_header_8;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_header_9 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_header_9 <= trans_1_io_pipe_phv_out_header_9;
    end else begin
      amplifier_0_0_header_9 <= trans_0_io_pipe_phv_out_header_9;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_header_10 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_header_10 <= trans_1_io_pipe_phv_out_header_10;
    end else begin
      amplifier_0_0_header_10 <= trans_0_io_pipe_phv_out_header_10;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_header_11 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_header_11 <= trans_1_io_pipe_phv_out_header_11;
    end else begin
      amplifier_0_0_header_11 <= trans_0_io_pipe_phv_out_header_11;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_header_12 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_header_12 <= trans_1_io_pipe_phv_out_header_12;
    end else begin
      amplifier_0_0_header_12 <= trans_0_io_pipe_phv_out_header_12;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_header_13 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_header_13 <= trans_1_io_pipe_phv_out_header_13;
    end else begin
      amplifier_0_0_header_13 <= trans_0_io_pipe_phv_out_header_13;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_header_14 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_header_14 <= trans_1_io_pipe_phv_out_header_14;
    end else begin
      amplifier_0_0_header_14 <= trans_0_io_pipe_phv_out_header_14;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_header_15 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_header_15 <= trans_1_io_pipe_phv_out_header_15;
    end else begin
      amplifier_0_0_header_15 <= trans_0_io_pipe_phv_out_header_15;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_parse_current_state <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_parse_current_state <= trans_1_io_pipe_phv_out_parse_current_state;
    end else begin
      amplifier_0_0_parse_current_state <= trans_0_io_pipe_phv_out_parse_current_state;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_parse_current_offset <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_parse_current_offset <= trans_1_io_pipe_phv_out_parse_current_offset;
    end else begin
      amplifier_0_0_parse_current_offset <= trans_0_io_pipe_phv_out_parse_current_offset;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_parse_transition_field <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_parse_transition_field <= trans_1_io_pipe_phv_out_parse_transition_field;
    end else begin
      amplifier_0_0_parse_transition_field <= trans_0_io_pipe_phv_out_parse_transition_field;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_next_processor_id <= init_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_next_processor_id <= trans_1_io_pipe_phv_out_next_processor_id;
    end else begin
      amplifier_0_0_next_processor_id <= trans_0_io_pipe_phv_out_next_processor_id;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_next_config_id <= 1'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_next_config_id <= trans_1_io_pipe_phv_out_next_config_id;
    end else begin
      amplifier_0_0_next_config_id <= trans_0_io_pipe_phv_out_next_config_id;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      amplifier_0_0_is_valid_processor <= 1'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 109:31]
      amplifier_0_0_is_valid_processor <= trans_1_io_pipe_phv_out_is_valid_processor;
    end else begin
      amplifier_0_0_is_valid_processor <= trans_0_io_pipe_phv_out_is_valid_processor;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_0 <= init_io_pipe_phv_out_data_0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_0 <= trans_0_io_pipe_phv_out_data_0;
    end else begin
      amplifier_0_1_data_0 <= trans_1_io_pipe_phv_out_data_0;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_1 <= init_io_pipe_phv_out_data_1; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_1 <= trans_0_io_pipe_phv_out_data_1;
    end else begin
      amplifier_0_1_data_1 <= trans_1_io_pipe_phv_out_data_1;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_2 <= init_io_pipe_phv_out_data_2; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_2 <= trans_0_io_pipe_phv_out_data_2;
    end else begin
      amplifier_0_1_data_2 <= trans_1_io_pipe_phv_out_data_2;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_3 <= init_io_pipe_phv_out_data_3; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_3 <= trans_0_io_pipe_phv_out_data_3;
    end else begin
      amplifier_0_1_data_3 <= trans_1_io_pipe_phv_out_data_3;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_4 <= init_io_pipe_phv_out_data_4; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_4 <= trans_0_io_pipe_phv_out_data_4;
    end else begin
      amplifier_0_1_data_4 <= trans_1_io_pipe_phv_out_data_4;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_5 <= init_io_pipe_phv_out_data_5; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_5 <= trans_0_io_pipe_phv_out_data_5;
    end else begin
      amplifier_0_1_data_5 <= trans_1_io_pipe_phv_out_data_5;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_6 <= init_io_pipe_phv_out_data_6; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_6 <= trans_0_io_pipe_phv_out_data_6;
    end else begin
      amplifier_0_1_data_6 <= trans_1_io_pipe_phv_out_data_6;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_7 <= init_io_pipe_phv_out_data_7; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_7 <= trans_0_io_pipe_phv_out_data_7;
    end else begin
      amplifier_0_1_data_7 <= trans_1_io_pipe_phv_out_data_7;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_8 <= init_io_pipe_phv_out_data_8; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_8 <= trans_0_io_pipe_phv_out_data_8;
    end else begin
      amplifier_0_1_data_8 <= trans_1_io_pipe_phv_out_data_8;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_9 <= init_io_pipe_phv_out_data_9; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_9 <= trans_0_io_pipe_phv_out_data_9;
    end else begin
      amplifier_0_1_data_9 <= trans_1_io_pipe_phv_out_data_9;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_10 <= init_io_pipe_phv_out_data_10; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_10 <= trans_0_io_pipe_phv_out_data_10;
    end else begin
      amplifier_0_1_data_10 <= trans_1_io_pipe_phv_out_data_10;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_11 <= init_io_pipe_phv_out_data_11; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_11 <= trans_0_io_pipe_phv_out_data_11;
    end else begin
      amplifier_0_1_data_11 <= trans_1_io_pipe_phv_out_data_11;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_12 <= init_io_pipe_phv_out_data_12; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_12 <= trans_0_io_pipe_phv_out_data_12;
    end else begin
      amplifier_0_1_data_12 <= trans_1_io_pipe_phv_out_data_12;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_13 <= init_io_pipe_phv_out_data_13; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_13 <= trans_0_io_pipe_phv_out_data_13;
    end else begin
      amplifier_0_1_data_13 <= trans_1_io_pipe_phv_out_data_13;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_14 <= init_io_pipe_phv_out_data_14; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_14 <= trans_0_io_pipe_phv_out_data_14;
    end else begin
      amplifier_0_1_data_14 <= trans_1_io_pipe_phv_out_data_14;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_15 <= init_io_pipe_phv_out_data_15; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_15 <= trans_0_io_pipe_phv_out_data_15;
    end else begin
      amplifier_0_1_data_15 <= trans_1_io_pipe_phv_out_data_15;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_16 <= init_io_pipe_phv_out_data_16; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_16 <= trans_0_io_pipe_phv_out_data_16;
    end else begin
      amplifier_0_1_data_16 <= trans_1_io_pipe_phv_out_data_16;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_17 <= init_io_pipe_phv_out_data_17; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_17 <= trans_0_io_pipe_phv_out_data_17;
    end else begin
      amplifier_0_1_data_17 <= trans_1_io_pipe_phv_out_data_17;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_18 <= init_io_pipe_phv_out_data_18; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_18 <= trans_0_io_pipe_phv_out_data_18;
    end else begin
      amplifier_0_1_data_18 <= trans_1_io_pipe_phv_out_data_18;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_19 <= init_io_pipe_phv_out_data_19; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_19 <= trans_0_io_pipe_phv_out_data_19;
    end else begin
      amplifier_0_1_data_19 <= trans_1_io_pipe_phv_out_data_19;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_20 <= init_io_pipe_phv_out_data_20; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_20 <= trans_0_io_pipe_phv_out_data_20;
    end else begin
      amplifier_0_1_data_20 <= trans_1_io_pipe_phv_out_data_20;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_21 <= init_io_pipe_phv_out_data_21; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_21 <= trans_0_io_pipe_phv_out_data_21;
    end else begin
      amplifier_0_1_data_21 <= trans_1_io_pipe_phv_out_data_21;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_22 <= init_io_pipe_phv_out_data_22; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_22 <= trans_0_io_pipe_phv_out_data_22;
    end else begin
      amplifier_0_1_data_22 <= trans_1_io_pipe_phv_out_data_22;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_23 <= init_io_pipe_phv_out_data_23; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_23 <= trans_0_io_pipe_phv_out_data_23;
    end else begin
      amplifier_0_1_data_23 <= trans_1_io_pipe_phv_out_data_23;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_24 <= init_io_pipe_phv_out_data_24; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_24 <= trans_0_io_pipe_phv_out_data_24;
    end else begin
      amplifier_0_1_data_24 <= trans_1_io_pipe_phv_out_data_24;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_25 <= init_io_pipe_phv_out_data_25; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_25 <= trans_0_io_pipe_phv_out_data_25;
    end else begin
      amplifier_0_1_data_25 <= trans_1_io_pipe_phv_out_data_25;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_26 <= init_io_pipe_phv_out_data_26; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_26 <= trans_0_io_pipe_phv_out_data_26;
    end else begin
      amplifier_0_1_data_26 <= trans_1_io_pipe_phv_out_data_26;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_27 <= init_io_pipe_phv_out_data_27; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_27 <= trans_0_io_pipe_phv_out_data_27;
    end else begin
      amplifier_0_1_data_27 <= trans_1_io_pipe_phv_out_data_27;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_28 <= init_io_pipe_phv_out_data_28; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_28 <= trans_0_io_pipe_phv_out_data_28;
    end else begin
      amplifier_0_1_data_28 <= trans_1_io_pipe_phv_out_data_28;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_29 <= init_io_pipe_phv_out_data_29; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_29 <= trans_0_io_pipe_phv_out_data_29;
    end else begin
      amplifier_0_1_data_29 <= trans_1_io_pipe_phv_out_data_29;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_30 <= init_io_pipe_phv_out_data_30; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_30 <= trans_0_io_pipe_phv_out_data_30;
    end else begin
      amplifier_0_1_data_30 <= trans_1_io_pipe_phv_out_data_30;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_31 <= init_io_pipe_phv_out_data_31; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_31 <= trans_0_io_pipe_phv_out_data_31;
    end else begin
      amplifier_0_1_data_31 <= trans_1_io_pipe_phv_out_data_31;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_32 <= init_io_pipe_phv_out_data_32; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_32 <= trans_0_io_pipe_phv_out_data_32;
    end else begin
      amplifier_0_1_data_32 <= trans_1_io_pipe_phv_out_data_32;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_33 <= init_io_pipe_phv_out_data_33; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_33 <= trans_0_io_pipe_phv_out_data_33;
    end else begin
      amplifier_0_1_data_33 <= trans_1_io_pipe_phv_out_data_33;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_34 <= init_io_pipe_phv_out_data_34; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_34 <= trans_0_io_pipe_phv_out_data_34;
    end else begin
      amplifier_0_1_data_34 <= trans_1_io_pipe_phv_out_data_34;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_35 <= init_io_pipe_phv_out_data_35; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_35 <= trans_0_io_pipe_phv_out_data_35;
    end else begin
      amplifier_0_1_data_35 <= trans_1_io_pipe_phv_out_data_35;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_36 <= init_io_pipe_phv_out_data_36; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_36 <= trans_0_io_pipe_phv_out_data_36;
    end else begin
      amplifier_0_1_data_36 <= trans_1_io_pipe_phv_out_data_36;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_37 <= init_io_pipe_phv_out_data_37; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_37 <= trans_0_io_pipe_phv_out_data_37;
    end else begin
      amplifier_0_1_data_37 <= trans_1_io_pipe_phv_out_data_37;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_38 <= init_io_pipe_phv_out_data_38; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_38 <= trans_0_io_pipe_phv_out_data_38;
    end else begin
      amplifier_0_1_data_38 <= trans_1_io_pipe_phv_out_data_38;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_39 <= init_io_pipe_phv_out_data_39; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_39 <= trans_0_io_pipe_phv_out_data_39;
    end else begin
      amplifier_0_1_data_39 <= trans_1_io_pipe_phv_out_data_39;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_40 <= init_io_pipe_phv_out_data_40; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_40 <= trans_0_io_pipe_phv_out_data_40;
    end else begin
      amplifier_0_1_data_40 <= trans_1_io_pipe_phv_out_data_40;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_41 <= init_io_pipe_phv_out_data_41; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_41 <= trans_0_io_pipe_phv_out_data_41;
    end else begin
      amplifier_0_1_data_41 <= trans_1_io_pipe_phv_out_data_41;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_42 <= init_io_pipe_phv_out_data_42; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_42 <= trans_0_io_pipe_phv_out_data_42;
    end else begin
      amplifier_0_1_data_42 <= trans_1_io_pipe_phv_out_data_42;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_43 <= init_io_pipe_phv_out_data_43; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_43 <= trans_0_io_pipe_phv_out_data_43;
    end else begin
      amplifier_0_1_data_43 <= trans_1_io_pipe_phv_out_data_43;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_44 <= init_io_pipe_phv_out_data_44; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_44 <= trans_0_io_pipe_phv_out_data_44;
    end else begin
      amplifier_0_1_data_44 <= trans_1_io_pipe_phv_out_data_44;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_45 <= init_io_pipe_phv_out_data_45; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_45 <= trans_0_io_pipe_phv_out_data_45;
    end else begin
      amplifier_0_1_data_45 <= trans_1_io_pipe_phv_out_data_45;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_46 <= init_io_pipe_phv_out_data_46; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_46 <= trans_0_io_pipe_phv_out_data_46;
    end else begin
      amplifier_0_1_data_46 <= trans_1_io_pipe_phv_out_data_46;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_47 <= init_io_pipe_phv_out_data_47; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_47 <= trans_0_io_pipe_phv_out_data_47;
    end else begin
      amplifier_0_1_data_47 <= trans_1_io_pipe_phv_out_data_47;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_48 <= init_io_pipe_phv_out_data_48; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_48 <= trans_0_io_pipe_phv_out_data_48;
    end else begin
      amplifier_0_1_data_48 <= trans_1_io_pipe_phv_out_data_48;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_49 <= init_io_pipe_phv_out_data_49; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_49 <= trans_0_io_pipe_phv_out_data_49;
    end else begin
      amplifier_0_1_data_49 <= trans_1_io_pipe_phv_out_data_49;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_50 <= init_io_pipe_phv_out_data_50; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_50 <= trans_0_io_pipe_phv_out_data_50;
    end else begin
      amplifier_0_1_data_50 <= trans_1_io_pipe_phv_out_data_50;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_51 <= init_io_pipe_phv_out_data_51; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_51 <= trans_0_io_pipe_phv_out_data_51;
    end else begin
      amplifier_0_1_data_51 <= trans_1_io_pipe_phv_out_data_51;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_52 <= init_io_pipe_phv_out_data_52; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_52 <= trans_0_io_pipe_phv_out_data_52;
    end else begin
      amplifier_0_1_data_52 <= trans_1_io_pipe_phv_out_data_52;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_53 <= init_io_pipe_phv_out_data_53; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_53 <= trans_0_io_pipe_phv_out_data_53;
    end else begin
      amplifier_0_1_data_53 <= trans_1_io_pipe_phv_out_data_53;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_54 <= init_io_pipe_phv_out_data_54; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_54 <= trans_0_io_pipe_phv_out_data_54;
    end else begin
      amplifier_0_1_data_54 <= trans_1_io_pipe_phv_out_data_54;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_55 <= init_io_pipe_phv_out_data_55; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_55 <= trans_0_io_pipe_phv_out_data_55;
    end else begin
      amplifier_0_1_data_55 <= trans_1_io_pipe_phv_out_data_55;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_56 <= init_io_pipe_phv_out_data_56; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_56 <= trans_0_io_pipe_phv_out_data_56;
    end else begin
      amplifier_0_1_data_56 <= trans_1_io_pipe_phv_out_data_56;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_57 <= init_io_pipe_phv_out_data_57; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_57 <= trans_0_io_pipe_phv_out_data_57;
    end else begin
      amplifier_0_1_data_57 <= trans_1_io_pipe_phv_out_data_57;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_58 <= init_io_pipe_phv_out_data_58; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_58 <= trans_0_io_pipe_phv_out_data_58;
    end else begin
      amplifier_0_1_data_58 <= trans_1_io_pipe_phv_out_data_58;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_59 <= init_io_pipe_phv_out_data_59; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_59 <= trans_0_io_pipe_phv_out_data_59;
    end else begin
      amplifier_0_1_data_59 <= trans_1_io_pipe_phv_out_data_59;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_60 <= init_io_pipe_phv_out_data_60; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_60 <= trans_0_io_pipe_phv_out_data_60;
    end else begin
      amplifier_0_1_data_60 <= trans_1_io_pipe_phv_out_data_60;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_61 <= init_io_pipe_phv_out_data_61; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_61 <= trans_0_io_pipe_phv_out_data_61;
    end else begin
      amplifier_0_1_data_61 <= trans_1_io_pipe_phv_out_data_61;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_62 <= init_io_pipe_phv_out_data_62; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_62 <= trans_0_io_pipe_phv_out_data_62;
    end else begin
      amplifier_0_1_data_62 <= trans_1_io_pipe_phv_out_data_62;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_63 <= init_io_pipe_phv_out_data_63; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_63 <= trans_0_io_pipe_phv_out_data_63;
    end else begin
      amplifier_0_1_data_63 <= trans_1_io_pipe_phv_out_data_63;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_64 <= init_io_pipe_phv_out_data_64; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_64 <= trans_0_io_pipe_phv_out_data_64;
    end else begin
      amplifier_0_1_data_64 <= trans_1_io_pipe_phv_out_data_64;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_65 <= init_io_pipe_phv_out_data_65; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_65 <= trans_0_io_pipe_phv_out_data_65;
    end else begin
      amplifier_0_1_data_65 <= trans_1_io_pipe_phv_out_data_65;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_66 <= init_io_pipe_phv_out_data_66; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_66 <= trans_0_io_pipe_phv_out_data_66;
    end else begin
      amplifier_0_1_data_66 <= trans_1_io_pipe_phv_out_data_66;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_67 <= init_io_pipe_phv_out_data_67; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_67 <= trans_0_io_pipe_phv_out_data_67;
    end else begin
      amplifier_0_1_data_67 <= trans_1_io_pipe_phv_out_data_67;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_68 <= init_io_pipe_phv_out_data_68; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_68 <= trans_0_io_pipe_phv_out_data_68;
    end else begin
      amplifier_0_1_data_68 <= trans_1_io_pipe_phv_out_data_68;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_69 <= init_io_pipe_phv_out_data_69; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_69 <= trans_0_io_pipe_phv_out_data_69;
    end else begin
      amplifier_0_1_data_69 <= trans_1_io_pipe_phv_out_data_69;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_70 <= init_io_pipe_phv_out_data_70; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_70 <= trans_0_io_pipe_phv_out_data_70;
    end else begin
      amplifier_0_1_data_70 <= trans_1_io_pipe_phv_out_data_70;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_71 <= init_io_pipe_phv_out_data_71; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_71 <= trans_0_io_pipe_phv_out_data_71;
    end else begin
      amplifier_0_1_data_71 <= trans_1_io_pipe_phv_out_data_71;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_72 <= init_io_pipe_phv_out_data_72; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_72 <= trans_0_io_pipe_phv_out_data_72;
    end else begin
      amplifier_0_1_data_72 <= trans_1_io_pipe_phv_out_data_72;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_73 <= init_io_pipe_phv_out_data_73; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_73 <= trans_0_io_pipe_phv_out_data_73;
    end else begin
      amplifier_0_1_data_73 <= trans_1_io_pipe_phv_out_data_73;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_74 <= init_io_pipe_phv_out_data_74; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_74 <= trans_0_io_pipe_phv_out_data_74;
    end else begin
      amplifier_0_1_data_74 <= trans_1_io_pipe_phv_out_data_74;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_75 <= init_io_pipe_phv_out_data_75; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_75 <= trans_0_io_pipe_phv_out_data_75;
    end else begin
      amplifier_0_1_data_75 <= trans_1_io_pipe_phv_out_data_75;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_76 <= init_io_pipe_phv_out_data_76; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_76 <= trans_0_io_pipe_phv_out_data_76;
    end else begin
      amplifier_0_1_data_76 <= trans_1_io_pipe_phv_out_data_76;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_77 <= init_io_pipe_phv_out_data_77; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_77 <= trans_0_io_pipe_phv_out_data_77;
    end else begin
      amplifier_0_1_data_77 <= trans_1_io_pipe_phv_out_data_77;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_78 <= init_io_pipe_phv_out_data_78; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_78 <= trans_0_io_pipe_phv_out_data_78;
    end else begin
      amplifier_0_1_data_78 <= trans_1_io_pipe_phv_out_data_78;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_79 <= init_io_pipe_phv_out_data_79; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_79 <= trans_0_io_pipe_phv_out_data_79;
    end else begin
      amplifier_0_1_data_79 <= trans_1_io_pipe_phv_out_data_79;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_80 <= init_io_pipe_phv_out_data_80; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_80 <= trans_0_io_pipe_phv_out_data_80;
    end else begin
      amplifier_0_1_data_80 <= trans_1_io_pipe_phv_out_data_80;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_81 <= init_io_pipe_phv_out_data_81; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_81 <= trans_0_io_pipe_phv_out_data_81;
    end else begin
      amplifier_0_1_data_81 <= trans_1_io_pipe_phv_out_data_81;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_82 <= init_io_pipe_phv_out_data_82; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_82 <= trans_0_io_pipe_phv_out_data_82;
    end else begin
      amplifier_0_1_data_82 <= trans_1_io_pipe_phv_out_data_82;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_83 <= init_io_pipe_phv_out_data_83; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_83 <= trans_0_io_pipe_phv_out_data_83;
    end else begin
      amplifier_0_1_data_83 <= trans_1_io_pipe_phv_out_data_83;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_84 <= init_io_pipe_phv_out_data_84; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_84 <= trans_0_io_pipe_phv_out_data_84;
    end else begin
      amplifier_0_1_data_84 <= trans_1_io_pipe_phv_out_data_84;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_85 <= init_io_pipe_phv_out_data_85; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_85 <= trans_0_io_pipe_phv_out_data_85;
    end else begin
      amplifier_0_1_data_85 <= trans_1_io_pipe_phv_out_data_85;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_86 <= init_io_pipe_phv_out_data_86; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_86 <= trans_0_io_pipe_phv_out_data_86;
    end else begin
      amplifier_0_1_data_86 <= trans_1_io_pipe_phv_out_data_86;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_87 <= init_io_pipe_phv_out_data_87; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_87 <= trans_0_io_pipe_phv_out_data_87;
    end else begin
      amplifier_0_1_data_87 <= trans_1_io_pipe_phv_out_data_87;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_88 <= init_io_pipe_phv_out_data_88; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_88 <= trans_0_io_pipe_phv_out_data_88;
    end else begin
      amplifier_0_1_data_88 <= trans_1_io_pipe_phv_out_data_88;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_89 <= init_io_pipe_phv_out_data_89; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_89 <= trans_0_io_pipe_phv_out_data_89;
    end else begin
      amplifier_0_1_data_89 <= trans_1_io_pipe_phv_out_data_89;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_90 <= init_io_pipe_phv_out_data_90; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_90 <= trans_0_io_pipe_phv_out_data_90;
    end else begin
      amplifier_0_1_data_90 <= trans_1_io_pipe_phv_out_data_90;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_91 <= init_io_pipe_phv_out_data_91; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_91 <= trans_0_io_pipe_phv_out_data_91;
    end else begin
      amplifier_0_1_data_91 <= trans_1_io_pipe_phv_out_data_91;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_92 <= init_io_pipe_phv_out_data_92; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_92 <= trans_0_io_pipe_phv_out_data_92;
    end else begin
      amplifier_0_1_data_92 <= trans_1_io_pipe_phv_out_data_92;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_93 <= init_io_pipe_phv_out_data_93; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_93 <= trans_0_io_pipe_phv_out_data_93;
    end else begin
      amplifier_0_1_data_93 <= trans_1_io_pipe_phv_out_data_93;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_94 <= init_io_pipe_phv_out_data_94; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_94 <= trans_0_io_pipe_phv_out_data_94;
    end else begin
      amplifier_0_1_data_94 <= trans_1_io_pipe_phv_out_data_94;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_95 <= init_io_pipe_phv_out_data_95; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_95 <= trans_0_io_pipe_phv_out_data_95;
    end else begin
      amplifier_0_1_data_95 <= trans_1_io_pipe_phv_out_data_95;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_96 <= init_io_pipe_phv_out_data_96; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_96 <= trans_0_io_pipe_phv_out_data_96;
    end else begin
      amplifier_0_1_data_96 <= trans_1_io_pipe_phv_out_data_96;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_97 <= init_io_pipe_phv_out_data_97; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_97 <= trans_0_io_pipe_phv_out_data_97;
    end else begin
      amplifier_0_1_data_97 <= trans_1_io_pipe_phv_out_data_97;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_98 <= init_io_pipe_phv_out_data_98; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_98 <= trans_0_io_pipe_phv_out_data_98;
    end else begin
      amplifier_0_1_data_98 <= trans_1_io_pipe_phv_out_data_98;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_99 <= init_io_pipe_phv_out_data_99; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_99 <= trans_0_io_pipe_phv_out_data_99;
    end else begin
      amplifier_0_1_data_99 <= trans_1_io_pipe_phv_out_data_99;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_100 <= init_io_pipe_phv_out_data_100; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_100 <= trans_0_io_pipe_phv_out_data_100;
    end else begin
      amplifier_0_1_data_100 <= trans_1_io_pipe_phv_out_data_100;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_101 <= init_io_pipe_phv_out_data_101; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_101 <= trans_0_io_pipe_phv_out_data_101;
    end else begin
      amplifier_0_1_data_101 <= trans_1_io_pipe_phv_out_data_101;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_102 <= init_io_pipe_phv_out_data_102; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_102 <= trans_0_io_pipe_phv_out_data_102;
    end else begin
      amplifier_0_1_data_102 <= trans_1_io_pipe_phv_out_data_102;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_103 <= init_io_pipe_phv_out_data_103; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_103 <= trans_0_io_pipe_phv_out_data_103;
    end else begin
      amplifier_0_1_data_103 <= trans_1_io_pipe_phv_out_data_103;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_104 <= init_io_pipe_phv_out_data_104; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_104 <= trans_0_io_pipe_phv_out_data_104;
    end else begin
      amplifier_0_1_data_104 <= trans_1_io_pipe_phv_out_data_104;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_105 <= init_io_pipe_phv_out_data_105; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_105 <= trans_0_io_pipe_phv_out_data_105;
    end else begin
      amplifier_0_1_data_105 <= trans_1_io_pipe_phv_out_data_105;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_106 <= init_io_pipe_phv_out_data_106; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_106 <= trans_0_io_pipe_phv_out_data_106;
    end else begin
      amplifier_0_1_data_106 <= trans_1_io_pipe_phv_out_data_106;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_107 <= init_io_pipe_phv_out_data_107; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_107 <= trans_0_io_pipe_phv_out_data_107;
    end else begin
      amplifier_0_1_data_107 <= trans_1_io_pipe_phv_out_data_107;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_108 <= init_io_pipe_phv_out_data_108; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_108 <= trans_0_io_pipe_phv_out_data_108;
    end else begin
      amplifier_0_1_data_108 <= trans_1_io_pipe_phv_out_data_108;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_109 <= init_io_pipe_phv_out_data_109; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_109 <= trans_0_io_pipe_phv_out_data_109;
    end else begin
      amplifier_0_1_data_109 <= trans_1_io_pipe_phv_out_data_109;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_110 <= init_io_pipe_phv_out_data_110; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_110 <= trans_0_io_pipe_phv_out_data_110;
    end else begin
      amplifier_0_1_data_110 <= trans_1_io_pipe_phv_out_data_110;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_111 <= init_io_pipe_phv_out_data_111; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_111 <= trans_0_io_pipe_phv_out_data_111;
    end else begin
      amplifier_0_1_data_111 <= trans_1_io_pipe_phv_out_data_111;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_112 <= init_io_pipe_phv_out_data_112; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_112 <= trans_0_io_pipe_phv_out_data_112;
    end else begin
      amplifier_0_1_data_112 <= trans_1_io_pipe_phv_out_data_112;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_113 <= init_io_pipe_phv_out_data_113; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_113 <= trans_0_io_pipe_phv_out_data_113;
    end else begin
      amplifier_0_1_data_113 <= trans_1_io_pipe_phv_out_data_113;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_114 <= init_io_pipe_phv_out_data_114; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_114 <= trans_0_io_pipe_phv_out_data_114;
    end else begin
      amplifier_0_1_data_114 <= trans_1_io_pipe_phv_out_data_114;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_115 <= init_io_pipe_phv_out_data_115; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_115 <= trans_0_io_pipe_phv_out_data_115;
    end else begin
      amplifier_0_1_data_115 <= trans_1_io_pipe_phv_out_data_115;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_116 <= init_io_pipe_phv_out_data_116; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_116 <= trans_0_io_pipe_phv_out_data_116;
    end else begin
      amplifier_0_1_data_116 <= trans_1_io_pipe_phv_out_data_116;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_117 <= init_io_pipe_phv_out_data_117; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_117 <= trans_0_io_pipe_phv_out_data_117;
    end else begin
      amplifier_0_1_data_117 <= trans_1_io_pipe_phv_out_data_117;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_118 <= init_io_pipe_phv_out_data_118; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_118 <= trans_0_io_pipe_phv_out_data_118;
    end else begin
      amplifier_0_1_data_118 <= trans_1_io_pipe_phv_out_data_118;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_119 <= init_io_pipe_phv_out_data_119; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_119 <= trans_0_io_pipe_phv_out_data_119;
    end else begin
      amplifier_0_1_data_119 <= trans_1_io_pipe_phv_out_data_119;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_120 <= init_io_pipe_phv_out_data_120; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_120 <= trans_0_io_pipe_phv_out_data_120;
    end else begin
      amplifier_0_1_data_120 <= trans_1_io_pipe_phv_out_data_120;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_121 <= init_io_pipe_phv_out_data_121; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_121 <= trans_0_io_pipe_phv_out_data_121;
    end else begin
      amplifier_0_1_data_121 <= trans_1_io_pipe_phv_out_data_121;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_122 <= init_io_pipe_phv_out_data_122; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_122 <= trans_0_io_pipe_phv_out_data_122;
    end else begin
      amplifier_0_1_data_122 <= trans_1_io_pipe_phv_out_data_122;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_123 <= init_io_pipe_phv_out_data_123; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_123 <= trans_0_io_pipe_phv_out_data_123;
    end else begin
      amplifier_0_1_data_123 <= trans_1_io_pipe_phv_out_data_123;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_124 <= init_io_pipe_phv_out_data_124; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_124 <= trans_0_io_pipe_phv_out_data_124;
    end else begin
      amplifier_0_1_data_124 <= trans_1_io_pipe_phv_out_data_124;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_125 <= init_io_pipe_phv_out_data_125; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_125 <= trans_0_io_pipe_phv_out_data_125;
    end else begin
      amplifier_0_1_data_125 <= trans_1_io_pipe_phv_out_data_125;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_126 <= init_io_pipe_phv_out_data_126; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_126 <= trans_0_io_pipe_phv_out_data_126;
    end else begin
      amplifier_0_1_data_126 <= trans_1_io_pipe_phv_out_data_126;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_127 <= init_io_pipe_phv_out_data_127; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_127 <= trans_0_io_pipe_phv_out_data_127;
    end else begin
      amplifier_0_1_data_127 <= trans_1_io_pipe_phv_out_data_127;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_128 <= init_io_pipe_phv_out_data_128; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_128 <= trans_0_io_pipe_phv_out_data_128;
    end else begin
      amplifier_0_1_data_128 <= trans_1_io_pipe_phv_out_data_128;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_129 <= init_io_pipe_phv_out_data_129; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_129 <= trans_0_io_pipe_phv_out_data_129;
    end else begin
      amplifier_0_1_data_129 <= trans_1_io_pipe_phv_out_data_129;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_130 <= init_io_pipe_phv_out_data_130; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_130 <= trans_0_io_pipe_phv_out_data_130;
    end else begin
      amplifier_0_1_data_130 <= trans_1_io_pipe_phv_out_data_130;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_131 <= init_io_pipe_phv_out_data_131; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_131 <= trans_0_io_pipe_phv_out_data_131;
    end else begin
      amplifier_0_1_data_131 <= trans_1_io_pipe_phv_out_data_131;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_132 <= init_io_pipe_phv_out_data_132; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_132 <= trans_0_io_pipe_phv_out_data_132;
    end else begin
      amplifier_0_1_data_132 <= trans_1_io_pipe_phv_out_data_132;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_133 <= init_io_pipe_phv_out_data_133; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_133 <= trans_0_io_pipe_phv_out_data_133;
    end else begin
      amplifier_0_1_data_133 <= trans_1_io_pipe_phv_out_data_133;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_134 <= init_io_pipe_phv_out_data_134; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_134 <= trans_0_io_pipe_phv_out_data_134;
    end else begin
      amplifier_0_1_data_134 <= trans_1_io_pipe_phv_out_data_134;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_135 <= init_io_pipe_phv_out_data_135; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_135 <= trans_0_io_pipe_phv_out_data_135;
    end else begin
      amplifier_0_1_data_135 <= trans_1_io_pipe_phv_out_data_135;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_136 <= init_io_pipe_phv_out_data_136; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_136 <= trans_0_io_pipe_phv_out_data_136;
    end else begin
      amplifier_0_1_data_136 <= trans_1_io_pipe_phv_out_data_136;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_137 <= init_io_pipe_phv_out_data_137; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_137 <= trans_0_io_pipe_phv_out_data_137;
    end else begin
      amplifier_0_1_data_137 <= trans_1_io_pipe_phv_out_data_137;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_138 <= init_io_pipe_phv_out_data_138; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_138 <= trans_0_io_pipe_phv_out_data_138;
    end else begin
      amplifier_0_1_data_138 <= trans_1_io_pipe_phv_out_data_138;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_139 <= init_io_pipe_phv_out_data_139; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_139 <= trans_0_io_pipe_phv_out_data_139;
    end else begin
      amplifier_0_1_data_139 <= trans_1_io_pipe_phv_out_data_139;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_140 <= init_io_pipe_phv_out_data_140; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_140 <= trans_0_io_pipe_phv_out_data_140;
    end else begin
      amplifier_0_1_data_140 <= trans_1_io_pipe_phv_out_data_140;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_141 <= init_io_pipe_phv_out_data_141; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_141 <= trans_0_io_pipe_phv_out_data_141;
    end else begin
      amplifier_0_1_data_141 <= trans_1_io_pipe_phv_out_data_141;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_142 <= init_io_pipe_phv_out_data_142; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_142 <= trans_0_io_pipe_phv_out_data_142;
    end else begin
      amplifier_0_1_data_142 <= trans_1_io_pipe_phv_out_data_142;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_143 <= init_io_pipe_phv_out_data_143; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_143 <= trans_0_io_pipe_phv_out_data_143;
    end else begin
      amplifier_0_1_data_143 <= trans_1_io_pipe_phv_out_data_143;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_144 <= init_io_pipe_phv_out_data_144; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_144 <= trans_0_io_pipe_phv_out_data_144;
    end else begin
      amplifier_0_1_data_144 <= trans_1_io_pipe_phv_out_data_144;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_145 <= init_io_pipe_phv_out_data_145; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_145 <= trans_0_io_pipe_phv_out_data_145;
    end else begin
      amplifier_0_1_data_145 <= trans_1_io_pipe_phv_out_data_145;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_146 <= init_io_pipe_phv_out_data_146; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_146 <= trans_0_io_pipe_phv_out_data_146;
    end else begin
      amplifier_0_1_data_146 <= trans_1_io_pipe_phv_out_data_146;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_147 <= init_io_pipe_phv_out_data_147; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_147 <= trans_0_io_pipe_phv_out_data_147;
    end else begin
      amplifier_0_1_data_147 <= trans_1_io_pipe_phv_out_data_147;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_148 <= init_io_pipe_phv_out_data_148; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_148 <= trans_0_io_pipe_phv_out_data_148;
    end else begin
      amplifier_0_1_data_148 <= trans_1_io_pipe_phv_out_data_148;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_149 <= init_io_pipe_phv_out_data_149; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_149 <= trans_0_io_pipe_phv_out_data_149;
    end else begin
      amplifier_0_1_data_149 <= trans_1_io_pipe_phv_out_data_149;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_150 <= init_io_pipe_phv_out_data_150; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_150 <= trans_0_io_pipe_phv_out_data_150;
    end else begin
      amplifier_0_1_data_150 <= trans_1_io_pipe_phv_out_data_150;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_151 <= init_io_pipe_phv_out_data_151; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_151 <= trans_0_io_pipe_phv_out_data_151;
    end else begin
      amplifier_0_1_data_151 <= trans_1_io_pipe_phv_out_data_151;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_152 <= init_io_pipe_phv_out_data_152; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_152 <= trans_0_io_pipe_phv_out_data_152;
    end else begin
      amplifier_0_1_data_152 <= trans_1_io_pipe_phv_out_data_152;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_153 <= init_io_pipe_phv_out_data_153; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_153 <= trans_0_io_pipe_phv_out_data_153;
    end else begin
      amplifier_0_1_data_153 <= trans_1_io_pipe_phv_out_data_153;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_154 <= init_io_pipe_phv_out_data_154; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_154 <= trans_0_io_pipe_phv_out_data_154;
    end else begin
      amplifier_0_1_data_154 <= trans_1_io_pipe_phv_out_data_154;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_155 <= init_io_pipe_phv_out_data_155; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_155 <= trans_0_io_pipe_phv_out_data_155;
    end else begin
      amplifier_0_1_data_155 <= trans_1_io_pipe_phv_out_data_155;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_156 <= init_io_pipe_phv_out_data_156; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_156 <= trans_0_io_pipe_phv_out_data_156;
    end else begin
      amplifier_0_1_data_156 <= trans_1_io_pipe_phv_out_data_156;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_157 <= init_io_pipe_phv_out_data_157; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_157 <= trans_0_io_pipe_phv_out_data_157;
    end else begin
      amplifier_0_1_data_157 <= trans_1_io_pipe_phv_out_data_157;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_158 <= init_io_pipe_phv_out_data_158; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_158 <= trans_0_io_pipe_phv_out_data_158;
    end else begin
      amplifier_0_1_data_158 <= trans_1_io_pipe_phv_out_data_158;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_159 <= init_io_pipe_phv_out_data_159; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_159 <= trans_0_io_pipe_phv_out_data_159;
    end else begin
      amplifier_0_1_data_159 <= trans_1_io_pipe_phv_out_data_159;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_160 <= init_io_pipe_phv_out_data_160; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_160 <= trans_0_io_pipe_phv_out_data_160;
    end else begin
      amplifier_0_1_data_160 <= trans_1_io_pipe_phv_out_data_160;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_161 <= init_io_pipe_phv_out_data_161; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_161 <= trans_0_io_pipe_phv_out_data_161;
    end else begin
      amplifier_0_1_data_161 <= trans_1_io_pipe_phv_out_data_161;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_162 <= init_io_pipe_phv_out_data_162; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_162 <= trans_0_io_pipe_phv_out_data_162;
    end else begin
      amplifier_0_1_data_162 <= trans_1_io_pipe_phv_out_data_162;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_163 <= init_io_pipe_phv_out_data_163; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_163 <= trans_0_io_pipe_phv_out_data_163;
    end else begin
      amplifier_0_1_data_163 <= trans_1_io_pipe_phv_out_data_163;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_164 <= init_io_pipe_phv_out_data_164; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_164 <= trans_0_io_pipe_phv_out_data_164;
    end else begin
      amplifier_0_1_data_164 <= trans_1_io_pipe_phv_out_data_164;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_165 <= init_io_pipe_phv_out_data_165; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_165 <= trans_0_io_pipe_phv_out_data_165;
    end else begin
      amplifier_0_1_data_165 <= trans_1_io_pipe_phv_out_data_165;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_166 <= init_io_pipe_phv_out_data_166; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_166 <= trans_0_io_pipe_phv_out_data_166;
    end else begin
      amplifier_0_1_data_166 <= trans_1_io_pipe_phv_out_data_166;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_167 <= init_io_pipe_phv_out_data_167; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_167 <= trans_0_io_pipe_phv_out_data_167;
    end else begin
      amplifier_0_1_data_167 <= trans_1_io_pipe_phv_out_data_167;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_168 <= init_io_pipe_phv_out_data_168; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_168 <= trans_0_io_pipe_phv_out_data_168;
    end else begin
      amplifier_0_1_data_168 <= trans_1_io_pipe_phv_out_data_168;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_169 <= init_io_pipe_phv_out_data_169; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_169 <= trans_0_io_pipe_phv_out_data_169;
    end else begin
      amplifier_0_1_data_169 <= trans_1_io_pipe_phv_out_data_169;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_170 <= init_io_pipe_phv_out_data_170; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_170 <= trans_0_io_pipe_phv_out_data_170;
    end else begin
      amplifier_0_1_data_170 <= trans_1_io_pipe_phv_out_data_170;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_171 <= init_io_pipe_phv_out_data_171; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_171 <= trans_0_io_pipe_phv_out_data_171;
    end else begin
      amplifier_0_1_data_171 <= trans_1_io_pipe_phv_out_data_171;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_172 <= init_io_pipe_phv_out_data_172; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_172 <= trans_0_io_pipe_phv_out_data_172;
    end else begin
      amplifier_0_1_data_172 <= trans_1_io_pipe_phv_out_data_172;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_173 <= init_io_pipe_phv_out_data_173; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_173 <= trans_0_io_pipe_phv_out_data_173;
    end else begin
      amplifier_0_1_data_173 <= trans_1_io_pipe_phv_out_data_173;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_174 <= init_io_pipe_phv_out_data_174; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_174 <= trans_0_io_pipe_phv_out_data_174;
    end else begin
      amplifier_0_1_data_174 <= trans_1_io_pipe_phv_out_data_174;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_175 <= init_io_pipe_phv_out_data_175; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_175 <= trans_0_io_pipe_phv_out_data_175;
    end else begin
      amplifier_0_1_data_175 <= trans_1_io_pipe_phv_out_data_175;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_176 <= init_io_pipe_phv_out_data_176; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_176 <= trans_0_io_pipe_phv_out_data_176;
    end else begin
      amplifier_0_1_data_176 <= trans_1_io_pipe_phv_out_data_176;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_177 <= init_io_pipe_phv_out_data_177; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_177 <= trans_0_io_pipe_phv_out_data_177;
    end else begin
      amplifier_0_1_data_177 <= trans_1_io_pipe_phv_out_data_177;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_178 <= init_io_pipe_phv_out_data_178; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_178 <= trans_0_io_pipe_phv_out_data_178;
    end else begin
      amplifier_0_1_data_178 <= trans_1_io_pipe_phv_out_data_178;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_179 <= init_io_pipe_phv_out_data_179; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_179 <= trans_0_io_pipe_phv_out_data_179;
    end else begin
      amplifier_0_1_data_179 <= trans_1_io_pipe_phv_out_data_179;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_180 <= init_io_pipe_phv_out_data_180; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_180 <= trans_0_io_pipe_phv_out_data_180;
    end else begin
      amplifier_0_1_data_180 <= trans_1_io_pipe_phv_out_data_180;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_181 <= init_io_pipe_phv_out_data_181; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_181 <= trans_0_io_pipe_phv_out_data_181;
    end else begin
      amplifier_0_1_data_181 <= trans_1_io_pipe_phv_out_data_181;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_182 <= init_io_pipe_phv_out_data_182; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_182 <= trans_0_io_pipe_phv_out_data_182;
    end else begin
      amplifier_0_1_data_182 <= trans_1_io_pipe_phv_out_data_182;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_183 <= init_io_pipe_phv_out_data_183; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_183 <= trans_0_io_pipe_phv_out_data_183;
    end else begin
      amplifier_0_1_data_183 <= trans_1_io_pipe_phv_out_data_183;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_184 <= init_io_pipe_phv_out_data_184; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_184 <= trans_0_io_pipe_phv_out_data_184;
    end else begin
      amplifier_0_1_data_184 <= trans_1_io_pipe_phv_out_data_184;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_185 <= init_io_pipe_phv_out_data_185; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_185 <= trans_0_io_pipe_phv_out_data_185;
    end else begin
      amplifier_0_1_data_185 <= trans_1_io_pipe_phv_out_data_185;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_186 <= init_io_pipe_phv_out_data_186; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_186 <= trans_0_io_pipe_phv_out_data_186;
    end else begin
      amplifier_0_1_data_186 <= trans_1_io_pipe_phv_out_data_186;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_187 <= init_io_pipe_phv_out_data_187; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_187 <= trans_0_io_pipe_phv_out_data_187;
    end else begin
      amplifier_0_1_data_187 <= trans_1_io_pipe_phv_out_data_187;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_188 <= init_io_pipe_phv_out_data_188; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_188 <= trans_0_io_pipe_phv_out_data_188;
    end else begin
      amplifier_0_1_data_188 <= trans_1_io_pipe_phv_out_data_188;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_189 <= init_io_pipe_phv_out_data_189; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_189 <= trans_0_io_pipe_phv_out_data_189;
    end else begin
      amplifier_0_1_data_189 <= trans_1_io_pipe_phv_out_data_189;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_190 <= init_io_pipe_phv_out_data_190; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_190 <= trans_0_io_pipe_phv_out_data_190;
    end else begin
      amplifier_0_1_data_190 <= trans_1_io_pipe_phv_out_data_190;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_191 <= init_io_pipe_phv_out_data_191; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_191 <= trans_0_io_pipe_phv_out_data_191;
    end else begin
      amplifier_0_1_data_191 <= trans_1_io_pipe_phv_out_data_191;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_192 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_192 <= trans_0_io_pipe_phv_out_data_192;
    end else begin
      amplifier_0_1_data_192 <= trans_1_io_pipe_phv_out_data_192;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_193 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_193 <= trans_0_io_pipe_phv_out_data_193;
    end else begin
      amplifier_0_1_data_193 <= trans_1_io_pipe_phv_out_data_193;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_194 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_194 <= trans_0_io_pipe_phv_out_data_194;
    end else begin
      amplifier_0_1_data_194 <= trans_1_io_pipe_phv_out_data_194;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_195 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_195 <= trans_0_io_pipe_phv_out_data_195;
    end else begin
      amplifier_0_1_data_195 <= trans_1_io_pipe_phv_out_data_195;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_196 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_196 <= trans_0_io_pipe_phv_out_data_196;
    end else begin
      amplifier_0_1_data_196 <= trans_1_io_pipe_phv_out_data_196;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_197 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_197 <= trans_0_io_pipe_phv_out_data_197;
    end else begin
      amplifier_0_1_data_197 <= trans_1_io_pipe_phv_out_data_197;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_198 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_198 <= trans_0_io_pipe_phv_out_data_198;
    end else begin
      amplifier_0_1_data_198 <= trans_1_io_pipe_phv_out_data_198;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_199 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_199 <= trans_0_io_pipe_phv_out_data_199;
    end else begin
      amplifier_0_1_data_199 <= trans_1_io_pipe_phv_out_data_199;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_200 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_200 <= trans_0_io_pipe_phv_out_data_200;
    end else begin
      amplifier_0_1_data_200 <= trans_1_io_pipe_phv_out_data_200;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_201 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_201 <= trans_0_io_pipe_phv_out_data_201;
    end else begin
      amplifier_0_1_data_201 <= trans_1_io_pipe_phv_out_data_201;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_202 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_202 <= trans_0_io_pipe_phv_out_data_202;
    end else begin
      amplifier_0_1_data_202 <= trans_1_io_pipe_phv_out_data_202;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_203 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_203 <= trans_0_io_pipe_phv_out_data_203;
    end else begin
      amplifier_0_1_data_203 <= trans_1_io_pipe_phv_out_data_203;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_204 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_204 <= trans_0_io_pipe_phv_out_data_204;
    end else begin
      amplifier_0_1_data_204 <= trans_1_io_pipe_phv_out_data_204;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_205 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_205 <= trans_0_io_pipe_phv_out_data_205;
    end else begin
      amplifier_0_1_data_205 <= trans_1_io_pipe_phv_out_data_205;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_206 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_206 <= trans_0_io_pipe_phv_out_data_206;
    end else begin
      amplifier_0_1_data_206 <= trans_1_io_pipe_phv_out_data_206;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_207 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_207 <= trans_0_io_pipe_phv_out_data_207;
    end else begin
      amplifier_0_1_data_207 <= trans_1_io_pipe_phv_out_data_207;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_208 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_208 <= trans_0_io_pipe_phv_out_data_208;
    end else begin
      amplifier_0_1_data_208 <= trans_1_io_pipe_phv_out_data_208;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_209 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_209 <= trans_0_io_pipe_phv_out_data_209;
    end else begin
      amplifier_0_1_data_209 <= trans_1_io_pipe_phv_out_data_209;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_210 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_210 <= trans_0_io_pipe_phv_out_data_210;
    end else begin
      amplifier_0_1_data_210 <= trans_1_io_pipe_phv_out_data_210;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_211 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_211 <= trans_0_io_pipe_phv_out_data_211;
    end else begin
      amplifier_0_1_data_211 <= trans_1_io_pipe_phv_out_data_211;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_212 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_212 <= trans_0_io_pipe_phv_out_data_212;
    end else begin
      amplifier_0_1_data_212 <= trans_1_io_pipe_phv_out_data_212;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_213 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_213 <= trans_0_io_pipe_phv_out_data_213;
    end else begin
      amplifier_0_1_data_213 <= trans_1_io_pipe_phv_out_data_213;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_214 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_214 <= trans_0_io_pipe_phv_out_data_214;
    end else begin
      amplifier_0_1_data_214 <= trans_1_io_pipe_phv_out_data_214;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_215 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_215 <= trans_0_io_pipe_phv_out_data_215;
    end else begin
      amplifier_0_1_data_215 <= trans_1_io_pipe_phv_out_data_215;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_216 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_216 <= trans_0_io_pipe_phv_out_data_216;
    end else begin
      amplifier_0_1_data_216 <= trans_1_io_pipe_phv_out_data_216;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_217 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_217 <= trans_0_io_pipe_phv_out_data_217;
    end else begin
      amplifier_0_1_data_217 <= trans_1_io_pipe_phv_out_data_217;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_218 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_218 <= trans_0_io_pipe_phv_out_data_218;
    end else begin
      amplifier_0_1_data_218 <= trans_1_io_pipe_phv_out_data_218;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_219 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_219 <= trans_0_io_pipe_phv_out_data_219;
    end else begin
      amplifier_0_1_data_219 <= trans_1_io_pipe_phv_out_data_219;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_220 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_220 <= trans_0_io_pipe_phv_out_data_220;
    end else begin
      amplifier_0_1_data_220 <= trans_1_io_pipe_phv_out_data_220;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_221 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_221 <= trans_0_io_pipe_phv_out_data_221;
    end else begin
      amplifier_0_1_data_221 <= trans_1_io_pipe_phv_out_data_221;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_222 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_222 <= trans_0_io_pipe_phv_out_data_222;
    end else begin
      amplifier_0_1_data_222 <= trans_1_io_pipe_phv_out_data_222;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_223 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_223 <= trans_0_io_pipe_phv_out_data_223;
    end else begin
      amplifier_0_1_data_223 <= trans_1_io_pipe_phv_out_data_223;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_224 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_224 <= trans_0_io_pipe_phv_out_data_224;
    end else begin
      amplifier_0_1_data_224 <= trans_1_io_pipe_phv_out_data_224;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_225 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_225 <= trans_0_io_pipe_phv_out_data_225;
    end else begin
      amplifier_0_1_data_225 <= trans_1_io_pipe_phv_out_data_225;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_226 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_226 <= trans_0_io_pipe_phv_out_data_226;
    end else begin
      amplifier_0_1_data_226 <= trans_1_io_pipe_phv_out_data_226;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_227 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_227 <= trans_0_io_pipe_phv_out_data_227;
    end else begin
      amplifier_0_1_data_227 <= trans_1_io_pipe_phv_out_data_227;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_228 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_228 <= trans_0_io_pipe_phv_out_data_228;
    end else begin
      amplifier_0_1_data_228 <= trans_1_io_pipe_phv_out_data_228;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_229 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_229 <= trans_0_io_pipe_phv_out_data_229;
    end else begin
      amplifier_0_1_data_229 <= trans_1_io_pipe_phv_out_data_229;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_230 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_230 <= trans_0_io_pipe_phv_out_data_230;
    end else begin
      amplifier_0_1_data_230 <= trans_1_io_pipe_phv_out_data_230;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_231 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_231 <= trans_0_io_pipe_phv_out_data_231;
    end else begin
      amplifier_0_1_data_231 <= trans_1_io_pipe_phv_out_data_231;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_232 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_232 <= trans_0_io_pipe_phv_out_data_232;
    end else begin
      amplifier_0_1_data_232 <= trans_1_io_pipe_phv_out_data_232;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_233 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_233 <= trans_0_io_pipe_phv_out_data_233;
    end else begin
      amplifier_0_1_data_233 <= trans_1_io_pipe_phv_out_data_233;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_234 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_234 <= trans_0_io_pipe_phv_out_data_234;
    end else begin
      amplifier_0_1_data_234 <= trans_1_io_pipe_phv_out_data_234;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_235 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_235 <= trans_0_io_pipe_phv_out_data_235;
    end else begin
      amplifier_0_1_data_235 <= trans_1_io_pipe_phv_out_data_235;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_236 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_236 <= trans_0_io_pipe_phv_out_data_236;
    end else begin
      amplifier_0_1_data_236 <= trans_1_io_pipe_phv_out_data_236;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_237 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_237 <= trans_0_io_pipe_phv_out_data_237;
    end else begin
      amplifier_0_1_data_237 <= trans_1_io_pipe_phv_out_data_237;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_238 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_238 <= trans_0_io_pipe_phv_out_data_238;
    end else begin
      amplifier_0_1_data_238 <= trans_1_io_pipe_phv_out_data_238;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_239 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_239 <= trans_0_io_pipe_phv_out_data_239;
    end else begin
      amplifier_0_1_data_239 <= trans_1_io_pipe_phv_out_data_239;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_240 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_240 <= trans_0_io_pipe_phv_out_data_240;
    end else begin
      amplifier_0_1_data_240 <= trans_1_io_pipe_phv_out_data_240;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_241 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_241 <= trans_0_io_pipe_phv_out_data_241;
    end else begin
      amplifier_0_1_data_241 <= trans_1_io_pipe_phv_out_data_241;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_242 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_242 <= trans_0_io_pipe_phv_out_data_242;
    end else begin
      amplifier_0_1_data_242 <= trans_1_io_pipe_phv_out_data_242;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_243 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_243 <= trans_0_io_pipe_phv_out_data_243;
    end else begin
      amplifier_0_1_data_243 <= trans_1_io_pipe_phv_out_data_243;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_244 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_244 <= trans_0_io_pipe_phv_out_data_244;
    end else begin
      amplifier_0_1_data_244 <= trans_1_io_pipe_phv_out_data_244;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_245 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_245 <= trans_0_io_pipe_phv_out_data_245;
    end else begin
      amplifier_0_1_data_245 <= trans_1_io_pipe_phv_out_data_245;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_246 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_246 <= trans_0_io_pipe_phv_out_data_246;
    end else begin
      amplifier_0_1_data_246 <= trans_1_io_pipe_phv_out_data_246;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_247 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_247 <= trans_0_io_pipe_phv_out_data_247;
    end else begin
      amplifier_0_1_data_247 <= trans_1_io_pipe_phv_out_data_247;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_248 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_248 <= trans_0_io_pipe_phv_out_data_248;
    end else begin
      amplifier_0_1_data_248 <= trans_1_io_pipe_phv_out_data_248;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_249 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_249 <= trans_0_io_pipe_phv_out_data_249;
    end else begin
      amplifier_0_1_data_249 <= trans_1_io_pipe_phv_out_data_249;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_250 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_250 <= trans_0_io_pipe_phv_out_data_250;
    end else begin
      amplifier_0_1_data_250 <= trans_1_io_pipe_phv_out_data_250;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_251 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_251 <= trans_0_io_pipe_phv_out_data_251;
    end else begin
      amplifier_0_1_data_251 <= trans_1_io_pipe_phv_out_data_251;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_252 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_252 <= trans_0_io_pipe_phv_out_data_252;
    end else begin
      amplifier_0_1_data_252 <= trans_1_io_pipe_phv_out_data_252;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_253 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_253 <= trans_0_io_pipe_phv_out_data_253;
    end else begin
      amplifier_0_1_data_253 <= trans_1_io_pipe_phv_out_data_253;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_254 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_254 <= trans_0_io_pipe_phv_out_data_254;
    end else begin
      amplifier_0_1_data_254 <= trans_1_io_pipe_phv_out_data_254;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_data_255 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_data_255 <= trans_0_io_pipe_phv_out_data_255;
    end else begin
      amplifier_0_1_data_255 <= trans_1_io_pipe_phv_out_data_255;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_header_0 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_header_0 <= trans_0_io_pipe_phv_out_header_0;
    end else begin
      amplifier_0_1_header_0 <= trans_1_io_pipe_phv_out_header_0;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_header_1 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_header_1 <= trans_0_io_pipe_phv_out_header_1;
    end else begin
      amplifier_0_1_header_1 <= trans_1_io_pipe_phv_out_header_1;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_header_2 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_header_2 <= trans_0_io_pipe_phv_out_header_2;
    end else begin
      amplifier_0_1_header_2 <= trans_1_io_pipe_phv_out_header_2;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_header_3 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_header_3 <= trans_0_io_pipe_phv_out_header_3;
    end else begin
      amplifier_0_1_header_3 <= trans_1_io_pipe_phv_out_header_3;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_header_4 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_header_4 <= trans_0_io_pipe_phv_out_header_4;
    end else begin
      amplifier_0_1_header_4 <= trans_1_io_pipe_phv_out_header_4;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_header_5 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_header_5 <= trans_0_io_pipe_phv_out_header_5;
    end else begin
      amplifier_0_1_header_5 <= trans_1_io_pipe_phv_out_header_5;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_header_6 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_header_6 <= trans_0_io_pipe_phv_out_header_6;
    end else begin
      amplifier_0_1_header_6 <= trans_1_io_pipe_phv_out_header_6;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_header_7 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_header_7 <= trans_0_io_pipe_phv_out_header_7;
    end else begin
      amplifier_0_1_header_7 <= trans_1_io_pipe_phv_out_header_7;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_header_8 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_header_8 <= trans_0_io_pipe_phv_out_header_8;
    end else begin
      amplifier_0_1_header_8 <= trans_1_io_pipe_phv_out_header_8;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_header_9 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_header_9 <= trans_0_io_pipe_phv_out_header_9;
    end else begin
      amplifier_0_1_header_9 <= trans_1_io_pipe_phv_out_header_9;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_header_10 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_header_10 <= trans_0_io_pipe_phv_out_header_10;
    end else begin
      amplifier_0_1_header_10 <= trans_1_io_pipe_phv_out_header_10;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_header_11 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_header_11 <= trans_0_io_pipe_phv_out_header_11;
    end else begin
      amplifier_0_1_header_11 <= trans_1_io_pipe_phv_out_header_11;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_header_12 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_header_12 <= trans_0_io_pipe_phv_out_header_12;
    end else begin
      amplifier_0_1_header_12 <= trans_1_io_pipe_phv_out_header_12;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_header_13 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_header_13 <= trans_0_io_pipe_phv_out_header_13;
    end else begin
      amplifier_0_1_header_13 <= trans_1_io_pipe_phv_out_header_13;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_header_14 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_header_14 <= trans_0_io_pipe_phv_out_header_14;
    end else begin
      amplifier_0_1_header_14 <= trans_1_io_pipe_phv_out_header_14;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_header_15 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_header_15 <= trans_0_io_pipe_phv_out_header_15;
    end else begin
      amplifier_0_1_header_15 <= trans_1_io_pipe_phv_out_header_15;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_parse_current_state <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_parse_current_state <= trans_0_io_pipe_phv_out_parse_current_state;
    end else begin
      amplifier_0_1_parse_current_state <= trans_1_io_pipe_phv_out_parse_current_state;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_parse_current_offset <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_parse_current_offset <= trans_0_io_pipe_phv_out_parse_current_offset;
    end else begin
      amplifier_0_1_parse_current_offset <= trans_1_io_pipe_phv_out_parse_current_offset;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_parse_transition_field <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_parse_transition_field <= trans_0_io_pipe_phv_out_parse_transition_field;
    end else begin
      amplifier_0_1_parse_transition_field <= trans_1_io_pipe_phv_out_parse_transition_field;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_next_processor_id <= init_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_next_processor_id <= trans_0_io_pipe_phv_out_next_processor_id;
    end else begin
      amplifier_0_1_next_processor_id <= trans_1_io_pipe_phv_out_next_processor_id;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_next_config_id <= 1'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_next_config_id <= trans_0_io_pipe_phv_out_next_config_id;
    end else begin
      amplifier_0_1_next_config_id <= trans_1_io_pipe_phv_out_next_config_id;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      amplifier_0_1_is_valid_processor <= 1'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 116:31]
      amplifier_0_1_is_valid_processor <= trans_0_io_pipe_phv_out_is_valid_processor;
    end else begin
      amplifier_0_1_is_valid_processor <= trans_1_io_pipe_phv_out_is_valid_processor;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_0 <= init_io_pipe_phv_out_data_0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_0 <= trans_3_io_pipe_phv_out_data_0;
    end else begin
      amplifier_0_2_data_0 <= trans_2_io_pipe_phv_out_data_0;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_1 <= init_io_pipe_phv_out_data_1; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_1 <= trans_3_io_pipe_phv_out_data_1;
    end else begin
      amplifier_0_2_data_1 <= trans_2_io_pipe_phv_out_data_1;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_2 <= init_io_pipe_phv_out_data_2; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_2 <= trans_3_io_pipe_phv_out_data_2;
    end else begin
      amplifier_0_2_data_2 <= trans_2_io_pipe_phv_out_data_2;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_3 <= init_io_pipe_phv_out_data_3; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_3 <= trans_3_io_pipe_phv_out_data_3;
    end else begin
      amplifier_0_2_data_3 <= trans_2_io_pipe_phv_out_data_3;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_4 <= init_io_pipe_phv_out_data_4; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_4 <= trans_3_io_pipe_phv_out_data_4;
    end else begin
      amplifier_0_2_data_4 <= trans_2_io_pipe_phv_out_data_4;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_5 <= init_io_pipe_phv_out_data_5; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_5 <= trans_3_io_pipe_phv_out_data_5;
    end else begin
      amplifier_0_2_data_5 <= trans_2_io_pipe_phv_out_data_5;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_6 <= init_io_pipe_phv_out_data_6; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_6 <= trans_3_io_pipe_phv_out_data_6;
    end else begin
      amplifier_0_2_data_6 <= trans_2_io_pipe_phv_out_data_6;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_7 <= init_io_pipe_phv_out_data_7; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_7 <= trans_3_io_pipe_phv_out_data_7;
    end else begin
      amplifier_0_2_data_7 <= trans_2_io_pipe_phv_out_data_7;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_8 <= init_io_pipe_phv_out_data_8; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_8 <= trans_3_io_pipe_phv_out_data_8;
    end else begin
      amplifier_0_2_data_8 <= trans_2_io_pipe_phv_out_data_8;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_9 <= init_io_pipe_phv_out_data_9; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_9 <= trans_3_io_pipe_phv_out_data_9;
    end else begin
      amplifier_0_2_data_9 <= trans_2_io_pipe_phv_out_data_9;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_10 <= init_io_pipe_phv_out_data_10; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_10 <= trans_3_io_pipe_phv_out_data_10;
    end else begin
      amplifier_0_2_data_10 <= trans_2_io_pipe_phv_out_data_10;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_11 <= init_io_pipe_phv_out_data_11; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_11 <= trans_3_io_pipe_phv_out_data_11;
    end else begin
      amplifier_0_2_data_11 <= trans_2_io_pipe_phv_out_data_11;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_12 <= init_io_pipe_phv_out_data_12; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_12 <= trans_3_io_pipe_phv_out_data_12;
    end else begin
      amplifier_0_2_data_12 <= trans_2_io_pipe_phv_out_data_12;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_13 <= init_io_pipe_phv_out_data_13; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_13 <= trans_3_io_pipe_phv_out_data_13;
    end else begin
      amplifier_0_2_data_13 <= trans_2_io_pipe_phv_out_data_13;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_14 <= init_io_pipe_phv_out_data_14; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_14 <= trans_3_io_pipe_phv_out_data_14;
    end else begin
      amplifier_0_2_data_14 <= trans_2_io_pipe_phv_out_data_14;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_15 <= init_io_pipe_phv_out_data_15; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_15 <= trans_3_io_pipe_phv_out_data_15;
    end else begin
      amplifier_0_2_data_15 <= trans_2_io_pipe_phv_out_data_15;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_16 <= init_io_pipe_phv_out_data_16; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_16 <= trans_3_io_pipe_phv_out_data_16;
    end else begin
      amplifier_0_2_data_16 <= trans_2_io_pipe_phv_out_data_16;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_17 <= init_io_pipe_phv_out_data_17; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_17 <= trans_3_io_pipe_phv_out_data_17;
    end else begin
      amplifier_0_2_data_17 <= trans_2_io_pipe_phv_out_data_17;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_18 <= init_io_pipe_phv_out_data_18; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_18 <= trans_3_io_pipe_phv_out_data_18;
    end else begin
      amplifier_0_2_data_18 <= trans_2_io_pipe_phv_out_data_18;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_19 <= init_io_pipe_phv_out_data_19; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_19 <= trans_3_io_pipe_phv_out_data_19;
    end else begin
      amplifier_0_2_data_19 <= trans_2_io_pipe_phv_out_data_19;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_20 <= init_io_pipe_phv_out_data_20; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_20 <= trans_3_io_pipe_phv_out_data_20;
    end else begin
      amplifier_0_2_data_20 <= trans_2_io_pipe_phv_out_data_20;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_21 <= init_io_pipe_phv_out_data_21; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_21 <= trans_3_io_pipe_phv_out_data_21;
    end else begin
      amplifier_0_2_data_21 <= trans_2_io_pipe_phv_out_data_21;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_22 <= init_io_pipe_phv_out_data_22; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_22 <= trans_3_io_pipe_phv_out_data_22;
    end else begin
      amplifier_0_2_data_22 <= trans_2_io_pipe_phv_out_data_22;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_23 <= init_io_pipe_phv_out_data_23; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_23 <= trans_3_io_pipe_phv_out_data_23;
    end else begin
      amplifier_0_2_data_23 <= trans_2_io_pipe_phv_out_data_23;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_24 <= init_io_pipe_phv_out_data_24; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_24 <= trans_3_io_pipe_phv_out_data_24;
    end else begin
      amplifier_0_2_data_24 <= trans_2_io_pipe_phv_out_data_24;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_25 <= init_io_pipe_phv_out_data_25; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_25 <= trans_3_io_pipe_phv_out_data_25;
    end else begin
      amplifier_0_2_data_25 <= trans_2_io_pipe_phv_out_data_25;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_26 <= init_io_pipe_phv_out_data_26; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_26 <= trans_3_io_pipe_phv_out_data_26;
    end else begin
      amplifier_0_2_data_26 <= trans_2_io_pipe_phv_out_data_26;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_27 <= init_io_pipe_phv_out_data_27; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_27 <= trans_3_io_pipe_phv_out_data_27;
    end else begin
      amplifier_0_2_data_27 <= trans_2_io_pipe_phv_out_data_27;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_28 <= init_io_pipe_phv_out_data_28; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_28 <= trans_3_io_pipe_phv_out_data_28;
    end else begin
      amplifier_0_2_data_28 <= trans_2_io_pipe_phv_out_data_28;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_29 <= init_io_pipe_phv_out_data_29; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_29 <= trans_3_io_pipe_phv_out_data_29;
    end else begin
      amplifier_0_2_data_29 <= trans_2_io_pipe_phv_out_data_29;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_30 <= init_io_pipe_phv_out_data_30; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_30 <= trans_3_io_pipe_phv_out_data_30;
    end else begin
      amplifier_0_2_data_30 <= trans_2_io_pipe_phv_out_data_30;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_31 <= init_io_pipe_phv_out_data_31; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_31 <= trans_3_io_pipe_phv_out_data_31;
    end else begin
      amplifier_0_2_data_31 <= trans_2_io_pipe_phv_out_data_31;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_32 <= init_io_pipe_phv_out_data_32; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_32 <= trans_3_io_pipe_phv_out_data_32;
    end else begin
      amplifier_0_2_data_32 <= trans_2_io_pipe_phv_out_data_32;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_33 <= init_io_pipe_phv_out_data_33; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_33 <= trans_3_io_pipe_phv_out_data_33;
    end else begin
      amplifier_0_2_data_33 <= trans_2_io_pipe_phv_out_data_33;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_34 <= init_io_pipe_phv_out_data_34; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_34 <= trans_3_io_pipe_phv_out_data_34;
    end else begin
      amplifier_0_2_data_34 <= trans_2_io_pipe_phv_out_data_34;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_35 <= init_io_pipe_phv_out_data_35; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_35 <= trans_3_io_pipe_phv_out_data_35;
    end else begin
      amplifier_0_2_data_35 <= trans_2_io_pipe_phv_out_data_35;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_36 <= init_io_pipe_phv_out_data_36; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_36 <= trans_3_io_pipe_phv_out_data_36;
    end else begin
      amplifier_0_2_data_36 <= trans_2_io_pipe_phv_out_data_36;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_37 <= init_io_pipe_phv_out_data_37; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_37 <= trans_3_io_pipe_phv_out_data_37;
    end else begin
      amplifier_0_2_data_37 <= trans_2_io_pipe_phv_out_data_37;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_38 <= init_io_pipe_phv_out_data_38; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_38 <= trans_3_io_pipe_phv_out_data_38;
    end else begin
      amplifier_0_2_data_38 <= trans_2_io_pipe_phv_out_data_38;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_39 <= init_io_pipe_phv_out_data_39; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_39 <= trans_3_io_pipe_phv_out_data_39;
    end else begin
      amplifier_0_2_data_39 <= trans_2_io_pipe_phv_out_data_39;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_40 <= init_io_pipe_phv_out_data_40; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_40 <= trans_3_io_pipe_phv_out_data_40;
    end else begin
      amplifier_0_2_data_40 <= trans_2_io_pipe_phv_out_data_40;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_41 <= init_io_pipe_phv_out_data_41; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_41 <= trans_3_io_pipe_phv_out_data_41;
    end else begin
      amplifier_0_2_data_41 <= trans_2_io_pipe_phv_out_data_41;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_42 <= init_io_pipe_phv_out_data_42; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_42 <= trans_3_io_pipe_phv_out_data_42;
    end else begin
      amplifier_0_2_data_42 <= trans_2_io_pipe_phv_out_data_42;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_43 <= init_io_pipe_phv_out_data_43; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_43 <= trans_3_io_pipe_phv_out_data_43;
    end else begin
      amplifier_0_2_data_43 <= trans_2_io_pipe_phv_out_data_43;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_44 <= init_io_pipe_phv_out_data_44; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_44 <= trans_3_io_pipe_phv_out_data_44;
    end else begin
      amplifier_0_2_data_44 <= trans_2_io_pipe_phv_out_data_44;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_45 <= init_io_pipe_phv_out_data_45; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_45 <= trans_3_io_pipe_phv_out_data_45;
    end else begin
      amplifier_0_2_data_45 <= trans_2_io_pipe_phv_out_data_45;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_46 <= init_io_pipe_phv_out_data_46; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_46 <= trans_3_io_pipe_phv_out_data_46;
    end else begin
      amplifier_0_2_data_46 <= trans_2_io_pipe_phv_out_data_46;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_47 <= init_io_pipe_phv_out_data_47; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_47 <= trans_3_io_pipe_phv_out_data_47;
    end else begin
      amplifier_0_2_data_47 <= trans_2_io_pipe_phv_out_data_47;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_48 <= init_io_pipe_phv_out_data_48; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_48 <= trans_3_io_pipe_phv_out_data_48;
    end else begin
      amplifier_0_2_data_48 <= trans_2_io_pipe_phv_out_data_48;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_49 <= init_io_pipe_phv_out_data_49; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_49 <= trans_3_io_pipe_phv_out_data_49;
    end else begin
      amplifier_0_2_data_49 <= trans_2_io_pipe_phv_out_data_49;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_50 <= init_io_pipe_phv_out_data_50; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_50 <= trans_3_io_pipe_phv_out_data_50;
    end else begin
      amplifier_0_2_data_50 <= trans_2_io_pipe_phv_out_data_50;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_51 <= init_io_pipe_phv_out_data_51; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_51 <= trans_3_io_pipe_phv_out_data_51;
    end else begin
      amplifier_0_2_data_51 <= trans_2_io_pipe_phv_out_data_51;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_52 <= init_io_pipe_phv_out_data_52; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_52 <= trans_3_io_pipe_phv_out_data_52;
    end else begin
      amplifier_0_2_data_52 <= trans_2_io_pipe_phv_out_data_52;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_53 <= init_io_pipe_phv_out_data_53; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_53 <= trans_3_io_pipe_phv_out_data_53;
    end else begin
      amplifier_0_2_data_53 <= trans_2_io_pipe_phv_out_data_53;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_54 <= init_io_pipe_phv_out_data_54; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_54 <= trans_3_io_pipe_phv_out_data_54;
    end else begin
      amplifier_0_2_data_54 <= trans_2_io_pipe_phv_out_data_54;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_55 <= init_io_pipe_phv_out_data_55; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_55 <= trans_3_io_pipe_phv_out_data_55;
    end else begin
      amplifier_0_2_data_55 <= trans_2_io_pipe_phv_out_data_55;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_56 <= init_io_pipe_phv_out_data_56; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_56 <= trans_3_io_pipe_phv_out_data_56;
    end else begin
      amplifier_0_2_data_56 <= trans_2_io_pipe_phv_out_data_56;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_57 <= init_io_pipe_phv_out_data_57; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_57 <= trans_3_io_pipe_phv_out_data_57;
    end else begin
      amplifier_0_2_data_57 <= trans_2_io_pipe_phv_out_data_57;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_58 <= init_io_pipe_phv_out_data_58; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_58 <= trans_3_io_pipe_phv_out_data_58;
    end else begin
      amplifier_0_2_data_58 <= trans_2_io_pipe_phv_out_data_58;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_59 <= init_io_pipe_phv_out_data_59; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_59 <= trans_3_io_pipe_phv_out_data_59;
    end else begin
      amplifier_0_2_data_59 <= trans_2_io_pipe_phv_out_data_59;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_60 <= init_io_pipe_phv_out_data_60; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_60 <= trans_3_io_pipe_phv_out_data_60;
    end else begin
      amplifier_0_2_data_60 <= trans_2_io_pipe_phv_out_data_60;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_61 <= init_io_pipe_phv_out_data_61; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_61 <= trans_3_io_pipe_phv_out_data_61;
    end else begin
      amplifier_0_2_data_61 <= trans_2_io_pipe_phv_out_data_61;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_62 <= init_io_pipe_phv_out_data_62; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_62 <= trans_3_io_pipe_phv_out_data_62;
    end else begin
      amplifier_0_2_data_62 <= trans_2_io_pipe_phv_out_data_62;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_63 <= init_io_pipe_phv_out_data_63; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_63 <= trans_3_io_pipe_phv_out_data_63;
    end else begin
      amplifier_0_2_data_63 <= trans_2_io_pipe_phv_out_data_63;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_64 <= init_io_pipe_phv_out_data_64; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_64 <= trans_3_io_pipe_phv_out_data_64;
    end else begin
      amplifier_0_2_data_64 <= trans_2_io_pipe_phv_out_data_64;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_65 <= init_io_pipe_phv_out_data_65; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_65 <= trans_3_io_pipe_phv_out_data_65;
    end else begin
      amplifier_0_2_data_65 <= trans_2_io_pipe_phv_out_data_65;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_66 <= init_io_pipe_phv_out_data_66; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_66 <= trans_3_io_pipe_phv_out_data_66;
    end else begin
      amplifier_0_2_data_66 <= trans_2_io_pipe_phv_out_data_66;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_67 <= init_io_pipe_phv_out_data_67; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_67 <= trans_3_io_pipe_phv_out_data_67;
    end else begin
      amplifier_0_2_data_67 <= trans_2_io_pipe_phv_out_data_67;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_68 <= init_io_pipe_phv_out_data_68; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_68 <= trans_3_io_pipe_phv_out_data_68;
    end else begin
      amplifier_0_2_data_68 <= trans_2_io_pipe_phv_out_data_68;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_69 <= init_io_pipe_phv_out_data_69; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_69 <= trans_3_io_pipe_phv_out_data_69;
    end else begin
      amplifier_0_2_data_69 <= trans_2_io_pipe_phv_out_data_69;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_70 <= init_io_pipe_phv_out_data_70; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_70 <= trans_3_io_pipe_phv_out_data_70;
    end else begin
      amplifier_0_2_data_70 <= trans_2_io_pipe_phv_out_data_70;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_71 <= init_io_pipe_phv_out_data_71; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_71 <= trans_3_io_pipe_phv_out_data_71;
    end else begin
      amplifier_0_2_data_71 <= trans_2_io_pipe_phv_out_data_71;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_72 <= init_io_pipe_phv_out_data_72; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_72 <= trans_3_io_pipe_phv_out_data_72;
    end else begin
      amplifier_0_2_data_72 <= trans_2_io_pipe_phv_out_data_72;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_73 <= init_io_pipe_phv_out_data_73; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_73 <= trans_3_io_pipe_phv_out_data_73;
    end else begin
      amplifier_0_2_data_73 <= trans_2_io_pipe_phv_out_data_73;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_74 <= init_io_pipe_phv_out_data_74; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_74 <= trans_3_io_pipe_phv_out_data_74;
    end else begin
      amplifier_0_2_data_74 <= trans_2_io_pipe_phv_out_data_74;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_75 <= init_io_pipe_phv_out_data_75; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_75 <= trans_3_io_pipe_phv_out_data_75;
    end else begin
      amplifier_0_2_data_75 <= trans_2_io_pipe_phv_out_data_75;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_76 <= init_io_pipe_phv_out_data_76; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_76 <= trans_3_io_pipe_phv_out_data_76;
    end else begin
      amplifier_0_2_data_76 <= trans_2_io_pipe_phv_out_data_76;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_77 <= init_io_pipe_phv_out_data_77; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_77 <= trans_3_io_pipe_phv_out_data_77;
    end else begin
      amplifier_0_2_data_77 <= trans_2_io_pipe_phv_out_data_77;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_78 <= init_io_pipe_phv_out_data_78; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_78 <= trans_3_io_pipe_phv_out_data_78;
    end else begin
      amplifier_0_2_data_78 <= trans_2_io_pipe_phv_out_data_78;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_79 <= init_io_pipe_phv_out_data_79; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_79 <= trans_3_io_pipe_phv_out_data_79;
    end else begin
      amplifier_0_2_data_79 <= trans_2_io_pipe_phv_out_data_79;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_80 <= init_io_pipe_phv_out_data_80; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_80 <= trans_3_io_pipe_phv_out_data_80;
    end else begin
      amplifier_0_2_data_80 <= trans_2_io_pipe_phv_out_data_80;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_81 <= init_io_pipe_phv_out_data_81; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_81 <= trans_3_io_pipe_phv_out_data_81;
    end else begin
      amplifier_0_2_data_81 <= trans_2_io_pipe_phv_out_data_81;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_82 <= init_io_pipe_phv_out_data_82; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_82 <= trans_3_io_pipe_phv_out_data_82;
    end else begin
      amplifier_0_2_data_82 <= trans_2_io_pipe_phv_out_data_82;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_83 <= init_io_pipe_phv_out_data_83; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_83 <= trans_3_io_pipe_phv_out_data_83;
    end else begin
      amplifier_0_2_data_83 <= trans_2_io_pipe_phv_out_data_83;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_84 <= init_io_pipe_phv_out_data_84; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_84 <= trans_3_io_pipe_phv_out_data_84;
    end else begin
      amplifier_0_2_data_84 <= trans_2_io_pipe_phv_out_data_84;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_85 <= init_io_pipe_phv_out_data_85; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_85 <= trans_3_io_pipe_phv_out_data_85;
    end else begin
      amplifier_0_2_data_85 <= trans_2_io_pipe_phv_out_data_85;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_86 <= init_io_pipe_phv_out_data_86; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_86 <= trans_3_io_pipe_phv_out_data_86;
    end else begin
      amplifier_0_2_data_86 <= trans_2_io_pipe_phv_out_data_86;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_87 <= init_io_pipe_phv_out_data_87; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_87 <= trans_3_io_pipe_phv_out_data_87;
    end else begin
      amplifier_0_2_data_87 <= trans_2_io_pipe_phv_out_data_87;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_88 <= init_io_pipe_phv_out_data_88; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_88 <= trans_3_io_pipe_phv_out_data_88;
    end else begin
      amplifier_0_2_data_88 <= trans_2_io_pipe_phv_out_data_88;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_89 <= init_io_pipe_phv_out_data_89; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_89 <= trans_3_io_pipe_phv_out_data_89;
    end else begin
      amplifier_0_2_data_89 <= trans_2_io_pipe_phv_out_data_89;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_90 <= init_io_pipe_phv_out_data_90; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_90 <= trans_3_io_pipe_phv_out_data_90;
    end else begin
      amplifier_0_2_data_90 <= trans_2_io_pipe_phv_out_data_90;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_91 <= init_io_pipe_phv_out_data_91; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_91 <= trans_3_io_pipe_phv_out_data_91;
    end else begin
      amplifier_0_2_data_91 <= trans_2_io_pipe_phv_out_data_91;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_92 <= init_io_pipe_phv_out_data_92; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_92 <= trans_3_io_pipe_phv_out_data_92;
    end else begin
      amplifier_0_2_data_92 <= trans_2_io_pipe_phv_out_data_92;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_93 <= init_io_pipe_phv_out_data_93; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_93 <= trans_3_io_pipe_phv_out_data_93;
    end else begin
      amplifier_0_2_data_93 <= trans_2_io_pipe_phv_out_data_93;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_94 <= init_io_pipe_phv_out_data_94; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_94 <= trans_3_io_pipe_phv_out_data_94;
    end else begin
      amplifier_0_2_data_94 <= trans_2_io_pipe_phv_out_data_94;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_95 <= init_io_pipe_phv_out_data_95; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_95 <= trans_3_io_pipe_phv_out_data_95;
    end else begin
      amplifier_0_2_data_95 <= trans_2_io_pipe_phv_out_data_95;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_96 <= init_io_pipe_phv_out_data_96; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_96 <= trans_3_io_pipe_phv_out_data_96;
    end else begin
      amplifier_0_2_data_96 <= trans_2_io_pipe_phv_out_data_96;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_97 <= init_io_pipe_phv_out_data_97; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_97 <= trans_3_io_pipe_phv_out_data_97;
    end else begin
      amplifier_0_2_data_97 <= trans_2_io_pipe_phv_out_data_97;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_98 <= init_io_pipe_phv_out_data_98; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_98 <= trans_3_io_pipe_phv_out_data_98;
    end else begin
      amplifier_0_2_data_98 <= trans_2_io_pipe_phv_out_data_98;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_99 <= init_io_pipe_phv_out_data_99; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_99 <= trans_3_io_pipe_phv_out_data_99;
    end else begin
      amplifier_0_2_data_99 <= trans_2_io_pipe_phv_out_data_99;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_100 <= init_io_pipe_phv_out_data_100; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_100 <= trans_3_io_pipe_phv_out_data_100;
    end else begin
      amplifier_0_2_data_100 <= trans_2_io_pipe_phv_out_data_100;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_101 <= init_io_pipe_phv_out_data_101; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_101 <= trans_3_io_pipe_phv_out_data_101;
    end else begin
      amplifier_0_2_data_101 <= trans_2_io_pipe_phv_out_data_101;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_102 <= init_io_pipe_phv_out_data_102; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_102 <= trans_3_io_pipe_phv_out_data_102;
    end else begin
      amplifier_0_2_data_102 <= trans_2_io_pipe_phv_out_data_102;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_103 <= init_io_pipe_phv_out_data_103; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_103 <= trans_3_io_pipe_phv_out_data_103;
    end else begin
      amplifier_0_2_data_103 <= trans_2_io_pipe_phv_out_data_103;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_104 <= init_io_pipe_phv_out_data_104; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_104 <= trans_3_io_pipe_phv_out_data_104;
    end else begin
      amplifier_0_2_data_104 <= trans_2_io_pipe_phv_out_data_104;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_105 <= init_io_pipe_phv_out_data_105; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_105 <= trans_3_io_pipe_phv_out_data_105;
    end else begin
      amplifier_0_2_data_105 <= trans_2_io_pipe_phv_out_data_105;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_106 <= init_io_pipe_phv_out_data_106; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_106 <= trans_3_io_pipe_phv_out_data_106;
    end else begin
      amplifier_0_2_data_106 <= trans_2_io_pipe_phv_out_data_106;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_107 <= init_io_pipe_phv_out_data_107; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_107 <= trans_3_io_pipe_phv_out_data_107;
    end else begin
      amplifier_0_2_data_107 <= trans_2_io_pipe_phv_out_data_107;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_108 <= init_io_pipe_phv_out_data_108; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_108 <= trans_3_io_pipe_phv_out_data_108;
    end else begin
      amplifier_0_2_data_108 <= trans_2_io_pipe_phv_out_data_108;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_109 <= init_io_pipe_phv_out_data_109; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_109 <= trans_3_io_pipe_phv_out_data_109;
    end else begin
      amplifier_0_2_data_109 <= trans_2_io_pipe_phv_out_data_109;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_110 <= init_io_pipe_phv_out_data_110; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_110 <= trans_3_io_pipe_phv_out_data_110;
    end else begin
      amplifier_0_2_data_110 <= trans_2_io_pipe_phv_out_data_110;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_111 <= init_io_pipe_phv_out_data_111; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_111 <= trans_3_io_pipe_phv_out_data_111;
    end else begin
      amplifier_0_2_data_111 <= trans_2_io_pipe_phv_out_data_111;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_112 <= init_io_pipe_phv_out_data_112; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_112 <= trans_3_io_pipe_phv_out_data_112;
    end else begin
      amplifier_0_2_data_112 <= trans_2_io_pipe_phv_out_data_112;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_113 <= init_io_pipe_phv_out_data_113; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_113 <= trans_3_io_pipe_phv_out_data_113;
    end else begin
      amplifier_0_2_data_113 <= trans_2_io_pipe_phv_out_data_113;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_114 <= init_io_pipe_phv_out_data_114; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_114 <= trans_3_io_pipe_phv_out_data_114;
    end else begin
      amplifier_0_2_data_114 <= trans_2_io_pipe_phv_out_data_114;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_115 <= init_io_pipe_phv_out_data_115; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_115 <= trans_3_io_pipe_phv_out_data_115;
    end else begin
      amplifier_0_2_data_115 <= trans_2_io_pipe_phv_out_data_115;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_116 <= init_io_pipe_phv_out_data_116; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_116 <= trans_3_io_pipe_phv_out_data_116;
    end else begin
      amplifier_0_2_data_116 <= trans_2_io_pipe_phv_out_data_116;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_117 <= init_io_pipe_phv_out_data_117; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_117 <= trans_3_io_pipe_phv_out_data_117;
    end else begin
      amplifier_0_2_data_117 <= trans_2_io_pipe_phv_out_data_117;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_118 <= init_io_pipe_phv_out_data_118; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_118 <= trans_3_io_pipe_phv_out_data_118;
    end else begin
      amplifier_0_2_data_118 <= trans_2_io_pipe_phv_out_data_118;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_119 <= init_io_pipe_phv_out_data_119; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_119 <= trans_3_io_pipe_phv_out_data_119;
    end else begin
      amplifier_0_2_data_119 <= trans_2_io_pipe_phv_out_data_119;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_120 <= init_io_pipe_phv_out_data_120; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_120 <= trans_3_io_pipe_phv_out_data_120;
    end else begin
      amplifier_0_2_data_120 <= trans_2_io_pipe_phv_out_data_120;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_121 <= init_io_pipe_phv_out_data_121; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_121 <= trans_3_io_pipe_phv_out_data_121;
    end else begin
      amplifier_0_2_data_121 <= trans_2_io_pipe_phv_out_data_121;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_122 <= init_io_pipe_phv_out_data_122; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_122 <= trans_3_io_pipe_phv_out_data_122;
    end else begin
      amplifier_0_2_data_122 <= trans_2_io_pipe_phv_out_data_122;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_123 <= init_io_pipe_phv_out_data_123; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_123 <= trans_3_io_pipe_phv_out_data_123;
    end else begin
      amplifier_0_2_data_123 <= trans_2_io_pipe_phv_out_data_123;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_124 <= init_io_pipe_phv_out_data_124; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_124 <= trans_3_io_pipe_phv_out_data_124;
    end else begin
      amplifier_0_2_data_124 <= trans_2_io_pipe_phv_out_data_124;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_125 <= init_io_pipe_phv_out_data_125; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_125 <= trans_3_io_pipe_phv_out_data_125;
    end else begin
      amplifier_0_2_data_125 <= trans_2_io_pipe_phv_out_data_125;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_126 <= init_io_pipe_phv_out_data_126; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_126 <= trans_3_io_pipe_phv_out_data_126;
    end else begin
      amplifier_0_2_data_126 <= trans_2_io_pipe_phv_out_data_126;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_127 <= init_io_pipe_phv_out_data_127; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_127 <= trans_3_io_pipe_phv_out_data_127;
    end else begin
      amplifier_0_2_data_127 <= trans_2_io_pipe_phv_out_data_127;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_128 <= init_io_pipe_phv_out_data_128; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_128 <= trans_3_io_pipe_phv_out_data_128;
    end else begin
      amplifier_0_2_data_128 <= trans_2_io_pipe_phv_out_data_128;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_129 <= init_io_pipe_phv_out_data_129; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_129 <= trans_3_io_pipe_phv_out_data_129;
    end else begin
      amplifier_0_2_data_129 <= trans_2_io_pipe_phv_out_data_129;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_130 <= init_io_pipe_phv_out_data_130; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_130 <= trans_3_io_pipe_phv_out_data_130;
    end else begin
      amplifier_0_2_data_130 <= trans_2_io_pipe_phv_out_data_130;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_131 <= init_io_pipe_phv_out_data_131; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_131 <= trans_3_io_pipe_phv_out_data_131;
    end else begin
      amplifier_0_2_data_131 <= trans_2_io_pipe_phv_out_data_131;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_132 <= init_io_pipe_phv_out_data_132; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_132 <= trans_3_io_pipe_phv_out_data_132;
    end else begin
      amplifier_0_2_data_132 <= trans_2_io_pipe_phv_out_data_132;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_133 <= init_io_pipe_phv_out_data_133; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_133 <= trans_3_io_pipe_phv_out_data_133;
    end else begin
      amplifier_0_2_data_133 <= trans_2_io_pipe_phv_out_data_133;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_134 <= init_io_pipe_phv_out_data_134; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_134 <= trans_3_io_pipe_phv_out_data_134;
    end else begin
      amplifier_0_2_data_134 <= trans_2_io_pipe_phv_out_data_134;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_135 <= init_io_pipe_phv_out_data_135; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_135 <= trans_3_io_pipe_phv_out_data_135;
    end else begin
      amplifier_0_2_data_135 <= trans_2_io_pipe_phv_out_data_135;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_136 <= init_io_pipe_phv_out_data_136; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_136 <= trans_3_io_pipe_phv_out_data_136;
    end else begin
      amplifier_0_2_data_136 <= trans_2_io_pipe_phv_out_data_136;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_137 <= init_io_pipe_phv_out_data_137; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_137 <= trans_3_io_pipe_phv_out_data_137;
    end else begin
      amplifier_0_2_data_137 <= trans_2_io_pipe_phv_out_data_137;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_138 <= init_io_pipe_phv_out_data_138; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_138 <= trans_3_io_pipe_phv_out_data_138;
    end else begin
      amplifier_0_2_data_138 <= trans_2_io_pipe_phv_out_data_138;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_139 <= init_io_pipe_phv_out_data_139; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_139 <= trans_3_io_pipe_phv_out_data_139;
    end else begin
      amplifier_0_2_data_139 <= trans_2_io_pipe_phv_out_data_139;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_140 <= init_io_pipe_phv_out_data_140; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_140 <= trans_3_io_pipe_phv_out_data_140;
    end else begin
      amplifier_0_2_data_140 <= trans_2_io_pipe_phv_out_data_140;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_141 <= init_io_pipe_phv_out_data_141; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_141 <= trans_3_io_pipe_phv_out_data_141;
    end else begin
      amplifier_0_2_data_141 <= trans_2_io_pipe_phv_out_data_141;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_142 <= init_io_pipe_phv_out_data_142; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_142 <= trans_3_io_pipe_phv_out_data_142;
    end else begin
      amplifier_0_2_data_142 <= trans_2_io_pipe_phv_out_data_142;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_143 <= init_io_pipe_phv_out_data_143; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_143 <= trans_3_io_pipe_phv_out_data_143;
    end else begin
      amplifier_0_2_data_143 <= trans_2_io_pipe_phv_out_data_143;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_144 <= init_io_pipe_phv_out_data_144; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_144 <= trans_3_io_pipe_phv_out_data_144;
    end else begin
      amplifier_0_2_data_144 <= trans_2_io_pipe_phv_out_data_144;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_145 <= init_io_pipe_phv_out_data_145; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_145 <= trans_3_io_pipe_phv_out_data_145;
    end else begin
      amplifier_0_2_data_145 <= trans_2_io_pipe_phv_out_data_145;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_146 <= init_io_pipe_phv_out_data_146; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_146 <= trans_3_io_pipe_phv_out_data_146;
    end else begin
      amplifier_0_2_data_146 <= trans_2_io_pipe_phv_out_data_146;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_147 <= init_io_pipe_phv_out_data_147; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_147 <= trans_3_io_pipe_phv_out_data_147;
    end else begin
      amplifier_0_2_data_147 <= trans_2_io_pipe_phv_out_data_147;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_148 <= init_io_pipe_phv_out_data_148; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_148 <= trans_3_io_pipe_phv_out_data_148;
    end else begin
      amplifier_0_2_data_148 <= trans_2_io_pipe_phv_out_data_148;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_149 <= init_io_pipe_phv_out_data_149; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_149 <= trans_3_io_pipe_phv_out_data_149;
    end else begin
      amplifier_0_2_data_149 <= trans_2_io_pipe_phv_out_data_149;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_150 <= init_io_pipe_phv_out_data_150; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_150 <= trans_3_io_pipe_phv_out_data_150;
    end else begin
      amplifier_0_2_data_150 <= trans_2_io_pipe_phv_out_data_150;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_151 <= init_io_pipe_phv_out_data_151; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_151 <= trans_3_io_pipe_phv_out_data_151;
    end else begin
      amplifier_0_2_data_151 <= trans_2_io_pipe_phv_out_data_151;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_152 <= init_io_pipe_phv_out_data_152; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_152 <= trans_3_io_pipe_phv_out_data_152;
    end else begin
      amplifier_0_2_data_152 <= trans_2_io_pipe_phv_out_data_152;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_153 <= init_io_pipe_phv_out_data_153; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_153 <= trans_3_io_pipe_phv_out_data_153;
    end else begin
      amplifier_0_2_data_153 <= trans_2_io_pipe_phv_out_data_153;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_154 <= init_io_pipe_phv_out_data_154; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_154 <= trans_3_io_pipe_phv_out_data_154;
    end else begin
      amplifier_0_2_data_154 <= trans_2_io_pipe_phv_out_data_154;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_155 <= init_io_pipe_phv_out_data_155; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_155 <= trans_3_io_pipe_phv_out_data_155;
    end else begin
      amplifier_0_2_data_155 <= trans_2_io_pipe_phv_out_data_155;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_156 <= init_io_pipe_phv_out_data_156; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_156 <= trans_3_io_pipe_phv_out_data_156;
    end else begin
      amplifier_0_2_data_156 <= trans_2_io_pipe_phv_out_data_156;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_157 <= init_io_pipe_phv_out_data_157; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_157 <= trans_3_io_pipe_phv_out_data_157;
    end else begin
      amplifier_0_2_data_157 <= trans_2_io_pipe_phv_out_data_157;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_158 <= init_io_pipe_phv_out_data_158; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_158 <= trans_3_io_pipe_phv_out_data_158;
    end else begin
      amplifier_0_2_data_158 <= trans_2_io_pipe_phv_out_data_158;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_159 <= init_io_pipe_phv_out_data_159; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_159 <= trans_3_io_pipe_phv_out_data_159;
    end else begin
      amplifier_0_2_data_159 <= trans_2_io_pipe_phv_out_data_159;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_160 <= init_io_pipe_phv_out_data_160; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_160 <= trans_3_io_pipe_phv_out_data_160;
    end else begin
      amplifier_0_2_data_160 <= trans_2_io_pipe_phv_out_data_160;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_161 <= init_io_pipe_phv_out_data_161; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_161 <= trans_3_io_pipe_phv_out_data_161;
    end else begin
      amplifier_0_2_data_161 <= trans_2_io_pipe_phv_out_data_161;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_162 <= init_io_pipe_phv_out_data_162; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_162 <= trans_3_io_pipe_phv_out_data_162;
    end else begin
      amplifier_0_2_data_162 <= trans_2_io_pipe_phv_out_data_162;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_163 <= init_io_pipe_phv_out_data_163; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_163 <= trans_3_io_pipe_phv_out_data_163;
    end else begin
      amplifier_0_2_data_163 <= trans_2_io_pipe_phv_out_data_163;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_164 <= init_io_pipe_phv_out_data_164; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_164 <= trans_3_io_pipe_phv_out_data_164;
    end else begin
      amplifier_0_2_data_164 <= trans_2_io_pipe_phv_out_data_164;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_165 <= init_io_pipe_phv_out_data_165; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_165 <= trans_3_io_pipe_phv_out_data_165;
    end else begin
      amplifier_0_2_data_165 <= trans_2_io_pipe_phv_out_data_165;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_166 <= init_io_pipe_phv_out_data_166; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_166 <= trans_3_io_pipe_phv_out_data_166;
    end else begin
      amplifier_0_2_data_166 <= trans_2_io_pipe_phv_out_data_166;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_167 <= init_io_pipe_phv_out_data_167; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_167 <= trans_3_io_pipe_phv_out_data_167;
    end else begin
      amplifier_0_2_data_167 <= trans_2_io_pipe_phv_out_data_167;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_168 <= init_io_pipe_phv_out_data_168; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_168 <= trans_3_io_pipe_phv_out_data_168;
    end else begin
      amplifier_0_2_data_168 <= trans_2_io_pipe_phv_out_data_168;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_169 <= init_io_pipe_phv_out_data_169; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_169 <= trans_3_io_pipe_phv_out_data_169;
    end else begin
      amplifier_0_2_data_169 <= trans_2_io_pipe_phv_out_data_169;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_170 <= init_io_pipe_phv_out_data_170; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_170 <= trans_3_io_pipe_phv_out_data_170;
    end else begin
      amplifier_0_2_data_170 <= trans_2_io_pipe_phv_out_data_170;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_171 <= init_io_pipe_phv_out_data_171; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_171 <= trans_3_io_pipe_phv_out_data_171;
    end else begin
      amplifier_0_2_data_171 <= trans_2_io_pipe_phv_out_data_171;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_172 <= init_io_pipe_phv_out_data_172; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_172 <= trans_3_io_pipe_phv_out_data_172;
    end else begin
      amplifier_0_2_data_172 <= trans_2_io_pipe_phv_out_data_172;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_173 <= init_io_pipe_phv_out_data_173; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_173 <= trans_3_io_pipe_phv_out_data_173;
    end else begin
      amplifier_0_2_data_173 <= trans_2_io_pipe_phv_out_data_173;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_174 <= init_io_pipe_phv_out_data_174; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_174 <= trans_3_io_pipe_phv_out_data_174;
    end else begin
      amplifier_0_2_data_174 <= trans_2_io_pipe_phv_out_data_174;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_175 <= init_io_pipe_phv_out_data_175; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_175 <= trans_3_io_pipe_phv_out_data_175;
    end else begin
      amplifier_0_2_data_175 <= trans_2_io_pipe_phv_out_data_175;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_176 <= init_io_pipe_phv_out_data_176; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_176 <= trans_3_io_pipe_phv_out_data_176;
    end else begin
      amplifier_0_2_data_176 <= trans_2_io_pipe_phv_out_data_176;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_177 <= init_io_pipe_phv_out_data_177; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_177 <= trans_3_io_pipe_phv_out_data_177;
    end else begin
      amplifier_0_2_data_177 <= trans_2_io_pipe_phv_out_data_177;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_178 <= init_io_pipe_phv_out_data_178; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_178 <= trans_3_io_pipe_phv_out_data_178;
    end else begin
      amplifier_0_2_data_178 <= trans_2_io_pipe_phv_out_data_178;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_179 <= init_io_pipe_phv_out_data_179; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_179 <= trans_3_io_pipe_phv_out_data_179;
    end else begin
      amplifier_0_2_data_179 <= trans_2_io_pipe_phv_out_data_179;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_180 <= init_io_pipe_phv_out_data_180; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_180 <= trans_3_io_pipe_phv_out_data_180;
    end else begin
      amplifier_0_2_data_180 <= trans_2_io_pipe_phv_out_data_180;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_181 <= init_io_pipe_phv_out_data_181; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_181 <= trans_3_io_pipe_phv_out_data_181;
    end else begin
      amplifier_0_2_data_181 <= trans_2_io_pipe_phv_out_data_181;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_182 <= init_io_pipe_phv_out_data_182; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_182 <= trans_3_io_pipe_phv_out_data_182;
    end else begin
      amplifier_0_2_data_182 <= trans_2_io_pipe_phv_out_data_182;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_183 <= init_io_pipe_phv_out_data_183; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_183 <= trans_3_io_pipe_phv_out_data_183;
    end else begin
      amplifier_0_2_data_183 <= trans_2_io_pipe_phv_out_data_183;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_184 <= init_io_pipe_phv_out_data_184; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_184 <= trans_3_io_pipe_phv_out_data_184;
    end else begin
      amplifier_0_2_data_184 <= trans_2_io_pipe_phv_out_data_184;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_185 <= init_io_pipe_phv_out_data_185; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_185 <= trans_3_io_pipe_phv_out_data_185;
    end else begin
      amplifier_0_2_data_185 <= trans_2_io_pipe_phv_out_data_185;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_186 <= init_io_pipe_phv_out_data_186; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_186 <= trans_3_io_pipe_phv_out_data_186;
    end else begin
      amplifier_0_2_data_186 <= trans_2_io_pipe_phv_out_data_186;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_187 <= init_io_pipe_phv_out_data_187; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_187 <= trans_3_io_pipe_phv_out_data_187;
    end else begin
      amplifier_0_2_data_187 <= trans_2_io_pipe_phv_out_data_187;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_188 <= init_io_pipe_phv_out_data_188; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_188 <= trans_3_io_pipe_phv_out_data_188;
    end else begin
      amplifier_0_2_data_188 <= trans_2_io_pipe_phv_out_data_188;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_189 <= init_io_pipe_phv_out_data_189; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_189 <= trans_3_io_pipe_phv_out_data_189;
    end else begin
      amplifier_0_2_data_189 <= trans_2_io_pipe_phv_out_data_189;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_190 <= init_io_pipe_phv_out_data_190; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_190 <= trans_3_io_pipe_phv_out_data_190;
    end else begin
      amplifier_0_2_data_190 <= trans_2_io_pipe_phv_out_data_190;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_191 <= init_io_pipe_phv_out_data_191; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_191 <= trans_3_io_pipe_phv_out_data_191;
    end else begin
      amplifier_0_2_data_191 <= trans_2_io_pipe_phv_out_data_191;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_192 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_192 <= trans_3_io_pipe_phv_out_data_192;
    end else begin
      amplifier_0_2_data_192 <= trans_2_io_pipe_phv_out_data_192;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_193 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_193 <= trans_3_io_pipe_phv_out_data_193;
    end else begin
      amplifier_0_2_data_193 <= trans_2_io_pipe_phv_out_data_193;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_194 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_194 <= trans_3_io_pipe_phv_out_data_194;
    end else begin
      amplifier_0_2_data_194 <= trans_2_io_pipe_phv_out_data_194;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_195 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_195 <= trans_3_io_pipe_phv_out_data_195;
    end else begin
      amplifier_0_2_data_195 <= trans_2_io_pipe_phv_out_data_195;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_196 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_196 <= trans_3_io_pipe_phv_out_data_196;
    end else begin
      amplifier_0_2_data_196 <= trans_2_io_pipe_phv_out_data_196;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_197 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_197 <= trans_3_io_pipe_phv_out_data_197;
    end else begin
      amplifier_0_2_data_197 <= trans_2_io_pipe_phv_out_data_197;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_198 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_198 <= trans_3_io_pipe_phv_out_data_198;
    end else begin
      amplifier_0_2_data_198 <= trans_2_io_pipe_phv_out_data_198;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_199 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_199 <= trans_3_io_pipe_phv_out_data_199;
    end else begin
      amplifier_0_2_data_199 <= trans_2_io_pipe_phv_out_data_199;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_200 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_200 <= trans_3_io_pipe_phv_out_data_200;
    end else begin
      amplifier_0_2_data_200 <= trans_2_io_pipe_phv_out_data_200;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_201 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_201 <= trans_3_io_pipe_phv_out_data_201;
    end else begin
      amplifier_0_2_data_201 <= trans_2_io_pipe_phv_out_data_201;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_202 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_202 <= trans_3_io_pipe_phv_out_data_202;
    end else begin
      amplifier_0_2_data_202 <= trans_2_io_pipe_phv_out_data_202;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_203 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_203 <= trans_3_io_pipe_phv_out_data_203;
    end else begin
      amplifier_0_2_data_203 <= trans_2_io_pipe_phv_out_data_203;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_204 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_204 <= trans_3_io_pipe_phv_out_data_204;
    end else begin
      amplifier_0_2_data_204 <= trans_2_io_pipe_phv_out_data_204;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_205 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_205 <= trans_3_io_pipe_phv_out_data_205;
    end else begin
      amplifier_0_2_data_205 <= trans_2_io_pipe_phv_out_data_205;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_206 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_206 <= trans_3_io_pipe_phv_out_data_206;
    end else begin
      amplifier_0_2_data_206 <= trans_2_io_pipe_phv_out_data_206;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_207 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_207 <= trans_3_io_pipe_phv_out_data_207;
    end else begin
      amplifier_0_2_data_207 <= trans_2_io_pipe_phv_out_data_207;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_208 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_208 <= trans_3_io_pipe_phv_out_data_208;
    end else begin
      amplifier_0_2_data_208 <= trans_2_io_pipe_phv_out_data_208;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_209 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_209 <= trans_3_io_pipe_phv_out_data_209;
    end else begin
      amplifier_0_2_data_209 <= trans_2_io_pipe_phv_out_data_209;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_210 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_210 <= trans_3_io_pipe_phv_out_data_210;
    end else begin
      amplifier_0_2_data_210 <= trans_2_io_pipe_phv_out_data_210;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_211 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_211 <= trans_3_io_pipe_phv_out_data_211;
    end else begin
      amplifier_0_2_data_211 <= trans_2_io_pipe_phv_out_data_211;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_212 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_212 <= trans_3_io_pipe_phv_out_data_212;
    end else begin
      amplifier_0_2_data_212 <= trans_2_io_pipe_phv_out_data_212;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_213 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_213 <= trans_3_io_pipe_phv_out_data_213;
    end else begin
      amplifier_0_2_data_213 <= trans_2_io_pipe_phv_out_data_213;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_214 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_214 <= trans_3_io_pipe_phv_out_data_214;
    end else begin
      amplifier_0_2_data_214 <= trans_2_io_pipe_phv_out_data_214;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_215 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_215 <= trans_3_io_pipe_phv_out_data_215;
    end else begin
      amplifier_0_2_data_215 <= trans_2_io_pipe_phv_out_data_215;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_216 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_216 <= trans_3_io_pipe_phv_out_data_216;
    end else begin
      amplifier_0_2_data_216 <= trans_2_io_pipe_phv_out_data_216;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_217 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_217 <= trans_3_io_pipe_phv_out_data_217;
    end else begin
      amplifier_0_2_data_217 <= trans_2_io_pipe_phv_out_data_217;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_218 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_218 <= trans_3_io_pipe_phv_out_data_218;
    end else begin
      amplifier_0_2_data_218 <= trans_2_io_pipe_phv_out_data_218;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_219 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_219 <= trans_3_io_pipe_phv_out_data_219;
    end else begin
      amplifier_0_2_data_219 <= trans_2_io_pipe_phv_out_data_219;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_220 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_220 <= trans_3_io_pipe_phv_out_data_220;
    end else begin
      amplifier_0_2_data_220 <= trans_2_io_pipe_phv_out_data_220;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_221 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_221 <= trans_3_io_pipe_phv_out_data_221;
    end else begin
      amplifier_0_2_data_221 <= trans_2_io_pipe_phv_out_data_221;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_222 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_222 <= trans_3_io_pipe_phv_out_data_222;
    end else begin
      amplifier_0_2_data_222 <= trans_2_io_pipe_phv_out_data_222;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_223 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_223 <= trans_3_io_pipe_phv_out_data_223;
    end else begin
      amplifier_0_2_data_223 <= trans_2_io_pipe_phv_out_data_223;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_224 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_224 <= trans_3_io_pipe_phv_out_data_224;
    end else begin
      amplifier_0_2_data_224 <= trans_2_io_pipe_phv_out_data_224;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_225 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_225 <= trans_3_io_pipe_phv_out_data_225;
    end else begin
      amplifier_0_2_data_225 <= trans_2_io_pipe_phv_out_data_225;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_226 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_226 <= trans_3_io_pipe_phv_out_data_226;
    end else begin
      amplifier_0_2_data_226 <= trans_2_io_pipe_phv_out_data_226;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_227 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_227 <= trans_3_io_pipe_phv_out_data_227;
    end else begin
      amplifier_0_2_data_227 <= trans_2_io_pipe_phv_out_data_227;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_228 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_228 <= trans_3_io_pipe_phv_out_data_228;
    end else begin
      amplifier_0_2_data_228 <= trans_2_io_pipe_phv_out_data_228;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_229 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_229 <= trans_3_io_pipe_phv_out_data_229;
    end else begin
      amplifier_0_2_data_229 <= trans_2_io_pipe_phv_out_data_229;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_230 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_230 <= trans_3_io_pipe_phv_out_data_230;
    end else begin
      amplifier_0_2_data_230 <= trans_2_io_pipe_phv_out_data_230;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_231 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_231 <= trans_3_io_pipe_phv_out_data_231;
    end else begin
      amplifier_0_2_data_231 <= trans_2_io_pipe_phv_out_data_231;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_232 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_232 <= trans_3_io_pipe_phv_out_data_232;
    end else begin
      amplifier_0_2_data_232 <= trans_2_io_pipe_phv_out_data_232;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_233 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_233 <= trans_3_io_pipe_phv_out_data_233;
    end else begin
      amplifier_0_2_data_233 <= trans_2_io_pipe_phv_out_data_233;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_234 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_234 <= trans_3_io_pipe_phv_out_data_234;
    end else begin
      amplifier_0_2_data_234 <= trans_2_io_pipe_phv_out_data_234;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_235 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_235 <= trans_3_io_pipe_phv_out_data_235;
    end else begin
      amplifier_0_2_data_235 <= trans_2_io_pipe_phv_out_data_235;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_236 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_236 <= trans_3_io_pipe_phv_out_data_236;
    end else begin
      amplifier_0_2_data_236 <= trans_2_io_pipe_phv_out_data_236;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_237 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_237 <= trans_3_io_pipe_phv_out_data_237;
    end else begin
      amplifier_0_2_data_237 <= trans_2_io_pipe_phv_out_data_237;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_238 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_238 <= trans_3_io_pipe_phv_out_data_238;
    end else begin
      amplifier_0_2_data_238 <= trans_2_io_pipe_phv_out_data_238;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_239 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_239 <= trans_3_io_pipe_phv_out_data_239;
    end else begin
      amplifier_0_2_data_239 <= trans_2_io_pipe_phv_out_data_239;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_240 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_240 <= trans_3_io_pipe_phv_out_data_240;
    end else begin
      amplifier_0_2_data_240 <= trans_2_io_pipe_phv_out_data_240;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_241 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_241 <= trans_3_io_pipe_phv_out_data_241;
    end else begin
      amplifier_0_2_data_241 <= trans_2_io_pipe_phv_out_data_241;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_242 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_242 <= trans_3_io_pipe_phv_out_data_242;
    end else begin
      amplifier_0_2_data_242 <= trans_2_io_pipe_phv_out_data_242;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_243 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_243 <= trans_3_io_pipe_phv_out_data_243;
    end else begin
      amplifier_0_2_data_243 <= trans_2_io_pipe_phv_out_data_243;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_244 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_244 <= trans_3_io_pipe_phv_out_data_244;
    end else begin
      amplifier_0_2_data_244 <= trans_2_io_pipe_phv_out_data_244;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_245 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_245 <= trans_3_io_pipe_phv_out_data_245;
    end else begin
      amplifier_0_2_data_245 <= trans_2_io_pipe_phv_out_data_245;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_246 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_246 <= trans_3_io_pipe_phv_out_data_246;
    end else begin
      amplifier_0_2_data_246 <= trans_2_io_pipe_phv_out_data_246;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_247 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_247 <= trans_3_io_pipe_phv_out_data_247;
    end else begin
      amplifier_0_2_data_247 <= trans_2_io_pipe_phv_out_data_247;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_248 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_248 <= trans_3_io_pipe_phv_out_data_248;
    end else begin
      amplifier_0_2_data_248 <= trans_2_io_pipe_phv_out_data_248;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_249 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_249 <= trans_3_io_pipe_phv_out_data_249;
    end else begin
      amplifier_0_2_data_249 <= trans_2_io_pipe_phv_out_data_249;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_250 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_250 <= trans_3_io_pipe_phv_out_data_250;
    end else begin
      amplifier_0_2_data_250 <= trans_2_io_pipe_phv_out_data_250;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_251 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_251 <= trans_3_io_pipe_phv_out_data_251;
    end else begin
      amplifier_0_2_data_251 <= trans_2_io_pipe_phv_out_data_251;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_252 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_252 <= trans_3_io_pipe_phv_out_data_252;
    end else begin
      amplifier_0_2_data_252 <= trans_2_io_pipe_phv_out_data_252;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_253 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_253 <= trans_3_io_pipe_phv_out_data_253;
    end else begin
      amplifier_0_2_data_253 <= trans_2_io_pipe_phv_out_data_253;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_254 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_254 <= trans_3_io_pipe_phv_out_data_254;
    end else begin
      amplifier_0_2_data_254 <= trans_2_io_pipe_phv_out_data_254;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_data_255 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_data_255 <= trans_3_io_pipe_phv_out_data_255;
    end else begin
      amplifier_0_2_data_255 <= trans_2_io_pipe_phv_out_data_255;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_header_0 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_header_0 <= trans_3_io_pipe_phv_out_header_0;
    end else begin
      amplifier_0_2_header_0 <= trans_2_io_pipe_phv_out_header_0;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_header_1 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_header_1 <= trans_3_io_pipe_phv_out_header_1;
    end else begin
      amplifier_0_2_header_1 <= trans_2_io_pipe_phv_out_header_1;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_header_2 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_header_2 <= trans_3_io_pipe_phv_out_header_2;
    end else begin
      amplifier_0_2_header_2 <= trans_2_io_pipe_phv_out_header_2;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_header_3 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_header_3 <= trans_3_io_pipe_phv_out_header_3;
    end else begin
      amplifier_0_2_header_3 <= trans_2_io_pipe_phv_out_header_3;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_header_4 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_header_4 <= trans_3_io_pipe_phv_out_header_4;
    end else begin
      amplifier_0_2_header_4 <= trans_2_io_pipe_phv_out_header_4;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_header_5 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_header_5 <= trans_3_io_pipe_phv_out_header_5;
    end else begin
      amplifier_0_2_header_5 <= trans_2_io_pipe_phv_out_header_5;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_header_6 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_header_6 <= trans_3_io_pipe_phv_out_header_6;
    end else begin
      amplifier_0_2_header_6 <= trans_2_io_pipe_phv_out_header_6;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_header_7 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_header_7 <= trans_3_io_pipe_phv_out_header_7;
    end else begin
      amplifier_0_2_header_7 <= trans_2_io_pipe_phv_out_header_7;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_header_8 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_header_8 <= trans_3_io_pipe_phv_out_header_8;
    end else begin
      amplifier_0_2_header_8 <= trans_2_io_pipe_phv_out_header_8;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_header_9 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_header_9 <= trans_3_io_pipe_phv_out_header_9;
    end else begin
      amplifier_0_2_header_9 <= trans_2_io_pipe_phv_out_header_9;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_header_10 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_header_10 <= trans_3_io_pipe_phv_out_header_10;
    end else begin
      amplifier_0_2_header_10 <= trans_2_io_pipe_phv_out_header_10;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_header_11 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_header_11 <= trans_3_io_pipe_phv_out_header_11;
    end else begin
      amplifier_0_2_header_11 <= trans_2_io_pipe_phv_out_header_11;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_header_12 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_header_12 <= trans_3_io_pipe_phv_out_header_12;
    end else begin
      amplifier_0_2_header_12 <= trans_2_io_pipe_phv_out_header_12;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_header_13 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_header_13 <= trans_3_io_pipe_phv_out_header_13;
    end else begin
      amplifier_0_2_header_13 <= trans_2_io_pipe_phv_out_header_13;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_header_14 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_header_14 <= trans_3_io_pipe_phv_out_header_14;
    end else begin
      amplifier_0_2_header_14 <= trans_2_io_pipe_phv_out_header_14;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_header_15 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_header_15 <= trans_3_io_pipe_phv_out_header_15;
    end else begin
      amplifier_0_2_header_15 <= trans_2_io_pipe_phv_out_header_15;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_parse_current_state <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_parse_current_state <= trans_3_io_pipe_phv_out_parse_current_state;
    end else begin
      amplifier_0_2_parse_current_state <= trans_2_io_pipe_phv_out_parse_current_state;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_parse_current_offset <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_parse_current_offset <= trans_3_io_pipe_phv_out_parse_current_offset;
    end else begin
      amplifier_0_2_parse_current_offset <= trans_2_io_pipe_phv_out_parse_current_offset;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_parse_transition_field <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_parse_transition_field <= trans_3_io_pipe_phv_out_parse_transition_field;
    end else begin
      amplifier_0_2_parse_transition_field <= trans_2_io_pipe_phv_out_parse_transition_field;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_next_processor_id <= init_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_next_processor_id <= trans_3_io_pipe_phv_out_next_processor_id;
    end else begin
      amplifier_0_2_next_processor_id <= trans_2_io_pipe_phv_out_next_processor_id;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_next_config_id <= 1'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_next_config_id <= trans_3_io_pipe_phv_out_next_config_id;
    end else begin
      amplifier_0_2_next_config_id <= trans_2_io_pipe_phv_out_next_config_id;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      amplifier_0_2_is_valid_processor <= 1'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 109:31]
      amplifier_0_2_is_valid_processor <= trans_3_io_pipe_phv_out_is_valid_processor;
    end else begin
      amplifier_0_2_is_valid_processor <= trans_2_io_pipe_phv_out_is_valid_processor;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_0 <= init_io_pipe_phv_out_data_0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_0 <= trans_2_io_pipe_phv_out_data_0;
    end else begin
      amplifier_0_3_data_0 <= trans_3_io_pipe_phv_out_data_0;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_1 <= init_io_pipe_phv_out_data_1; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_1 <= trans_2_io_pipe_phv_out_data_1;
    end else begin
      amplifier_0_3_data_1 <= trans_3_io_pipe_phv_out_data_1;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_2 <= init_io_pipe_phv_out_data_2; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_2 <= trans_2_io_pipe_phv_out_data_2;
    end else begin
      amplifier_0_3_data_2 <= trans_3_io_pipe_phv_out_data_2;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_3 <= init_io_pipe_phv_out_data_3; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_3 <= trans_2_io_pipe_phv_out_data_3;
    end else begin
      amplifier_0_3_data_3 <= trans_3_io_pipe_phv_out_data_3;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_4 <= init_io_pipe_phv_out_data_4; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_4 <= trans_2_io_pipe_phv_out_data_4;
    end else begin
      amplifier_0_3_data_4 <= trans_3_io_pipe_phv_out_data_4;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_5 <= init_io_pipe_phv_out_data_5; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_5 <= trans_2_io_pipe_phv_out_data_5;
    end else begin
      amplifier_0_3_data_5 <= trans_3_io_pipe_phv_out_data_5;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_6 <= init_io_pipe_phv_out_data_6; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_6 <= trans_2_io_pipe_phv_out_data_6;
    end else begin
      amplifier_0_3_data_6 <= trans_3_io_pipe_phv_out_data_6;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_7 <= init_io_pipe_phv_out_data_7; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_7 <= trans_2_io_pipe_phv_out_data_7;
    end else begin
      amplifier_0_3_data_7 <= trans_3_io_pipe_phv_out_data_7;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_8 <= init_io_pipe_phv_out_data_8; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_8 <= trans_2_io_pipe_phv_out_data_8;
    end else begin
      amplifier_0_3_data_8 <= trans_3_io_pipe_phv_out_data_8;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_9 <= init_io_pipe_phv_out_data_9; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_9 <= trans_2_io_pipe_phv_out_data_9;
    end else begin
      amplifier_0_3_data_9 <= trans_3_io_pipe_phv_out_data_9;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_10 <= init_io_pipe_phv_out_data_10; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_10 <= trans_2_io_pipe_phv_out_data_10;
    end else begin
      amplifier_0_3_data_10 <= trans_3_io_pipe_phv_out_data_10;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_11 <= init_io_pipe_phv_out_data_11; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_11 <= trans_2_io_pipe_phv_out_data_11;
    end else begin
      amplifier_0_3_data_11 <= trans_3_io_pipe_phv_out_data_11;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_12 <= init_io_pipe_phv_out_data_12; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_12 <= trans_2_io_pipe_phv_out_data_12;
    end else begin
      amplifier_0_3_data_12 <= trans_3_io_pipe_phv_out_data_12;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_13 <= init_io_pipe_phv_out_data_13; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_13 <= trans_2_io_pipe_phv_out_data_13;
    end else begin
      amplifier_0_3_data_13 <= trans_3_io_pipe_phv_out_data_13;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_14 <= init_io_pipe_phv_out_data_14; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_14 <= trans_2_io_pipe_phv_out_data_14;
    end else begin
      amplifier_0_3_data_14 <= trans_3_io_pipe_phv_out_data_14;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_15 <= init_io_pipe_phv_out_data_15; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_15 <= trans_2_io_pipe_phv_out_data_15;
    end else begin
      amplifier_0_3_data_15 <= trans_3_io_pipe_phv_out_data_15;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_16 <= init_io_pipe_phv_out_data_16; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_16 <= trans_2_io_pipe_phv_out_data_16;
    end else begin
      amplifier_0_3_data_16 <= trans_3_io_pipe_phv_out_data_16;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_17 <= init_io_pipe_phv_out_data_17; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_17 <= trans_2_io_pipe_phv_out_data_17;
    end else begin
      amplifier_0_3_data_17 <= trans_3_io_pipe_phv_out_data_17;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_18 <= init_io_pipe_phv_out_data_18; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_18 <= trans_2_io_pipe_phv_out_data_18;
    end else begin
      amplifier_0_3_data_18 <= trans_3_io_pipe_phv_out_data_18;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_19 <= init_io_pipe_phv_out_data_19; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_19 <= trans_2_io_pipe_phv_out_data_19;
    end else begin
      amplifier_0_3_data_19 <= trans_3_io_pipe_phv_out_data_19;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_20 <= init_io_pipe_phv_out_data_20; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_20 <= trans_2_io_pipe_phv_out_data_20;
    end else begin
      amplifier_0_3_data_20 <= trans_3_io_pipe_phv_out_data_20;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_21 <= init_io_pipe_phv_out_data_21; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_21 <= trans_2_io_pipe_phv_out_data_21;
    end else begin
      amplifier_0_3_data_21 <= trans_3_io_pipe_phv_out_data_21;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_22 <= init_io_pipe_phv_out_data_22; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_22 <= trans_2_io_pipe_phv_out_data_22;
    end else begin
      amplifier_0_3_data_22 <= trans_3_io_pipe_phv_out_data_22;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_23 <= init_io_pipe_phv_out_data_23; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_23 <= trans_2_io_pipe_phv_out_data_23;
    end else begin
      amplifier_0_3_data_23 <= trans_3_io_pipe_phv_out_data_23;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_24 <= init_io_pipe_phv_out_data_24; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_24 <= trans_2_io_pipe_phv_out_data_24;
    end else begin
      amplifier_0_3_data_24 <= trans_3_io_pipe_phv_out_data_24;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_25 <= init_io_pipe_phv_out_data_25; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_25 <= trans_2_io_pipe_phv_out_data_25;
    end else begin
      amplifier_0_3_data_25 <= trans_3_io_pipe_phv_out_data_25;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_26 <= init_io_pipe_phv_out_data_26; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_26 <= trans_2_io_pipe_phv_out_data_26;
    end else begin
      amplifier_0_3_data_26 <= trans_3_io_pipe_phv_out_data_26;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_27 <= init_io_pipe_phv_out_data_27; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_27 <= trans_2_io_pipe_phv_out_data_27;
    end else begin
      amplifier_0_3_data_27 <= trans_3_io_pipe_phv_out_data_27;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_28 <= init_io_pipe_phv_out_data_28; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_28 <= trans_2_io_pipe_phv_out_data_28;
    end else begin
      amplifier_0_3_data_28 <= trans_3_io_pipe_phv_out_data_28;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_29 <= init_io_pipe_phv_out_data_29; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_29 <= trans_2_io_pipe_phv_out_data_29;
    end else begin
      amplifier_0_3_data_29 <= trans_3_io_pipe_phv_out_data_29;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_30 <= init_io_pipe_phv_out_data_30; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_30 <= trans_2_io_pipe_phv_out_data_30;
    end else begin
      amplifier_0_3_data_30 <= trans_3_io_pipe_phv_out_data_30;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_31 <= init_io_pipe_phv_out_data_31; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_31 <= trans_2_io_pipe_phv_out_data_31;
    end else begin
      amplifier_0_3_data_31 <= trans_3_io_pipe_phv_out_data_31;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_32 <= init_io_pipe_phv_out_data_32; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_32 <= trans_2_io_pipe_phv_out_data_32;
    end else begin
      amplifier_0_3_data_32 <= trans_3_io_pipe_phv_out_data_32;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_33 <= init_io_pipe_phv_out_data_33; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_33 <= trans_2_io_pipe_phv_out_data_33;
    end else begin
      amplifier_0_3_data_33 <= trans_3_io_pipe_phv_out_data_33;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_34 <= init_io_pipe_phv_out_data_34; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_34 <= trans_2_io_pipe_phv_out_data_34;
    end else begin
      amplifier_0_3_data_34 <= trans_3_io_pipe_phv_out_data_34;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_35 <= init_io_pipe_phv_out_data_35; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_35 <= trans_2_io_pipe_phv_out_data_35;
    end else begin
      amplifier_0_3_data_35 <= trans_3_io_pipe_phv_out_data_35;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_36 <= init_io_pipe_phv_out_data_36; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_36 <= trans_2_io_pipe_phv_out_data_36;
    end else begin
      amplifier_0_3_data_36 <= trans_3_io_pipe_phv_out_data_36;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_37 <= init_io_pipe_phv_out_data_37; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_37 <= trans_2_io_pipe_phv_out_data_37;
    end else begin
      amplifier_0_3_data_37 <= trans_3_io_pipe_phv_out_data_37;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_38 <= init_io_pipe_phv_out_data_38; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_38 <= trans_2_io_pipe_phv_out_data_38;
    end else begin
      amplifier_0_3_data_38 <= trans_3_io_pipe_phv_out_data_38;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_39 <= init_io_pipe_phv_out_data_39; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_39 <= trans_2_io_pipe_phv_out_data_39;
    end else begin
      amplifier_0_3_data_39 <= trans_3_io_pipe_phv_out_data_39;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_40 <= init_io_pipe_phv_out_data_40; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_40 <= trans_2_io_pipe_phv_out_data_40;
    end else begin
      amplifier_0_3_data_40 <= trans_3_io_pipe_phv_out_data_40;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_41 <= init_io_pipe_phv_out_data_41; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_41 <= trans_2_io_pipe_phv_out_data_41;
    end else begin
      amplifier_0_3_data_41 <= trans_3_io_pipe_phv_out_data_41;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_42 <= init_io_pipe_phv_out_data_42; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_42 <= trans_2_io_pipe_phv_out_data_42;
    end else begin
      amplifier_0_3_data_42 <= trans_3_io_pipe_phv_out_data_42;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_43 <= init_io_pipe_phv_out_data_43; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_43 <= trans_2_io_pipe_phv_out_data_43;
    end else begin
      amplifier_0_3_data_43 <= trans_3_io_pipe_phv_out_data_43;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_44 <= init_io_pipe_phv_out_data_44; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_44 <= trans_2_io_pipe_phv_out_data_44;
    end else begin
      amplifier_0_3_data_44 <= trans_3_io_pipe_phv_out_data_44;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_45 <= init_io_pipe_phv_out_data_45; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_45 <= trans_2_io_pipe_phv_out_data_45;
    end else begin
      amplifier_0_3_data_45 <= trans_3_io_pipe_phv_out_data_45;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_46 <= init_io_pipe_phv_out_data_46; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_46 <= trans_2_io_pipe_phv_out_data_46;
    end else begin
      amplifier_0_3_data_46 <= trans_3_io_pipe_phv_out_data_46;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_47 <= init_io_pipe_phv_out_data_47; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_47 <= trans_2_io_pipe_phv_out_data_47;
    end else begin
      amplifier_0_3_data_47 <= trans_3_io_pipe_phv_out_data_47;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_48 <= init_io_pipe_phv_out_data_48; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_48 <= trans_2_io_pipe_phv_out_data_48;
    end else begin
      amplifier_0_3_data_48 <= trans_3_io_pipe_phv_out_data_48;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_49 <= init_io_pipe_phv_out_data_49; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_49 <= trans_2_io_pipe_phv_out_data_49;
    end else begin
      amplifier_0_3_data_49 <= trans_3_io_pipe_phv_out_data_49;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_50 <= init_io_pipe_phv_out_data_50; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_50 <= trans_2_io_pipe_phv_out_data_50;
    end else begin
      amplifier_0_3_data_50 <= trans_3_io_pipe_phv_out_data_50;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_51 <= init_io_pipe_phv_out_data_51; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_51 <= trans_2_io_pipe_phv_out_data_51;
    end else begin
      amplifier_0_3_data_51 <= trans_3_io_pipe_phv_out_data_51;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_52 <= init_io_pipe_phv_out_data_52; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_52 <= trans_2_io_pipe_phv_out_data_52;
    end else begin
      amplifier_0_3_data_52 <= trans_3_io_pipe_phv_out_data_52;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_53 <= init_io_pipe_phv_out_data_53; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_53 <= trans_2_io_pipe_phv_out_data_53;
    end else begin
      amplifier_0_3_data_53 <= trans_3_io_pipe_phv_out_data_53;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_54 <= init_io_pipe_phv_out_data_54; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_54 <= trans_2_io_pipe_phv_out_data_54;
    end else begin
      amplifier_0_3_data_54 <= trans_3_io_pipe_phv_out_data_54;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_55 <= init_io_pipe_phv_out_data_55; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_55 <= trans_2_io_pipe_phv_out_data_55;
    end else begin
      amplifier_0_3_data_55 <= trans_3_io_pipe_phv_out_data_55;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_56 <= init_io_pipe_phv_out_data_56; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_56 <= trans_2_io_pipe_phv_out_data_56;
    end else begin
      amplifier_0_3_data_56 <= trans_3_io_pipe_phv_out_data_56;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_57 <= init_io_pipe_phv_out_data_57; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_57 <= trans_2_io_pipe_phv_out_data_57;
    end else begin
      amplifier_0_3_data_57 <= trans_3_io_pipe_phv_out_data_57;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_58 <= init_io_pipe_phv_out_data_58; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_58 <= trans_2_io_pipe_phv_out_data_58;
    end else begin
      amplifier_0_3_data_58 <= trans_3_io_pipe_phv_out_data_58;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_59 <= init_io_pipe_phv_out_data_59; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_59 <= trans_2_io_pipe_phv_out_data_59;
    end else begin
      amplifier_0_3_data_59 <= trans_3_io_pipe_phv_out_data_59;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_60 <= init_io_pipe_phv_out_data_60; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_60 <= trans_2_io_pipe_phv_out_data_60;
    end else begin
      amplifier_0_3_data_60 <= trans_3_io_pipe_phv_out_data_60;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_61 <= init_io_pipe_phv_out_data_61; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_61 <= trans_2_io_pipe_phv_out_data_61;
    end else begin
      amplifier_0_3_data_61 <= trans_3_io_pipe_phv_out_data_61;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_62 <= init_io_pipe_phv_out_data_62; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_62 <= trans_2_io_pipe_phv_out_data_62;
    end else begin
      amplifier_0_3_data_62 <= trans_3_io_pipe_phv_out_data_62;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_63 <= init_io_pipe_phv_out_data_63; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_63 <= trans_2_io_pipe_phv_out_data_63;
    end else begin
      amplifier_0_3_data_63 <= trans_3_io_pipe_phv_out_data_63;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_64 <= init_io_pipe_phv_out_data_64; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_64 <= trans_2_io_pipe_phv_out_data_64;
    end else begin
      amplifier_0_3_data_64 <= trans_3_io_pipe_phv_out_data_64;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_65 <= init_io_pipe_phv_out_data_65; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_65 <= trans_2_io_pipe_phv_out_data_65;
    end else begin
      amplifier_0_3_data_65 <= trans_3_io_pipe_phv_out_data_65;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_66 <= init_io_pipe_phv_out_data_66; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_66 <= trans_2_io_pipe_phv_out_data_66;
    end else begin
      amplifier_0_3_data_66 <= trans_3_io_pipe_phv_out_data_66;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_67 <= init_io_pipe_phv_out_data_67; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_67 <= trans_2_io_pipe_phv_out_data_67;
    end else begin
      amplifier_0_3_data_67 <= trans_3_io_pipe_phv_out_data_67;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_68 <= init_io_pipe_phv_out_data_68; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_68 <= trans_2_io_pipe_phv_out_data_68;
    end else begin
      amplifier_0_3_data_68 <= trans_3_io_pipe_phv_out_data_68;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_69 <= init_io_pipe_phv_out_data_69; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_69 <= trans_2_io_pipe_phv_out_data_69;
    end else begin
      amplifier_0_3_data_69 <= trans_3_io_pipe_phv_out_data_69;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_70 <= init_io_pipe_phv_out_data_70; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_70 <= trans_2_io_pipe_phv_out_data_70;
    end else begin
      amplifier_0_3_data_70 <= trans_3_io_pipe_phv_out_data_70;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_71 <= init_io_pipe_phv_out_data_71; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_71 <= trans_2_io_pipe_phv_out_data_71;
    end else begin
      amplifier_0_3_data_71 <= trans_3_io_pipe_phv_out_data_71;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_72 <= init_io_pipe_phv_out_data_72; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_72 <= trans_2_io_pipe_phv_out_data_72;
    end else begin
      amplifier_0_3_data_72 <= trans_3_io_pipe_phv_out_data_72;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_73 <= init_io_pipe_phv_out_data_73; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_73 <= trans_2_io_pipe_phv_out_data_73;
    end else begin
      amplifier_0_3_data_73 <= trans_3_io_pipe_phv_out_data_73;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_74 <= init_io_pipe_phv_out_data_74; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_74 <= trans_2_io_pipe_phv_out_data_74;
    end else begin
      amplifier_0_3_data_74 <= trans_3_io_pipe_phv_out_data_74;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_75 <= init_io_pipe_phv_out_data_75; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_75 <= trans_2_io_pipe_phv_out_data_75;
    end else begin
      amplifier_0_3_data_75 <= trans_3_io_pipe_phv_out_data_75;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_76 <= init_io_pipe_phv_out_data_76; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_76 <= trans_2_io_pipe_phv_out_data_76;
    end else begin
      amplifier_0_3_data_76 <= trans_3_io_pipe_phv_out_data_76;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_77 <= init_io_pipe_phv_out_data_77; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_77 <= trans_2_io_pipe_phv_out_data_77;
    end else begin
      amplifier_0_3_data_77 <= trans_3_io_pipe_phv_out_data_77;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_78 <= init_io_pipe_phv_out_data_78; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_78 <= trans_2_io_pipe_phv_out_data_78;
    end else begin
      amplifier_0_3_data_78 <= trans_3_io_pipe_phv_out_data_78;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_79 <= init_io_pipe_phv_out_data_79; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_79 <= trans_2_io_pipe_phv_out_data_79;
    end else begin
      amplifier_0_3_data_79 <= trans_3_io_pipe_phv_out_data_79;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_80 <= init_io_pipe_phv_out_data_80; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_80 <= trans_2_io_pipe_phv_out_data_80;
    end else begin
      amplifier_0_3_data_80 <= trans_3_io_pipe_phv_out_data_80;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_81 <= init_io_pipe_phv_out_data_81; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_81 <= trans_2_io_pipe_phv_out_data_81;
    end else begin
      amplifier_0_3_data_81 <= trans_3_io_pipe_phv_out_data_81;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_82 <= init_io_pipe_phv_out_data_82; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_82 <= trans_2_io_pipe_phv_out_data_82;
    end else begin
      amplifier_0_3_data_82 <= trans_3_io_pipe_phv_out_data_82;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_83 <= init_io_pipe_phv_out_data_83; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_83 <= trans_2_io_pipe_phv_out_data_83;
    end else begin
      amplifier_0_3_data_83 <= trans_3_io_pipe_phv_out_data_83;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_84 <= init_io_pipe_phv_out_data_84; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_84 <= trans_2_io_pipe_phv_out_data_84;
    end else begin
      amplifier_0_3_data_84 <= trans_3_io_pipe_phv_out_data_84;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_85 <= init_io_pipe_phv_out_data_85; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_85 <= trans_2_io_pipe_phv_out_data_85;
    end else begin
      amplifier_0_3_data_85 <= trans_3_io_pipe_phv_out_data_85;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_86 <= init_io_pipe_phv_out_data_86; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_86 <= trans_2_io_pipe_phv_out_data_86;
    end else begin
      amplifier_0_3_data_86 <= trans_3_io_pipe_phv_out_data_86;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_87 <= init_io_pipe_phv_out_data_87; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_87 <= trans_2_io_pipe_phv_out_data_87;
    end else begin
      amplifier_0_3_data_87 <= trans_3_io_pipe_phv_out_data_87;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_88 <= init_io_pipe_phv_out_data_88; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_88 <= trans_2_io_pipe_phv_out_data_88;
    end else begin
      amplifier_0_3_data_88 <= trans_3_io_pipe_phv_out_data_88;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_89 <= init_io_pipe_phv_out_data_89; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_89 <= trans_2_io_pipe_phv_out_data_89;
    end else begin
      amplifier_0_3_data_89 <= trans_3_io_pipe_phv_out_data_89;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_90 <= init_io_pipe_phv_out_data_90; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_90 <= trans_2_io_pipe_phv_out_data_90;
    end else begin
      amplifier_0_3_data_90 <= trans_3_io_pipe_phv_out_data_90;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_91 <= init_io_pipe_phv_out_data_91; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_91 <= trans_2_io_pipe_phv_out_data_91;
    end else begin
      amplifier_0_3_data_91 <= trans_3_io_pipe_phv_out_data_91;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_92 <= init_io_pipe_phv_out_data_92; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_92 <= trans_2_io_pipe_phv_out_data_92;
    end else begin
      amplifier_0_3_data_92 <= trans_3_io_pipe_phv_out_data_92;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_93 <= init_io_pipe_phv_out_data_93; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_93 <= trans_2_io_pipe_phv_out_data_93;
    end else begin
      amplifier_0_3_data_93 <= trans_3_io_pipe_phv_out_data_93;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_94 <= init_io_pipe_phv_out_data_94; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_94 <= trans_2_io_pipe_phv_out_data_94;
    end else begin
      amplifier_0_3_data_94 <= trans_3_io_pipe_phv_out_data_94;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_95 <= init_io_pipe_phv_out_data_95; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_95 <= trans_2_io_pipe_phv_out_data_95;
    end else begin
      amplifier_0_3_data_95 <= trans_3_io_pipe_phv_out_data_95;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_96 <= init_io_pipe_phv_out_data_96; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_96 <= trans_2_io_pipe_phv_out_data_96;
    end else begin
      amplifier_0_3_data_96 <= trans_3_io_pipe_phv_out_data_96;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_97 <= init_io_pipe_phv_out_data_97; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_97 <= trans_2_io_pipe_phv_out_data_97;
    end else begin
      amplifier_0_3_data_97 <= trans_3_io_pipe_phv_out_data_97;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_98 <= init_io_pipe_phv_out_data_98; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_98 <= trans_2_io_pipe_phv_out_data_98;
    end else begin
      amplifier_0_3_data_98 <= trans_3_io_pipe_phv_out_data_98;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_99 <= init_io_pipe_phv_out_data_99; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_99 <= trans_2_io_pipe_phv_out_data_99;
    end else begin
      amplifier_0_3_data_99 <= trans_3_io_pipe_phv_out_data_99;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_100 <= init_io_pipe_phv_out_data_100; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_100 <= trans_2_io_pipe_phv_out_data_100;
    end else begin
      amplifier_0_3_data_100 <= trans_3_io_pipe_phv_out_data_100;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_101 <= init_io_pipe_phv_out_data_101; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_101 <= trans_2_io_pipe_phv_out_data_101;
    end else begin
      amplifier_0_3_data_101 <= trans_3_io_pipe_phv_out_data_101;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_102 <= init_io_pipe_phv_out_data_102; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_102 <= trans_2_io_pipe_phv_out_data_102;
    end else begin
      amplifier_0_3_data_102 <= trans_3_io_pipe_phv_out_data_102;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_103 <= init_io_pipe_phv_out_data_103; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_103 <= trans_2_io_pipe_phv_out_data_103;
    end else begin
      amplifier_0_3_data_103 <= trans_3_io_pipe_phv_out_data_103;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_104 <= init_io_pipe_phv_out_data_104; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_104 <= trans_2_io_pipe_phv_out_data_104;
    end else begin
      amplifier_0_3_data_104 <= trans_3_io_pipe_phv_out_data_104;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_105 <= init_io_pipe_phv_out_data_105; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_105 <= trans_2_io_pipe_phv_out_data_105;
    end else begin
      amplifier_0_3_data_105 <= trans_3_io_pipe_phv_out_data_105;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_106 <= init_io_pipe_phv_out_data_106; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_106 <= trans_2_io_pipe_phv_out_data_106;
    end else begin
      amplifier_0_3_data_106 <= trans_3_io_pipe_phv_out_data_106;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_107 <= init_io_pipe_phv_out_data_107; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_107 <= trans_2_io_pipe_phv_out_data_107;
    end else begin
      amplifier_0_3_data_107 <= trans_3_io_pipe_phv_out_data_107;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_108 <= init_io_pipe_phv_out_data_108; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_108 <= trans_2_io_pipe_phv_out_data_108;
    end else begin
      amplifier_0_3_data_108 <= trans_3_io_pipe_phv_out_data_108;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_109 <= init_io_pipe_phv_out_data_109; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_109 <= trans_2_io_pipe_phv_out_data_109;
    end else begin
      amplifier_0_3_data_109 <= trans_3_io_pipe_phv_out_data_109;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_110 <= init_io_pipe_phv_out_data_110; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_110 <= trans_2_io_pipe_phv_out_data_110;
    end else begin
      amplifier_0_3_data_110 <= trans_3_io_pipe_phv_out_data_110;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_111 <= init_io_pipe_phv_out_data_111; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_111 <= trans_2_io_pipe_phv_out_data_111;
    end else begin
      amplifier_0_3_data_111 <= trans_3_io_pipe_phv_out_data_111;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_112 <= init_io_pipe_phv_out_data_112; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_112 <= trans_2_io_pipe_phv_out_data_112;
    end else begin
      amplifier_0_3_data_112 <= trans_3_io_pipe_phv_out_data_112;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_113 <= init_io_pipe_phv_out_data_113; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_113 <= trans_2_io_pipe_phv_out_data_113;
    end else begin
      amplifier_0_3_data_113 <= trans_3_io_pipe_phv_out_data_113;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_114 <= init_io_pipe_phv_out_data_114; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_114 <= trans_2_io_pipe_phv_out_data_114;
    end else begin
      amplifier_0_3_data_114 <= trans_3_io_pipe_phv_out_data_114;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_115 <= init_io_pipe_phv_out_data_115; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_115 <= trans_2_io_pipe_phv_out_data_115;
    end else begin
      amplifier_0_3_data_115 <= trans_3_io_pipe_phv_out_data_115;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_116 <= init_io_pipe_phv_out_data_116; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_116 <= trans_2_io_pipe_phv_out_data_116;
    end else begin
      amplifier_0_3_data_116 <= trans_3_io_pipe_phv_out_data_116;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_117 <= init_io_pipe_phv_out_data_117; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_117 <= trans_2_io_pipe_phv_out_data_117;
    end else begin
      amplifier_0_3_data_117 <= trans_3_io_pipe_phv_out_data_117;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_118 <= init_io_pipe_phv_out_data_118; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_118 <= trans_2_io_pipe_phv_out_data_118;
    end else begin
      amplifier_0_3_data_118 <= trans_3_io_pipe_phv_out_data_118;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_119 <= init_io_pipe_phv_out_data_119; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_119 <= trans_2_io_pipe_phv_out_data_119;
    end else begin
      amplifier_0_3_data_119 <= trans_3_io_pipe_phv_out_data_119;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_120 <= init_io_pipe_phv_out_data_120; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_120 <= trans_2_io_pipe_phv_out_data_120;
    end else begin
      amplifier_0_3_data_120 <= trans_3_io_pipe_phv_out_data_120;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_121 <= init_io_pipe_phv_out_data_121; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_121 <= trans_2_io_pipe_phv_out_data_121;
    end else begin
      amplifier_0_3_data_121 <= trans_3_io_pipe_phv_out_data_121;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_122 <= init_io_pipe_phv_out_data_122; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_122 <= trans_2_io_pipe_phv_out_data_122;
    end else begin
      amplifier_0_3_data_122 <= trans_3_io_pipe_phv_out_data_122;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_123 <= init_io_pipe_phv_out_data_123; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_123 <= trans_2_io_pipe_phv_out_data_123;
    end else begin
      amplifier_0_3_data_123 <= trans_3_io_pipe_phv_out_data_123;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_124 <= init_io_pipe_phv_out_data_124; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_124 <= trans_2_io_pipe_phv_out_data_124;
    end else begin
      amplifier_0_3_data_124 <= trans_3_io_pipe_phv_out_data_124;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_125 <= init_io_pipe_phv_out_data_125; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_125 <= trans_2_io_pipe_phv_out_data_125;
    end else begin
      amplifier_0_3_data_125 <= trans_3_io_pipe_phv_out_data_125;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_126 <= init_io_pipe_phv_out_data_126; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_126 <= trans_2_io_pipe_phv_out_data_126;
    end else begin
      amplifier_0_3_data_126 <= trans_3_io_pipe_phv_out_data_126;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_127 <= init_io_pipe_phv_out_data_127; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_127 <= trans_2_io_pipe_phv_out_data_127;
    end else begin
      amplifier_0_3_data_127 <= trans_3_io_pipe_phv_out_data_127;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_128 <= init_io_pipe_phv_out_data_128; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_128 <= trans_2_io_pipe_phv_out_data_128;
    end else begin
      amplifier_0_3_data_128 <= trans_3_io_pipe_phv_out_data_128;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_129 <= init_io_pipe_phv_out_data_129; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_129 <= trans_2_io_pipe_phv_out_data_129;
    end else begin
      amplifier_0_3_data_129 <= trans_3_io_pipe_phv_out_data_129;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_130 <= init_io_pipe_phv_out_data_130; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_130 <= trans_2_io_pipe_phv_out_data_130;
    end else begin
      amplifier_0_3_data_130 <= trans_3_io_pipe_phv_out_data_130;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_131 <= init_io_pipe_phv_out_data_131; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_131 <= trans_2_io_pipe_phv_out_data_131;
    end else begin
      amplifier_0_3_data_131 <= trans_3_io_pipe_phv_out_data_131;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_132 <= init_io_pipe_phv_out_data_132; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_132 <= trans_2_io_pipe_phv_out_data_132;
    end else begin
      amplifier_0_3_data_132 <= trans_3_io_pipe_phv_out_data_132;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_133 <= init_io_pipe_phv_out_data_133; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_133 <= trans_2_io_pipe_phv_out_data_133;
    end else begin
      amplifier_0_3_data_133 <= trans_3_io_pipe_phv_out_data_133;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_134 <= init_io_pipe_phv_out_data_134; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_134 <= trans_2_io_pipe_phv_out_data_134;
    end else begin
      amplifier_0_3_data_134 <= trans_3_io_pipe_phv_out_data_134;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_135 <= init_io_pipe_phv_out_data_135; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_135 <= trans_2_io_pipe_phv_out_data_135;
    end else begin
      amplifier_0_3_data_135 <= trans_3_io_pipe_phv_out_data_135;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_136 <= init_io_pipe_phv_out_data_136; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_136 <= trans_2_io_pipe_phv_out_data_136;
    end else begin
      amplifier_0_3_data_136 <= trans_3_io_pipe_phv_out_data_136;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_137 <= init_io_pipe_phv_out_data_137; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_137 <= trans_2_io_pipe_phv_out_data_137;
    end else begin
      amplifier_0_3_data_137 <= trans_3_io_pipe_phv_out_data_137;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_138 <= init_io_pipe_phv_out_data_138; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_138 <= trans_2_io_pipe_phv_out_data_138;
    end else begin
      amplifier_0_3_data_138 <= trans_3_io_pipe_phv_out_data_138;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_139 <= init_io_pipe_phv_out_data_139; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_139 <= trans_2_io_pipe_phv_out_data_139;
    end else begin
      amplifier_0_3_data_139 <= trans_3_io_pipe_phv_out_data_139;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_140 <= init_io_pipe_phv_out_data_140; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_140 <= trans_2_io_pipe_phv_out_data_140;
    end else begin
      amplifier_0_3_data_140 <= trans_3_io_pipe_phv_out_data_140;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_141 <= init_io_pipe_phv_out_data_141; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_141 <= trans_2_io_pipe_phv_out_data_141;
    end else begin
      amplifier_0_3_data_141 <= trans_3_io_pipe_phv_out_data_141;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_142 <= init_io_pipe_phv_out_data_142; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_142 <= trans_2_io_pipe_phv_out_data_142;
    end else begin
      amplifier_0_3_data_142 <= trans_3_io_pipe_phv_out_data_142;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_143 <= init_io_pipe_phv_out_data_143; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_143 <= trans_2_io_pipe_phv_out_data_143;
    end else begin
      amplifier_0_3_data_143 <= trans_3_io_pipe_phv_out_data_143;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_144 <= init_io_pipe_phv_out_data_144; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_144 <= trans_2_io_pipe_phv_out_data_144;
    end else begin
      amplifier_0_3_data_144 <= trans_3_io_pipe_phv_out_data_144;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_145 <= init_io_pipe_phv_out_data_145; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_145 <= trans_2_io_pipe_phv_out_data_145;
    end else begin
      amplifier_0_3_data_145 <= trans_3_io_pipe_phv_out_data_145;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_146 <= init_io_pipe_phv_out_data_146; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_146 <= trans_2_io_pipe_phv_out_data_146;
    end else begin
      amplifier_0_3_data_146 <= trans_3_io_pipe_phv_out_data_146;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_147 <= init_io_pipe_phv_out_data_147; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_147 <= trans_2_io_pipe_phv_out_data_147;
    end else begin
      amplifier_0_3_data_147 <= trans_3_io_pipe_phv_out_data_147;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_148 <= init_io_pipe_phv_out_data_148; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_148 <= trans_2_io_pipe_phv_out_data_148;
    end else begin
      amplifier_0_3_data_148 <= trans_3_io_pipe_phv_out_data_148;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_149 <= init_io_pipe_phv_out_data_149; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_149 <= trans_2_io_pipe_phv_out_data_149;
    end else begin
      amplifier_0_3_data_149 <= trans_3_io_pipe_phv_out_data_149;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_150 <= init_io_pipe_phv_out_data_150; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_150 <= trans_2_io_pipe_phv_out_data_150;
    end else begin
      amplifier_0_3_data_150 <= trans_3_io_pipe_phv_out_data_150;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_151 <= init_io_pipe_phv_out_data_151; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_151 <= trans_2_io_pipe_phv_out_data_151;
    end else begin
      amplifier_0_3_data_151 <= trans_3_io_pipe_phv_out_data_151;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_152 <= init_io_pipe_phv_out_data_152; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_152 <= trans_2_io_pipe_phv_out_data_152;
    end else begin
      amplifier_0_3_data_152 <= trans_3_io_pipe_phv_out_data_152;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_153 <= init_io_pipe_phv_out_data_153; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_153 <= trans_2_io_pipe_phv_out_data_153;
    end else begin
      amplifier_0_3_data_153 <= trans_3_io_pipe_phv_out_data_153;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_154 <= init_io_pipe_phv_out_data_154; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_154 <= trans_2_io_pipe_phv_out_data_154;
    end else begin
      amplifier_0_3_data_154 <= trans_3_io_pipe_phv_out_data_154;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_155 <= init_io_pipe_phv_out_data_155; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_155 <= trans_2_io_pipe_phv_out_data_155;
    end else begin
      amplifier_0_3_data_155 <= trans_3_io_pipe_phv_out_data_155;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_156 <= init_io_pipe_phv_out_data_156; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_156 <= trans_2_io_pipe_phv_out_data_156;
    end else begin
      amplifier_0_3_data_156 <= trans_3_io_pipe_phv_out_data_156;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_157 <= init_io_pipe_phv_out_data_157; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_157 <= trans_2_io_pipe_phv_out_data_157;
    end else begin
      amplifier_0_3_data_157 <= trans_3_io_pipe_phv_out_data_157;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_158 <= init_io_pipe_phv_out_data_158; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_158 <= trans_2_io_pipe_phv_out_data_158;
    end else begin
      amplifier_0_3_data_158 <= trans_3_io_pipe_phv_out_data_158;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_159 <= init_io_pipe_phv_out_data_159; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_159 <= trans_2_io_pipe_phv_out_data_159;
    end else begin
      amplifier_0_3_data_159 <= trans_3_io_pipe_phv_out_data_159;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_160 <= init_io_pipe_phv_out_data_160; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_160 <= trans_2_io_pipe_phv_out_data_160;
    end else begin
      amplifier_0_3_data_160 <= trans_3_io_pipe_phv_out_data_160;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_161 <= init_io_pipe_phv_out_data_161; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_161 <= trans_2_io_pipe_phv_out_data_161;
    end else begin
      amplifier_0_3_data_161 <= trans_3_io_pipe_phv_out_data_161;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_162 <= init_io_pipe_phv_out_data_162; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_162 <= trans_2_io_pipe_phv_out_data_162;
    end else begin
      amplifier_0_3_data_162 <= trans_3_io_pipe_phv_out_data_162;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_163 <= init_io_pipe_phv_out_data_163; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_163 <= trans_2_io_pipe_phv_out_data_163;
    end else begin
      amplifier_0_3_data_163 <= trans_3_io_pipe_phv_out_data_163;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_164 <= init_io_pipe_phv_out_data_164; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_164 <= trans_2_io_pipe_phv_out_data_164;
    end else begin
      amplifier_0_3_data_164 <= trans_3_io_pipe_phv_out_data_164;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_165 <= init_io_pipe_phv_out_data_165; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_165 <= trans_2_io_pipe_phv_out_data_165;
    end else begin
      amplifier_0_3_data_165 <= trans_3_io_pipe_phv_out_data_165;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_166 <= init_io_pipe_phv_out_data_166; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_166 <= trans_2_io_pipe_phv_out_data_166;
    end else begin
      amplifier_0_3_data_166 <= trans_3_io_pipe_phv_out_data_166;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_167 <= init_io_pipe_phv_out_data_167; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_167 <= trans_2_io_pipe_phv_out_data_167;
    end else begin
      amplifier_0_3_data_167 <= trans_3_io_pipe_phv_out_data_167;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_168 <= init_io_pipe_phv_out_data_168; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_168 <= trans_2_io_pipe_phv_out_data_168;
    end else begin
      amplifier_0_3_data_168 <= trans_3_io_pipe_phv_out_data_168;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_169 <= init_io_pipe_phv_out_data_169; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_169 <= trans_2_io_pipe_phv_out_data_169;
    end else begin
      amplifier_0_3_data_169 <= trans_3_io_pipe_phv_out_data_169;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_170 <= init_io_pipe_phv_out_data_170; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_170 <= trans_2_io_pipe_phv_out_data_170;
    end else begin
      amplifier_0_3_data_170 <= trans_3_io_pipe_phv_out_data_170;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_171 <= init_io_pipe_phv_out_data_171; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_171 <= trans_2_io_pipe_phv_out_data_171;
    end else begin
      amplifier_0_3_data_171 <= trans_3_io_pipe_phv_out_data_171;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_172 <= init_io_pipe_phv_out_data_172; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_172 <= trans_2_io_pipe_phv_out_data_172;
    end else begin
      amplifier_0_3_data_172 <= trans_3_io_pipe_phv_out_data_172;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_173 <= init_io_pipe_phv_out_data_173; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_173 <= trans_2_io_pipe_phv_out_data_173;
    end else begin
      amplifier_0_3_data_173 <= trans_3_io_pipe_phv_out_data_173;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_174 <= init_io_pipe_phv_out_data_174; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_174 <= trans_2_io_pipe_phv_out_data_174;
    end else begin
      amplifier_0_3_data_174 <= trans_3_io_pipe_phv_out_data_174;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_175 <= init_io_pipe_phv_out_data_175; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_175 <= trans_2_io_pipe_phv_out_data_175;
    end else begin
      amplifier_0_3_data_175 <= trans_3_io_pipe_phv_out_data_175;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_176 <= init_io_pipe_phv_out_data_176; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_176 <= trans_2_io_pipe_phv_out_data_176;
    end else begin
      amplifier_0_3_data_176 <= trans_3_io_pipe_phv_out_data_176;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_177 <= init_io_pipe_phv_out_data_177; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_177 <= trans_2_io_pipe_phv_out_data_177;
    end else begin
      amplifier_0_3_data_177 <= trans_3_io_pipe_phv_out_data_177;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_178 <= init_io_pipe_phv_out_data_178; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_178 <= trans_2_io_pipe_phv_out_data_178;
    end else begin
      amplifier_0_3_data_178 <= trans_3_io_pipe_phv_out_data_178;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_179 <= init_io_pipe_phv_out_data_179; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_179 <= trans_2_io_pipe_phv_out_data_179;
    end else begin
      amplifier_0_3_data_179 <= trans_3_io_pipe_phv_out_data_179;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_180 <= init_io_pipe_phv_out_data_180; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_180 <= trans_2_io_pipe_phv_out_data_180;
    end else begin
      amplifier_0_3_data_180 <= trans_3_io_pipe_phv_out_data_180;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_181 <= init_io_pipe_phv_out_data_181; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_181 <= trans_2_io_pipe_phv_out_data_181;
    end else begin
      amplifier_0_3_data_181 <= trans_3_io_pipe_phv_out_data_181;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_182 <= init_io_pipe_phv_out_data_182; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_182 <= trans_2_io_pipe_phv_out_data_182;
    end else begin
      amplifier_0_3_data_182 <= trans_3_io_pipe_phv_out_data_182;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_183 <= init_io_pipe_phv_out_data_183; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_183 <= trans_2_io_pipe_phv_out_data_183;
    end else begin
      amplifier_0_3_data_183 <= trans_3_io_pipe_phv_out_data_183;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_184 <= init_io_pipe_phv_out_data_184; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_184 <= trans_2_io_pipe_phv_out_data_184;
    end else begin
      amplifier_0_3_data_184 <= trans_3_io_pipe_phv_out_data_184;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_185 <= init_io_pipe_phv_out_data_185; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_185 <= trans_2_io_pipe_phv_out_data_185;
    end else begin
      amplifier_0_3_data_185 <= trans_3_io_pipe_phv_out_data_185;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_186 <= init_io_pipe_phv_out_data_186; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_186 <= trans_2_io_pipe_phv_out_data_186;
    end else begin
      amplifier_0_3_data_186 <= trans_3_io_pipe_phv_out_data_186;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_187 <= init_io_pipe_phv_out_data_187; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_187 <= trans_2_io_pipe_phv_out_data_187;
    end else begin
      amplifier_0_3_data_187 <= trans_3_io_pipe_phv_out_data_187;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_188 <= init_io_pipe_phv_out_data_188; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_188 <= trans_2_io_pipe_phv_out_data_188;
    end else begin
      amplifier_0_3_data_188 <= trans_3_io_pipe_phv_out_data_188;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_189 <= init_io_pipe_phv_out_data_189; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_189 <= trans_2_io_pipe_phv_out_data_189;
    end else begin
      amplifier_0_3_data_189 <= trans_3_io_pipe_phv_out_data_189;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_190 <= init_io_pipe_phv_out_data_190; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_190 <= trans_2_io_pipe_phv_out_data_190;
    end else begin
      amplifier_0_3_data_190 <= trans_3_io_pipe_phv_out_data_190;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_191 <= init_io_pipe_phv_out_data_191; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_191 <= trans_2_io_pipe_phv_out_data_191;
    end else begin
      amplifier_0_3_data_191 <= trans_3_io_pipe_phv_out_data_191;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_192 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_192 <= trans_2_io_pipe_phv_out_data_192;
    end else begin
      amplifier_0_3_data_192 <= trans_3_io_pipe_phv_out_data_192;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_193 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_193 <= trans_2_io_pipe_phv_out_data_193;
    end else begin
      amplifier_0_3_data_193 <= trans_3_io_pipe_phv_out_data_193;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_194 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_194 <= trans_2_io_pipe_phv_out_data_194;
    end else begin
      amplifier_0_3_data_194 <= trans_3_io_pipe_phv_out_data_194;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_195 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_195 <= trans_2_io_pipe_phv_out_data_195;
    end else begin
      amplifier_0_3_data_195 <= trans_3_io_pipe_phv_out_data_195;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_196 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_196 <= trans_2_io_pipe_phv_out_data_196;
    end else begin
      amplifier_0_3_data_196 <= trans_3_io_pipe_phv_out_data_196;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_197 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_197 <= trans_2_io_pipe_phv_out_data_197;
    end else begin
      amplifier_0_3_data_197 <= trans_3_io_pipe_phv_out_data_197;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_198 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_198 <= trans_2_io_pipe_phv_out_data_198;
    end else begin
      amplifier_0_3_data_198 <= trans_3_io_pipe_phv_out_data_198;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_199 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_199 <= trans_2_io_pipe_phv_out_data_199;
    end else begin
      amplifier_0_3_data_199 <= trans_3_io_pipe_phv_out_data_199;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_200 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_200 <= trans_2_io_pipe_phv_out_data_200;
    end else begin
      amplifier_0_3_data_200 <= trans_3_io_pipe_phv_out_data_200;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_201 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_201 <= trans_2_io_pipe_phv_out_data_201;
    end else begin
      amplifier_0_3_data_201 <= trans_3_io_pipe_phv_out_data_201;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_202 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_202 <= trans_2_io_pipe_phv_out_data_202;
    end else begin
      amplifier_0_3_data_202 <= trans_3_io_pipe_phv_out_data_202;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_203 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_203 <= trans_2_io_pipe_phv_out_data_203;
    end else begin
      amplifier_0_3_data_203 <= trans_3_io_pipe_phv_out_data_203;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_204 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_204 <= trans_2_io_pipe_phv_out_data_204;
    end else begin
      amplifier_0_3_data_204 <= trans_3_io_pipe_phv_out_data_204;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_205 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_205 <= trans_2_io_pipe_phv_out_data_205;
    end else begin
      amplifier_0_3_data_205 <= trans_3_io_pipe_phv_out_data_205;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_206 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_206 <= trans_2_io_pipe_phv_out_data_206;
    end else begin
      amplifier_0_3_data_206 <= trans_3_io_pipe_phv_out_data_206;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_207 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_207 <= trans_2_io_pipe_phv_out_data_207;
    end else begin
      amplifier_0_3_data_207 <= trans_3_io_pipe_phv_out_data_207;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_208 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_208 <= trans_2_io_pipe_phv_out_data_208;
    end else begin
      amplifier_0_3_data_208 <= trans_3_io_pipe_phv_out_data_208;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_209 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_209 <= trans_2_io_pipe_phv_out_data_209;
    end else begin
      amplifier_0_3_data_209 <= trans_3_io_pipe_phv_out_data_209;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_210 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_210 <= trans_2_io_pipe_phv_out_data_210;
    end else begin
      amplifier_0_3_data_210 <= trans_3_io_pipe_phv_out_data_210;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_211 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_211 <= trans_2_io_pipe_phv_out_data_211;
    end else begin
      amplifier_0_3_data_211 <= trans_3_io_pipe_phv_out_data_211;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_212 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_212 <= trans_2_io_pipe_phv_out_data_212;
    end else begin
      amplifier_0_3_data_212 <= trans_3_io_pipe_phv_out_data_212;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_213 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_213 <= trans_2_io_pipe_phv_out_data_213;
    end else begin
      amplifier_0_3_data_213 <= trans_3_io_pipe_phv_out_data_213;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_214 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_214 <= trans_2_io_pipe_phv_out_data_214;
    end else begin
      amplifier_0_3_data_214 <= trans_3_io_pipe_phv_out_data_214;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_215 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_215 <= trans_2_io_pipe_phv_out_data_215;
    end else begin
      amplifier_0_3_data_215 <= trans_3_io_pipe_phv_out_data_215;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_216 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_216 <= trans_2_io_pipe_phv_out_data_216;
    end else begin
      amplifier_0_3_data_216 <= trans_3_io_pipe_phv_out_data_216;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_217 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_217 <= trans_2_io_pipe_phv_out_data_217;
    end else begin
      amplifier_0_3_data_217 <= trans_3_io_pipe_phv_out_data_217;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_218 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_218 <= trans_2_io_pipe_phv_out_data_218;
    end else begin
      amplifier_0_3_data_218 <= trans_3_io_pipe_phv_out_data_218;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_219 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_219 <= trans_2_io_pipe_phv_out_data_219;
    end else begin
      amplifier_0_3_data_219 <= trans_3_io_pipe_phv_out_data_219;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_220 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_220 <= trans_2_io_pipe_phv_out_data_220;
    end else begin
      amplifier_0_3_data_220 <= trans_3_io_pipe_phv_out_data_220;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_221 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_221 <= trans_2_io_pipe_phv_out_data_221;
    end else begin
      amplifier_0_3_data_221 <= trans_3_io_pipe_phv_out_data_221;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_222 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_222 <= trans_2_io_pipe_phv_out_data_222;
    end else begin
      amplifier_0_3_data_222 <= trans_3_io_pipe_phv_out_data_222;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_223 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_223 <= trans_2_io_pipe_phv_out_data_223;
    end else begin
      amplifier_0_3_data_223 <= trans_3_io_pipe_phv_out_data_223;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_224 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_224 <= trans_2_io_pipe_phv_out_data_224;
    end else begin
      amplifier_0_3_data_224 <= trans_3_io_pipe_phv_out_data_224;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_225 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_225 <= trans_2_io_pipe_phv_out_data_225;
    end else begin
      amplifier_0_3_data_225 <= trans_3_io_pipe_phv_out_data_225;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_226 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_226 <= trans_2_io_pipe_phv_out_data_226;
    end else begin
      amplifier_0_3_data_226 <= trans_3_io_pipe_phv_out_data_226;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_227 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_227 <= trans_2_io_pipe_phv_out_data_227;
    end else begin
      amplifier_0_3_data_227 <= trans_3_io_pipe_phv_out_data_227;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_228 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_228 <= trans_2_io_pipe_phv_out_data_228;
    end else begin
      amplifier_0_3_data_228 <= trans_3_io_pipe_phv_out_data_228;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_229 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_229 <= trans_2_io_pipe_phv_out_data_229;
    end else begin
      amplifier_0_3_data_229 <= trans_3_io_pipe_phv_out_data_229;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_230 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_230 <= trans_2_io_pipe_phv_out_data_230;
    end else begin
      amplifier_0_3_data_230 <= trans_3_io_pipe_phv_out_data_230;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_231 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_231 <= trans_2_io_pipe_phv_out_data_231;
    end else begin
      amplifier_0_3_data_231 <= trans_3_io_pipe_phv_out_data_231;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_232 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_232 <= trans_2_io_pipe_phv_out_data_232;
    end else begin
      amplifier_0_3_data_232 <= trans_3_io_pipe_phv_out_data_232;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_233 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_233 <= trans_2_io_pipe_phv_out_data_233;
    end else begin
      amplifier_0_3_data_233 <= trans_3_io_pipe_phv_out_data_233;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_234 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_234 <= trans_2_io_pipe_phv_out_data_234;
    end else begin
      amplifier_0_3_data_234 <= trans_3_io_pipe_phv_out_data_234;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_235 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_235 <= trans_2_io_pipe_phv_out_data_235;
    end else begin
      amplifier_0_3_data_235 <= trans_3_io_pipe_phv_out_data_235;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_236 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_236 <= trans_2_io_pipe_phv_out_data_236;
    end else begin
      amplifier_0_3_data_236 <= trans_3_io_pipe_phv_out_data_236;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_237 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_237 <= trans_2_io_pipe_phv_out_data_237;
    end else begin
      amplifier_0_3_data_237 <= trans_3_io_pipe_phv_out_data_237;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_238 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_238 <= trans_2_io_pipe_phv_out_data_238;
    end else begin
      amplifier_0_3_data_238 <= trans_3_io_pipe_phv_out_data_238;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_239 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_239 <= trans_2_io_pipe_phv_out_data_239;
    end else begin
      amplifier_0_3_data_239 <= trans_3_io_pipe_phv_out_data_239;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_240 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_240 <= trans_2_io_pipe_phv_out_data_240;
    end else begin
      amplifier_0_3_data_240 <= trans_3_io_pipe_phv_out_data_240;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_241 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_241 <= trans_2_io_pipe_phv_out_data_241;
    end else begin
      amplifier_0_3_data_241 <= trans_3_io_pipe_phv_out_data_241;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_242 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_242 <= trans_2_io_pipe_phv_out_data_242;
    end else begin
      amplifier_0_3_data_242 <= trans_3_io_pipe_phv_out_data_242;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_243 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_243 <= trans_2_io_pipe_phv_out_data_243;
    end else begin
      amplifier_0_3_data_243 <= trans_3_io_pipe_phv_out_data_243;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_244 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_244 <= trans_2_io_pipe_phv_out_data_244;
    end else begin
      amplifier_0_3_data_244 <= trans_3_io_pipe_phv_out_data_244;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_245 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_245 <= trans_2_io_pipe_phv_out_data_245;
    end else begin
      amplifier_0_3_data_245 <= trans_3_io_pipe_phv_out_data_245;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_246 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_246 <= trans_2_io_pipe_phv_out_data_246;
    end else begin
      amplifier_0_3_data_246 <= trans_3_io_pipe_phv_out_data_246;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_247 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_247 <= trans_2_io_pipe_phv_out_data_247;
    end else begin
      amplifier_0_3_data_247 <= trans_3_io_pipe_phv_out_data_247;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_248 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_248 <= trans_2_io_pipe_phv_out_data_248;
    end else begin
      amplifier_0_3_data_248 <= trans_3_io_pipe_phv_out_data_248;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_249 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_249 <= trans_2_io_pipe_phv_out_data_249;
    end else begin
      amplifier_0_3_data_249 <= trans_3_io_pipe_phv_out_data_249;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_250 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_250 <= trans_2_io_pipe_phv_out_data_250;
    end else begin
      amplifier_0_3_data_250 <= trans_3_io_pipe_phv_out_data_250;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_251 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_251 <= trans_2_io_pipe_phv_out_data_251;
    end else begin
      amplifier_0_3_data_251 <= trans_3_io_pipe_phv_out_data_251;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_252 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_252 <= trans_2_io_pipe_phv_out_data_252;
    end else begin
      amplifier_0_3_data_252 <= trans_3_io_pipe_phv_out_data_252;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_253 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_253 <= trans_2_io_pipe_phv_out_data_253;
    end else begin
      amplifier_0_3_data_253 <= trans_3_io_pipe_phv_out_data_253;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_254 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_254 <= trans_2_io_pipe_phv_out_data_254;
    end else begin
      amplifier_0_3_data_254 <= trans_3_io_pipe_phv_out_data_254;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_data_255 <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_data_255 <= trans_2_io_pipe_phv_out_data_255;
    end else begin
      amplifier_0_3_data_255 <= trans_3_io_pipe_phv_out_data_255;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_header_0 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_header_0 <= trans_2_io_pipe_phv_out_header_0;
    end else begin
      amplifier_0_3_header_0 <= trans_3_io_pipe_phv_out_header_0;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_header_1 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_header_1 <= trans_2_io_pipe_phv_out_header_1;
    end else begin
      amplifier_0_3_header_1 <= trans_3_io_pipe_phv_out_header_1;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_header_2 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_header_2 <= trans_2_io_pipe_phv_out_header_2;
    end else begin
      amplifier_0_3_header_2 <= trans_3_io_pipe_phv_out_header_2;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_header_3 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_header_3 <= trans_2_io_pipe_phv_out_header_3;
    end else begin
      amplifier_0_3_header_3 <= trans_3_io_pipe_phv_out_header_3;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_header_4 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_header_4 <= trans_2_io_pipe_phv_out_header_4;
    end else begin
      amplifier_0_3_header_4 <= trans_3_io_pipe_phv_out_header_4;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_header_5 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_header_5 <= trans_2_io_pipe_phv_out_header_5;
    end else begin
      amplifier_0_3_header_5 <= trans_3_io_pipe_phv_out_header_5;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_header_6 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_header_6 <= trans_2_io_pipe_phv_out_header_6;
    end else begin
      amplifier_0_3_header_6 <= trans_3_io_pipe_phv_out_header_6;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_header_7 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_header_7 <= trans_2_io_pipe_phv_out_header_7;
    end else begin
      amplifier_0_3_header_7 <= trans_3_io_pipe_phv_out_header_7;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_header_8 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_header_8 <= trans_2_io_pipe_phv_out_header_8;
    end else begin
      amplifier_0_3_header_8 <= trans_3_io_pipe_phv_out_header_8;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_header_9 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_header_9 <= trans_2_io_pipe_phv_out_header_9;
    end else begin
      amplifier_0_3_header_9 <= trans_3_io_pipe_phv_out_header_9;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_header_10 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_header_10 <= trans_2_io_pipe_phv_out_header_10;
    end else begin
      amplifier_0_3_header_10 <= trans_3_io_pipe_phv_out_header_10;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_header_11 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_header_11 <= trans_2_io_pipe_phv_out_header_11;
    end else begin
      amplifier_0_3_header_11 <= trans_3_io_pipe_phv_out_header_11;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_header_12 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_header_12 <= trans_2_io_pipe_phv_out_header_12;
    end else begin
      amplifier_0_3_header_12 <= trans_3_io_pipe_phv_out_header_12;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_header_13 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_header_13 <= trans_2_io_pipe_phv_out_header_13;
    end else begin
      amplifier_0_3_header_13 <= trans_3_io_pipe_phv_out_header_13;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_header_14 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_header_14 <= trans_2_io_pipe_phv_out_header_14;
    end else begin
      amplifier_0_3_header_14 <= trans_3_io_pipe_phv_out_header_14;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_header_15 <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_header_15 <= trans_2_io_pipe_phv_out_header_15;
    end else begin
      amplifier_0_3_header_15 <= trans_3_io_pipe_phv_out_header_15;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_parse_current_state <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_parse_current_state <= trans_2_io_pipe_phv_out_parse_current_state;
    end else begin
      amplifier_0_3_parse_current_state <= trans_3_io_pipe_phv_out_parse_current_state;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_parse_current_offset <= 8'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_parse_current_offset <= trans_2_io_pipe_phv_out_parse_current_offset;
    end else begin
      amplifier_0_3_parse_current_offset <= trans_3_io_pipe_phv_out_parse_current_offset;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_parse_transition_field <= 16'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_parse_transition_field <= trans_2_io_pipe_phv_out_parse_transition_field;
    end else begin
      amplifier_0_3_parse_transition_field <= trans_3_io_pipe_phv_out_parse_transition_field;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_next_processor_id <= init_io_pipe_phv_out_next_processor_id; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_next_processor_id <= trans_2_io_pipe_phv_out_next_processor_id;
    end else begin
      amplifier_0_3_next_processor_id <= trans_3_io_pipe_phv_out_next_processor_id;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_next_config_id <= 1'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_next_config_id <= trans_2_io_pipe_phv_out_next_config_id;
    end else begin
      amplifier_0_3_next_config_id <= trans_3_io_pipe_phv_out_next_config_id;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      amplifier_0_3_is_valid_processor <= 1'h0; // @[ipsa.scala 127:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 116:31]
      amplifier_0_3_is_valid_processor <= trans_2_io_pipe_phv_out_is_valid_processor;
    end else begin
      amplifier_0_3_is_valid_processor <= trans_3_io_pipe_phv_out_is_valid_processor;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_0 <= amplifier_0_2_data_0;
    end else begin
      amplifier_1_0_data_0 <= amplifier_0_0_data_0;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_1 <= amplifier_0_2_data_1;
    end else begin
      amplifier_1_0_data_1 <= amplifier_0_0_data_1;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_2 <= amplifier_0_2_data_2;
    end else begin
      amplifier_1_0_data_2 <= amplifier_0_0_data_2;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_3 <= amplifier_0_2_data_3;
    end else begin
      amplifier_1_0_data_3 <= amplifier_0_0_data_3;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_4 <= amplifier_0_2_data_4;
    end else begin
      amplifier_1_0_data_4 <= amplifier_0_0_data_4;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_5 <= amplifier_0_2_data_5;
    end else begin
      amplifier_1_0_data_5 <= amplifier_0_0_data_5;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_6 <= amplifier_0_2_data_6;
    end else begin
      amplifier_1_0_data_6 <= amplifier_0_0_data_6;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_7 <= amplifier_0_2_data_7;
    end else begin
      amplifier_1_0_data_7 <= amplifier_0_0_data_7;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_8 <= amplifier_0_2_data_8;
    end else begin
      amplifier_1_0_data_8 <= amplifier_0_0_data_8;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_9 <= amplifier_0_2_data_9;
    end else begin
      amplifier_1_0_data_9 <= amplifier_0_0_data_9;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_10 <= amplifier_0_2_data_10;
    end else begin
      amplifier_1_0_data_10 <= amplifier_0_0_data_10;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_11 <= amplifier_0_2_data_11;
    end else begin
      amplifier_1_0_data_11 <= amplifier_0_0_data_11;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_12 <= amplifier_0_2_data_12;
    end else begin
      amplifier_1_0_data_12 <= amplifier_0_0_data_12;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_13 <= amplifier_0_2_data_13;
    end else begin
      amplifier_1_0_data_13 <= amplifier_0_0_data_13;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_14 <= amplifier_0_2_data_14;
    end else begin
      amplifier_1_0_data_14 <= amplifier_0_0_data_14;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_15 <= amplifier_0_2_data_15;
    end else begin
      amplifier_1_0_data_15 <= amplifier_0_0_data_15;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_16 <= amplifier_0_2_data_16;
    end else begin
      amplifier_1_0_data_16 <= amplifier_0_0_data_16;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_17 <= amplifier_0_2_data_17;
    end else begin
      amplifier_1_0_data_17 <= amplifier_0_0_data_17;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_18 <= amplifier_0_2_data_18;
    end else begin
      amplifier_1_0_data_18 <= amplifier_0_0_data_18;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_19 <= amplifier_0_2_data_19;
    end else begin
      amplifier_1_0_data_19 <= amplifier_0_0_data_19;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_20 <= amplifier_0_2_data_20;
    end else begin
      amplifier_1_0_data_20 <= amplifier_0_0_data_20;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_21 <= amplifier_0_2_data_21;
    end else begin
      amplifier_1_0_data_21 <= amplifier_0_0_data_21;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_22 <= amplifier_0_2_data_22;
    end else begin
      amplifier_1_0_data_22 <= amplifier_0_0_data_22;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_23 <= amplifier_0_2_data_23;
    end else begin
      amplifier_1_0_data_23 <= amplifier_0_0_data_23;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_24 <= amplifier_0_2_data_24;
    end else begin
      amplifier_1_0_data_24 <= amplifier_0_0_data_24;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_25 <= amplifier_0_2_data_25;
    end else begin
      amplifier_1_0_data_25 <= amplifier_0_0_data_25;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_26 <= amplifier_0_2_data_26;
    end else begin
      amplifier_1_0_data_26 <= amplifier_0_0_data_26;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_27 <= amplifier_0_2_data_27;
    end else begin
      amplifier_1_0_data_27 <= amplifier_0_0_data_27;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_28 <= amplifier_0_2_data_28;
    end else begin
      amplifier_1_0_data_28 <= amplifier_0_0_data_28;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_29 <= amplifier_0_2_data_29;
    end else begin
      amplifier_1_0_data_29 <= amplifier_0_0_data_29;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_30 <= amplifier_0_2_data_30;
    end else begin
      amplifier_1_0_data_30 <= amplifier_0_0_data_30;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_31 <= amplifier_0_2_data_31;
    end else begin
      amplifier_1_0_data_31 <= amplifier_0_0_data_31;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_32 <= amplifier_0_2_data_32;
    end else begin
      amplifier_1_0_data_32 <= amplifier_0_0_data_32;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_33 <= amplifier_0_2_data_33;
    end else begin
      amplifier_1_0_data_33 <= amplifier_0_0_data_33;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_34 <= amplifier_0_2_data_34;
    end else begin
      amplifier_1_0_data_34 <= amplifier_0_0_data_34;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_35 <= amplifier_0_2_data_35;
    end else begin
      amplifier_1_0_data_35 <= amplifier_0_0_data_35;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_36 <= amplifier_0_2_data_36;
    end else begin
      amplifier_1_0_data_36 <= amplifier_0_0_data_36;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_37 <= amplifier_0_2_data_37;
    end else begin
      amplifier_1_0_data_37 <= amplifier_0_0_data_37;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_38 <= amplifier_0_2_data_38;
    end else begin
      amplifier_1_0_data_38 <= amplifier_0_0_data_38;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_39 <= amplifier_0_2_data_39;
    end else begin
      amplifier_1_0_data_39 <= amplifier_0_0_data_39;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_40 <= amplifier_0_2_data_40;
    end else begin
      amplifier_1_0_data_40 <= amplifier_0_0_data_40;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_41 <= amplifier_0_2_data_41;
    end else begin
      amplifier_1_0_data_41 <= amplifier_0_0_data_41;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_42 <= amplifier_0_2_data_42;
    end else begin
      amplifier_1_0_data_42 <= amplifier_0_0_data_42;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_43 <= amplifier_0_2_data_43;
    end else begin
      amplifier_1_0_data_43 <= amplifier_0_0_data_43;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_44 <= amplifier_0_2_data_44;
    end else begin
      amplifier_1_0_data_44 <= amplifier_0_0_data_44;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_45 <= amplifier_0_2_data_45;
    end else begin
      amplifier_1_0_data_45 <= amplifier_0_0_data_45;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_46 <= amplifier_0_2_data_46;
    end else begin
      amplifier_1_0_data_46 <= amplifier_0_0_data_46;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_47 <= amplifier_0_2_data_47;
    end else begin
      amplifier_1_0_data_47 <= amplifier_0_0_data_47;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_48 <= amplifier_0_2_data_48;
    end else begin
      amplifier_1_0_data_48 <= amplifier_0_0_data_48;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_49 <= amplifier_0_2_data_49;
    end else begin
      amplifier_1_0_data_49 <= amplifier_0_0_data_49;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_50 <= amplifier_0_2_data_50;
    end else begin
      amplifier_1_0_data_50 <= amplifier_0_0_data_50;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_51 <= amplifier_0_2_data_51;
    end else begin
      amplifier_1_0_data_51 <= amplifier_0_0_data_51;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_52 <= amplifier_0_2_data_52;
    end else begin
      amplifier_1_0_data_52 <= amplifier_0_0_data_52;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_53 <= amplifier_0_2_data_53;
    end else begin
      amplifier_1_0_data_53 <= amplifier_0_0_data_53;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_54 <= amplifier_0_2_data_54;
    end else begin
      amplifier_1_0_data_54 <= amplifier_0_0_data_54;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_55 <= amplifier_0_2_data_55;
    end else begin
      amplifier_1_0_data_55 <= amplifier_0_0_data_55;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_56 <= amplifier_0_2_data_56;
    end else begin
      amplifier_1_0_data_56 <= amplifier_0_0_data_56;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_57 <= amplifier_0_2_data_57;
    end else begin
      amplifier_1_0_data_57 <= amplifier_0_0_data_57;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_58 <= amplifier_0_2_data_58;
    end else begin
      amplifier_1_0_data_58 <= amplifier_0_0_data_58;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_59 <= amplifier_0_2_data_59;
    end else begin
      amplifier_1_0_data_59 <= amplifier_0_0_data_59;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_60 <= amplifier_0_2_data_60;
    end else begin
      amplifier_1_0_data_60 <= amplifier_0_0_data_60;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_61 <= amplifier_0_2_data_61;
    end else begin
      amplifier_1_0_data_61 <= amplifier_0_0_data_61;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_62 <= amplifier_0_2_data_62;
    end else begin
      amplifier_1_0_data_62 <= amplifier_0_0_data_62;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_63 <= amplifier_0_2_data_63;
    end else begin
      amplifier_1_0_data_63 <= amplifier_0_0_data_63;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_64 <= amplifier_0_2_data_64;
    end else begin
      amplifier_1_0_data_64 <= amplifier_0_0_data_64;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_65 <= amplifier_0_2_data_65;
    end else begin
      amplifier_1_0_data_65 <= amplifier_0_0_data_65;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_66 <= amplifier_0_2_data_66;
    end else begin
      amplifier_1_0_data_66 <= amplifier_0_0_data_66;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_67 <= amplifier_0_2_data_67;
    end else begin
      amplifier_1_0_data_67 <= amplifier_0_0_data_67;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_68 <= amplifier_0_2_data_68;
    end else begin
      amplifier_1_0_data_68 <= amplifier_0_0_data_68;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_69 <= amplifier_0_2_data_69;
    end else begin
      amplifier_1_0_data_69 <= amplifier_0_0_data_69;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_70 <= amplifier_0_2_data_70;
    end else begin
      amplifier_1_0_data_70 <= amplifier_0_0_data_70;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_71 <= amplifier_0_2_data_71;
    end else begin
      amplifier_1_0_data_71 <= amplifier_0_0_data_71;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_72 <= amplifier_0_2_data_72;
    end else begin
      amplifier_1_0_data_72 <= amplifier_0_0_data_72;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_73 <= amplifier_0_2_data_73;
    end else begin
      amplifier_1_0_data_73 <= amplifier_0_0_data_73;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_74 <= amplifier_0_2_data_74;
    end else begin
      amplifier_1_0_data_74 <= amplifier_0_0_data_74;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_75 <= amplifier_0_2_data_75;
    end else begin
      amplifier_1_0_data_75 <= amplifier_0_0_data_75;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_76 <= amplifier_0_2_data_76;
    end else begin
      amplifier_1_0_data_76 <= amplifier_0_0_data_76;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_77 <= amplifier_0_2_data_77;
    end else begin
      amplifier_1_0_data_77 <= amplifier_0_0_data_77;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_78 <= amplifier_0_2_data_78;
    end else begin
      amplifier_1_0_data_78 <= amplifier_0_0_data_78;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_79 <= amplifier_0_2_data_79;
    end else begin
      amplifier_1_0_data_79 <= amplifier_0_0_data_79;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_80 <= amplifier_0_2_data_80;
    end else begin
      amplifier_1_0_data_80 <= amplifier_0_0_data_80;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_81 <= amplifier_0_2_data_81;
    end else begin
      amplifier_1_0_data_81 <= amplifier_0_0_data_81;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_82 <= amplifier_0_2_data_82;
    end else begin
      amplifier_1_0_data_82 <= amplifier_0_0_data_82;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_83 <= amplifier_0_2_data_83;
    end else begin
      amplifier_1_0_data_83 <= amplifier_0_0_data_83;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_84 <= amplifier_0_2_data_84;
    end else begin
      amplifier_1_0_data_84 <= amplifier_0_0_data_84;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_85 <= amplifier_0_2_data_85;
    end else begin
      amplifier_1_0_data_85 <= amplifier_0_0_data_85;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_86 <= amplifier_0_2_data_86;
    end else begin
      amplifier_1_0_data_86 <= amplifier_0_0_data_86;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_87 <= amplifier_0_2_data_87;
    end else begin
      amplifier_1_0_data_87 <= amplifier_0_0_data_87;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_88 <= amplifier_0_2_data_88;
    end else begin
      amplifier_1_0_data_88 <= amplifier_0_0_data_88;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_89 <= amplifier_0_2_data_89;
    end else begin
      amplifier_1_0_data_89 <= amplifier_0_0_data_89;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_90 <= amplifier_0_2_data_90;
    end else begin
      amplifier_1_0_data_90 <= amplifier_0_0_data_90;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_91 <= amplifier_0_2_data_91;
    end else begin
      amplifier_1_0_data_91 <= amplifier_0_0_data_91;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_92 <= amplifier_0_2_data_92;
    end else begin
      amplifier_1_0_data_92 <= amplifier_0_0_data_92;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_93 <= amplifier_0_2_data_93;
    end else begin
      amplifier_1_0_data_93 <= amplifier_0_0_data_93;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_94 <= amplifier_0_2_data_94;
    end else begin
      amplifier_1_0_data_94 <= amplifier_0_0_data_94;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_95 <= amplifier_0_2_data_95;
    end else begin
      amplifier_1_0_data_95 <= amplifier_0_0_data_95;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_96 <= amplifier_0_2_data_96;
    end else begin
      amplifier_1_0_data_96 <= amplifier_0_0_data_96;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_97 <= amplifier_0_2_data_97;
    end else begin
      amplifier_1_0_data_97 <= amplifier_0_0_data_97;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_98 <= amplifier_0_2_data_98;
    end else begin
      amplifier_1_0_data_98 <= amplifier_0_0_data_98;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_99 <= amplifier_0_2_data_99;
    end else begin
      amplifier_1_0_data_99 <= amplifier_0_0_data_99;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_100 <= amplifier_0_2_data_100;
    end else begin
      amplifier_1_0_data_100 <= amplifier_0_0_data_100;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_101 <= amplifier_0_2_data_101;
    end else begin
      amplifier_1_0_data_101 <= amplifier_0_0_data_101;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_102 <= amplifier_0_2_data_102;
    end else begin
      amplifier_1_0_data_102 <= amplifier_0_0_data_102;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_103 <= amplifier_0_2_data_103;
    end else begin
      amplifier_1_0_data_103 <= amplifier_0_0_data_103;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_104 <= amplifier_0_2_data_104;
    end else begin
      amplifier_1_0_data_104 <= amplifier_0_0_data_104;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_105 <= amplifier_0_2_data_105;
    end else begin
      amplifier_1_0_data_105 <= amplifier_0_0_data_105;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_106 <= amplifier_0_2_data_106;
    end else begin
      amplifier_1_0_data_106 <= amplifier_0_0_data_106;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_107 <= amplifier_0_2_data_107;
    end else begin
      amplifier_1_0_data_107 <= amplifier_0_0_data_107;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_108 <= amplifier_0_2_data_108;
    end else begin
      amplifier_1_0_data_108 <= amplifier_0_0_data_108;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_109 <= amplifier_0_2_data_109;
    end else begin
      amplifier_1_0_data_109 <= amplifier_0_0_data_109;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_110 <= amplifier_0_2_data_110;
    end else begin
      amplifier_1_0_data_110 <= amplifier_0_0_data_110;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_111 <= amplifier_0_2_data_111;
    end else begin
      amplifier_1_0_data_111 <= amplifier_0_0_data_111;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_112 <= amplifier_0_2_data_112;
    end else begin
      amplifier_1_0_data_112 <= amplifier_0_0_data_112;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_113 <= amplifier_0_2_data_113;
    end else begin
      amplifier_1_0_data_113 <= amplifier_0_0_data_113;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_114 <= amplifier_0_2_data_114;
    end else begin
      amplifier_1_0_data_114 <= amplifier_0_0_data_114;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_115 <= amplifier_0_2_data_115;
    end else begin
      amplifier_1_0_data_115 <= amplifier_0_0_data_115;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_116 <= amplifier_0_2_data_116;
    end else begin
      amplifier_1_0_data_116 <= amplifier_0_0_data_116;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_117 <= amplifier_0_2_data_117;
    end else begin
      amplifier_1_0_data_117 <= amplifier_0_0_data_117;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_118 <= amplifier_0_2_data_118;
    end else begin
      amplifier_1_0_data_118 <= amplifier_0_0_data_118;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_119 <= amplifier_0_2_data_119;
    end else begin
      amplifier_1_0_data_119 <= amplifier_0_0_data_119;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_120 <= amplifier_0_2_data_120;
    end else begin
      amplifier_1_0_data_120 <= amplifier_0_0_data_120;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_121 <= amplifier_0_2_data_121;
    end else begin
      amplifier_1_0_data_121 <= amplifier_0_0_data_121;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_122 <= amplifier_0_2_data_122;
    end else begin
      amplifier_1_0_data_122 <= amplifier_0_0_data_122;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_123 <= amplifier_0_2_data_123;
    end else begin
      amplifier_1_0_data_123 <= amplifier_0_0_data_123;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_124 <= amplifier_0_2_data_124;
    end else begin
      amplifier_1_0_data_124 <= amplifier_0_0_data_124;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_125 <= amplifier_0_2_data_125;
    end else begin
      amplifier_1_0_data_125 <= amplifier_0_0_data_125;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_126 <= amplifier_0_2_data_126;
    end else begin
      amplifier_1_0_data_126 <= amplifier_0_0_data_126;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_127 <= amplifier_0_2_data_127;
    end else begin
      amplifier_1_0_data_127 <= amplifier_0_0_data_127;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_128 <= amplifier_0_2_data_128;
    end else begin
      amplifier_1_0_data_128 <= amplifier_0_0_data_128;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_129 <= amplifier_0_2_data_129;
    end else begin
      amplifier_1_0_data_129 <= amplifier_0_0_data_129;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_130 <= amplifier_0_2_data_130;
    end else begin
      amplifier_1_0_data_130 <= amplifier_0_0_data_130;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_131 <= amplifier_0_2_data_131;
    end else begin
      amplifier_1_0_data_131 <= amplifier_0_0_data_131;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_132 <= amplifier_0_2_data_132;
    end else begin
      amplifier_1_0_data_132 <= amplifier_0_0_data_132;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_133 <= amplifier_0_2_data_133;
    end else begin
      amplifier_1_0_data_133 <= amplifier_0_0_data_133;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_134 <= amplifier_0_2_data_134;
    end else begin
      amplifier_1_0_data_134 <= amplifier_0_0_data_134;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_135 <= amplifier_0_2_data_135;
    end else begin
      amplifier_1_0_data_135 <= amplifier_0_0_data_135;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_136 <= amplifier_0_2_data_136;
    end else begin
      amplifier_1_0_data_136 <= amplifier_0_0_data_136;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_137 <= amplifier_0_2_data_137;
    end else begin
      amplifier_1_0_data_137 <= amplifier_0_0_data_137;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_138 <= amplifier_0_2_data_138;
    end else begin
      amplifier_1_0_data_138 <= amplifier_0_0_data_138;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_139 <= amplifier_0_2_data_139;
    end else begin
      amplifier_1_0_data_139 <= amplifier_0_0_data_139;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_140 <= amplifier_0_2_data_140;
    end else begin
      amplifier_1_0_data_140 <= amplifier_0_0_data_140;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_141 <= amplifier_0_2_data_141;
    end else begin
      amplifier_1_0_data_141 <= amplifier_0_0_data_141;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_142 <= amplifier_0_2_data_142;
    end else begin
      amplifier_1_0_data_142 <= amplifier_0_0_data_142;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_143 <= amplifier_0_2_data_143;
    end else begin
      amplifier_1_0_data_143 <= amplifier_0_0_data_143;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_144 <= amplifier_0_2_data_144;
    end else begin
      amplifier_1_0_data_144 <= amplifier_0_0_data_144;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_145 <= amplifier_0_2_data_145;
    end else begin
      amplifier_1_0_data_145 <= amplifier_0_0_data_145;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_146 <= amplifier_0_2_data_146;
    end else begin
      amplifier_1_0_data_146 <= amplifier_0_0_data_146;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_147 <= amplifier_0_2_data_147;
    end else begin
      amplifier_1_0_data_147 <= amplifier_0_0_data_147;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_148 <= amplifier_0_2_data_148;
    end else begin
      amplifier_1_0_data_148 <= amplifier_0_0_data_148;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_149 <= amplifier_0_2_data_149;
    end else begin
      amplifier_1_0_data_149 <= amplifier_0_0_data_149;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_150 <= amplifier_0_2_data_150;
    end else begin
      amplifier_1_0_data_150 <= amplifier_0_0_data_150;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_151 <= amplifier_0_2_data_151;
    end else begin
      amplifier_1_0_data_151 <= amplifier_0_0_data_151;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_152 <= amplifier_0_2_data_152;
    end else begin
      amplifier_1_0_data_152 <= amplifier_0_0_data_152;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_153 <= amplifier_0_2_data_153;
    end else begin
      amplifier_1_0_data_153 <= amplifier_0_0_data_153;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_154 <= amplifier_0_2_data_154;
    end else begin
      amplifier_1_0_data_154 <= amplifier_0_0_data_154;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_155 <= amplifier_0_2_data_155;
    end else begin
      amplifier_1_0_data_155 <= amplifier_0_0_data_155;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_156 <= amplifier_0_2_data_156;
    end else begin
      amplifier_1_0_data_156 <= amplifier_0_0_data_156;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_157 <= amplifier_0_2_data_157;
    end else begin
      amplifier_1_0_data_157 <= amplifier_0_0_data_157;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_158 <= amplifier_0_2_data_158;
    end else begin
      amplifier_1_0_data_158 <= amplifier_0_0_data_158;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_159 <= amplifier_0_2_data_159;
    end else begin
      amplifier_1_0_data_159 <= amplifier_0_0_data_159;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_160 <= amplifier_0_2_data_160;
    end else begin
      amplifier_1_0_data_160 <= amplifier_0_0_data_160;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_161 <= amplifier_0_2_data_161;
    end else begin
      amplifier_1_0_data_161 <= amplifier_0_0_data_161;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_162 <= amplifier_0_2_data_162;
    end else begin
      amplifier_1_0_data_162 <= amplifier_0_0_data_162;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_163 <= amplifier_0_2_data_163;
    end else begin
      amplifier_1_0_data_163 <= amplifier_0_0_data_163;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_164 <= amplifier_0_2_data_164;
    end else begin
      amplifier_1_0_data_164 <= amplifier_0_0_data_164;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_165 <= amplifier_0_2_data_165;
    end else begin
      amplifier_1_0_data_165 <= amplifier_0_0_data_165;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_166 <= amplifier_0_2_data_166;
    end else begin
      amplifier_1_0_data_166 <= amplifier_0_0_data_166;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_167 <= amplifier_0_2_data_167;
    end else begin
      amplifier_1_0_data_167 <= amplifier_0_0_data_167;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_168 <= amplifier_0_2_data_168;
    end else begin
      amplifier_1_0_data_168 <= amplifier_0_0_data_168;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_169 <= amplifier_0_2_data_169;
    end else begin
      amplifier_1_0_data_169 <= amplifier_0_0_data_169;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_170 <= amplifier_0_2_data_170;
    end else begin
      amplifier_1_0_data_170 <= amplifier_0_0_data_170;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_171 <= amplifier_0_2_data_171;
    end else begin
      amplifier_1_0_data_171 <= amplifier_0_0_data_171;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_172 <= amplifier_0_2_data_172;
    end else begin
      amplifier_1_0_data_172 <= amplifier_0_0_data_172;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_173 <= amplifier_0_2_data_173;
    end else begin
      amplifier_1_0_data_173 <= amplifier_0_0_data_173;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_174 <= amplifier_0_2_data_174;
    end else begin
      amplifier_1_0_data_174 <= amplifier_0_0_data_174;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_175 <= amplifier_0_2_data_175;
    end else begin
      amplifier_1_0_data_175 <= amplifier_0_0_data_175;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_176 <= amplifier_0_2_data_176;
    end else begin
      amplifier_1_0_data_176 <= amplifier_0_0_data_176;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_177 <= amplifier_0_2_data_177;
    end else begin
      amplifier_1_0_data_177 <= amplifier_0_0_data_177;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_178 <= amplifier_0_2_data_178;
    end else begin
      amplifier_1_0_data_178 <= amplifier_0_0_data_178;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_179 <= amplifier_0_2_data_179;
    end else begin
      amplifier_1_0_data_179 <= amplifier_0_0_data_179;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_180 <= amplifier_0_2_data_180;
    end else begin
      amplifier_1_0_data_180 <= amplifier_0_0_data_180;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_181 <= amplifier_0_2_data_181;
    end else begin
      amplifier_1_0_data_181 <= amplifier_0_0_data_181;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_182 <= amplifier_0_2_data_182;
    end else begin
      amplifier_1_0_data_182 <= amplifier_0_0_data_182;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_183 <= amplifier_0_2_data_183;
    end else begin
      amplifier_1_0_data_183 <= amplifier_0_0_data_183;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_184 <= amplifier_0_2_data_184;
    end else begin
      amplifier_1_0_data_184 <= amplifier_0_0_data_184;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_185 <= amplifier_0_2_data_185;
    end else begin
      amplifier_1_0_data_185 <= amplifier_0_0_data_185;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_186 <= amplifier_0_2_data_186;
    end else begin
      amplifier_1_0_data_186 <= amplifier_0_0_data_186;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_187 <= amplifier_0_2_data_187;
    end else begin
      amplifier_1_0_data_187 <= amplifier_0_0_data_187;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_188 <= amplifier_0_2_data_188;
    end else begin
      amplifier_1_0_data_188 <= amplifier_0_0_data_188;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_189 <= amplifier_0_2_data_189;
    end else begin
      amplifier_1_0_data_189 <= amplifier_0_0_data_189;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_190 <= amplifier_0_2_data_190;
    end else begin
      amplifier_1_0_data_190 <= amplifier_0_0_data_190;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_191 <= amplifier_0_2_data_191;
    end else begin
      amplifier_1_0_data_191 <= amplifier_0_0_data_191;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_192 <= amplifier_0_2_data_192;
    end else begin
      amplifier_1_0_data_192 <= amplifier_0_0_data_192;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_193 <= amplifier_0_2_data_193;
    end else begin
      amplifier_1_0_data_193 <= amplifier_0_0_data_193;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_194 <= amplifier_0_2_data_194;
    end else begin
      amplifier_1_0_data_194 <= amplifier_0_0_data_194;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_195 <= amplifier_0_2_data_195;
    end else begin
      amplifier_1_0_data_195 <= amplifier_0_0_data_195;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_196 <= amplifier_0_2_data_196;
    end else begin
      amplifier_1_0_data_196 <= amplifier_0_0_data_196;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_197 <= amplifier_0_2_data_197;
    end else begin
      amplifier_1_0_data_197 <= amplifier_0_0_data_197;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_198 <= amplifier_0_2_data_198;
    end else begin
      amplifier_1_0_data_198 <= amplifier_0_0_data_198;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_199 <= amplifier_0_2_data_199;
    end else begin
      amplifier_1_0_data_199 <= amplifier_0_0_data_199;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_200 <= amplifier_0_2_data_200;
    end else begin
      amplifier_1_0_data_200 <= amplifier_0_0_data_200;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_201 <= amplifier_0_2_data_201;
    end else begin
      amplifier_1_0_data_201 <= amplifier_0_0_data_201;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_202 <= amplifier_0_2_data_202;
    end else begin
      amplifier_1_0_data_202 <= amplifier_0_0_data_202;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_203 <= amplifier_0_2_data_203;
    end else begin
      amplifier_1_0_data_203 <= amplifier_0_0_data_203;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_204 <= amplifier_0_2_data_204;
    end else begin
      amplifier_1_0_data_204 <= amplifier_0_0_data_204;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_205 <= amplifier_0_2_data_205;
    end else begin
      amplifier_1_0_data_205 <= amplifier_0_0_data_205;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_206 <= amplifier_0_2_data_206;
    end else begin
      amplifier_1_0_data_206 <= amplifier_0_0_data_206;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_207 <= amplifier_0_2_data_207;
    end else begin
      amplifier_1_0_data_207 <= amplifier_0_0_data_207;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_208 <= amplifier_0_2_data_208;
    end else begin
      amplifier_1_0_data_208 <= amplifier_0_0_data_208;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_209 <= amplifier_0_2_data_209;
    end else begin
      amplifier_1_0_data_209 <= amplifier_0_0_data_209;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_210 <= amplifier_0_2_data_210;
    end else begin
      amplifier_1_0_data_210 <= amplifier_0_0_data_210;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_211 <= amplifier_0_2_data_211;
    end else begin
      amplifier_1_0_data_211 <= amplifier_0_0_data_211;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_212 <= amplifier_0_2_data_212;
    end else begin
      amplifier_1_0_data_212 <= amplifier_0_0_data_212;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_213 <= amplifier_0_2_data_213;
    end else begin
      amplifier_1_0_data_213 <= amplifier_0_0_data_213;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_214 <= amplifier_0_2_data_214;
    end else begin
      amplifier_1_0_data_214 <= amplifier_0_0_data_214;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_215 <= amplifier_0_2_data_215;
    end else begin
      amplifier_1_0_data_215 <= amplifier_0_0_data_215;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_216 <= amplifier_0_2_data_216;
    end else begin
      amplifier_1_0_data_216 <= amplifier_0_0_data_216;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_217 <= amplifier_0_2_data_217;
    end else begin
      amplifier_1_0_data_217 <= amplifier_0_0_data_217;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_218 <= amplifier_0_2_data_218;
    end else begin
      amplifier_1_0_data_218 <= amplifier_0_0_data_218;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_219 <= amplifier_0_2_data_219;
    end else begin
      amplifier_1_0_data_219 <= amplifier_0_0_data_219;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_220 <= amplifier_0_2_data_220;
    end else begin
      amplifier_1_0_data_220 <= amplifier_0_0_data_220;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_221 <= amplifier_0_2_data_221;
    end else begin
      amplifier_1_0_data_221 <= amplifier_0_0_data_221;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_222 <= amplifier_0_2_data_222;
    end else begin
      amplifier_1_0_data_222 <= amplifier_0_0_data_222;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_223 <= amplifier_0_2_data_223;
    end else begin
      amplifier_1_0_data_223 <= amplifier_0_0_data_223;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_224 <= amplifier_0_2_data_224;
    end else begin
      amplifier_1_0_data_224 <= amplifier_0_0_data_224;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_225 <= amplifier_0_2_data_225;
    end else begin
      amplifier_1_0_data_225 <= amplifier_0_0_data_225;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_226 <= amplifier_0_2_data_226;
    end else begin
      amplifier_1_0_data_226 <= amplifier_0_0_data_226;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_227 <= amplifier_0_2_data_227;
    end else begin
      amplifier_1_0_data_227 <= amplifier_0_0_data_227;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_228 <= amplifier_0_2_data_228;
    end else begin
      amplifier_1_0_data_228 <= amplifier_0_0_data_228;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_229 <= amplifier_0_2_data_229;
    end else begin
      amplifier_1_0_data_229 <= amplifier_0_0_data_229;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_230 <= amplifier_0_2_data_230;
    end else begin
      amplifier_1_0_data_230 <= amplifier_0_0_data_230;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_231 <= amplifier_0_2_data_231;
    end else begin
      amplifier_1_0_data_231 <= amplifier_0_0_data_231;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_232 <= amplifier_0_2_data_232;
    end else begin
      amplifier_1_0_data_232 <= amplifier_0_0_data_232;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_233 <= amplifier_0_2_data_233;
    end else begin
      amplifier_1_0_data_233 <= amplifier_0_0_data_233;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_234 <= amplifier_0_2_data_234;
    end else begin
      amplifier_1_0_data_234 <= amplifier_0_0_data_234;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_235 <= amplifier_0_2_data_235;
    end else begin
      amplifier_1_0_data_235 <= amplifier_0_0_data_235;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_236 <= amplifier_0_2_data_236;
    end else begin
      amplifier_1_0_data_236 <= amplifier_0_0_data_236;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_237 <= amplifier_0_2_data_237;
    end else begin
      amplifier_1_0_data_237 <= amplifier_0_0_data_237;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_238 <= amplifier_0_2_data_238;
    end else begin
      amplifier_1_0_data_238 <= amplifier_0_0_data_238;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_239 <= amplifier_0_2_data_239;
    end else begin
      amplifier_1_0_data_239 <= amplifier_0_0_data_239;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_240 <= amplifier_0_2_data_240;
    end else begin
      amplifier_1_0_data_240 <= amplifier_0_0_data_240;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_241 <= amplifier_0_2_data_241;
    end else begin
      amplifier_1_0_data_241 <= amplifier_0_0_data_241;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_242 <= amplifier_0_2_data_242;
    end else begin
      amplifier_1_0_data_242 <= amplifier_0_0_data_242;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_243 <= amplifier_0_2_data_243;
    end else begin
      amplifier_1_0_data_243 <= amplifier_0_0_data_243;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_244 <= amplifier_0_2_data_244;
    end else begin
      amplifier_1_0_data_244 <= amplifier_0_0_data_244;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_245 <= amplifier_0_2_data_245;
    end else begin
      amplifier_1_0_data_245 <= amplifier_0_0_data_245;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_246 <= amplifier_0_2_data_246;
    end else begin
      amplifier_1_0_data_246 <= amplifier_0_0_data_246;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_247 <= amplifier_0_2_data_247;
    end else begin
      amplifier_1_0_data_247 <= amplifier_0_0_data_247;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_248 <= amplifier_0_2_data_248;
    end else begin
      amplifier_1_0_data_248 <= amplifier_0_0_data_248;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_249 <= amplifier_0_2_data_249;
    end else begin
      amplifier_1_0_data_249 <= amplifier_0_0_data_249;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_250 <= amplifier_0_2_data_250;
    end else begin
      amplifier_1_0_data_250 <= amplifier_0_0_data_250;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_251 <= amplifier_0_2_data_251;
    end else begin
      amplifier_1_0_data_251 <= amplifier_0_0_data_251;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_252 <= amplifier_0_2_data_252;
    end else begin
      amplifier_1_0_data_252 <= amplifier_0_0_data_252;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_253 <= amplifier_0_2_data_253;
    end else begin
      amplifier_1_0_data_253 <= amplifier_0_0_data_253;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_254 <= amplifier_0_2_data_254;
    end else begin
      amplifier_1_0_data_254 <= amplifier_0_0_data_254;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_data_255 <= amplifier_0_2_data_255;
    end else begin
      amplifier_1_0_data_255 <= amplifier_0_0_data_255;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_header_0 <= amplifier_0_2_header_0;
    end else begin
      amplifier_1_0_header_0 <= amplifier_0_0_header_0;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_header_1 <= amplifier_0_2_header_1;
    end else begin
      amplifier_1_0_header_1 <= amplifier_0_0_header_1;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_header_2 <= amplifier_0_2_header_2;
    end else begin
      amplifier_1_0_header_2 <= amplifier_0_0_header_2;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_header_3 <= amplifier_0_2_header_3;
    end else begin
      amplifier_1_0_header_3 <= amplifier_0_0_header_3;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_header_4 <= amplifier_0_2_header_4;
    end else begin
      amplifier_1_0_header_4 <= amplifier_0_0_header_4;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_header_5 <= amplifier_0_2_header_5;
    end else begin
      amplifier_1_0_header_5 <= amplifier_0_0_header_5;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_header_6 <= amplifier_0_2_header_6;
    end else begin
      amplifier_1_0_header_6 <= amplifier_0_0_header_6;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_header_7 <= amplifier_0_2_header_7;
    end else begin
      amplifier_1_0_header_7 <= amplifier_0_0_header_7;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_header_8 <= amplifier_0_2_header_8;
    end else begin
      amplifier_1_0_header_8 <= amplifier_0_0_header_8;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_header_9 <= amplifier_0_2_header_9;
    end else begin
      amplifier_1_0_header_9 <= amplifier_0_0_header_9;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_header_10 <= amplifier_0_2_header_10;
    end else begin
      amplifier_1_0_header_10 <= amplifier_0_0_header_10;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_header_11 <= amplifier_0_2_header_11;
    end else begin
      amplifier_1_0_header_11 <= amplifier_0_0_header_11;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_header_12 <= amplifier_0_2_header_12;
    end else begin
      amplifier_1_0_header_12 <= amplifier_0_0_header_12;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_header_13 <= amplifier_0_2_header_13;
    end else begin
      amplifier_1_0_header_13 <= amplifier_0_0_header_13;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_header_14 <= amplifier_0_2_header_14;
    end else begin
      amplifier_1_0_header_14 <= amplifier_0_0_header_14;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_header_15 <= amplifier_0_2_header_15;
    end else begin
      amplifier_1_0_header_15 <= amplifier_0_0_header_15;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_parse_current_state <= amplifier_0_2_parse_current_state;
    end else begin
      amplifier_1_0_parse_current_state <= amplifier_0_0_parse_current_state;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_parse_current_offset <= amplifier_0_2_parse_current_offset;
    end else begin
      amplifier_1_0_parse_current_offset <= amplifier_0_0_parse_current_offset;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_parse_transition_field <= amplifier_0_2_parse_transition_field;
    end else begin
      amplifier_1_0_parse_transition_field <= amplifier_0_0_parse_transition_field;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_next_processor_id <= amplifier_0_2_next_processor_id;
    end else begin
      amplifier_1_0_next_processor_id <= amplifier_0_0_next_processor_id;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_next_config_id <= amplifier_0_2_next_config_id;
    end else begin
      amplifier_1_0_next_config_id <= amplifier_0_0_next_config_id;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 135:31]
      amplifier_1_0_is_valid_processor <= amplifier_0_2_is_valid_processor;
    end else begin
      amplifier_1_0_is_valid_processor <= amplifier_0_0_is_valid_processor;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_0 <= amplifier_0_3_data_0;
    end else begin
      amplifier_1_1_data_0 <= amplifier_0_1_data_0;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_1 <= amplifier_0_3_data_1;
    end else begin
      amplifier_1_1_data_1 <= amplifier_0_1_data_1;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_2 <= amplifier_0_3_data_2;
    end else begin
      amplifier_1_1_data_2 <= amplifier_0_1_data_2;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_3 <= amplifier_0_3_data_3;
    end else begin
      amplifier_1_1_data_3 <= amplifier_0_1_data_3;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_4 <= amplifier_0_3_data_4;
    end else begin
      amplifier_1_1_data_4 <= amplifier_0_1_data_4;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_5 <= amplifier_0_3_data_5;
    end else begin
      amplifier_1_1_data_5 <= amplifier_0_1_data_5;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_6 <= amplifier_0_3_data_6;
    end else begin
      amplifier_1_1_data_6 <= amplifier_0_1_data_6;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_7 <= amplifier_0_3_data_7;
    end else begin
      amplifier_1_1_data_7 <= amplifier_0_1_data_7;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_8 <= amplifier_0_3_data_8;
    end else begin
      amplifier_1_1_data_8 <= amplifier_0_1_data_8;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_9 <= amplifier_0_3_data_9;
    end else begin
      amplifier_1_1_data_9 <= amplifier_0_1_data_9;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_10 <= amplifier_0_3_data_10;
    end else begin
      amplifier_1_1_data_10 <= amplifier_0_1_data_10;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_11 <= amplifier_0_3_data_11;
    end else begin
      amplifier_1_1_data_11 <= amplifier_0_1_data_11;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_12 <= amplifier_0_3_data_12;
    end else begin
      amplifier_1_1_data_12 <= amplifier_0_1_data_12;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_13 <= amplifier_0_3_data_13;
    end else begin
      amplifier_1_1_data_13 <= amplifier_0_1_data_13;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_14 <= amplifier_0_3_data_14;
    end else begin
      amplifier_1_1_data_14 <= amplifier_0_1_data_14;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_15 <= amplifier_0_3_data_15;
    end else begin
      amplifier_1_1_data_15 <= amplifier_0_1_data_15;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_16 <= amplifier_0_3_data_16;
    end else begin
      amplifier_1_1_data_16 <= amplifier_0_1_data_16;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_17 <= amplifier_0_3_data_17;
    end else begin
      amplifier_1_1_data_17 <= amplifier_0_1_data_17;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_18 <= amplifier_0_3_data_18;
    end else begin
      amplifier_1_1_data_18 <= amplifier_0_1_data_18;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_19 <= amplifier_0_3_data_19;
    end else begin
      amplifier_1_1_data_19 <= amplifier_0_1_data_19;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_20 <= amplifier_0_3_data_20;
    end else begin
      amplifier_1_1_data_20 <= amplifier_0_1_data_20;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_21 <= amplifier_0_3_data_21;
    end else begin
      amplifier_1_1_data_21 <= amplifier_0_1_data_21;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_22 <= amplifier_0_3_data_22;
    end else begin
      amplifier_1_1_data_22 <= amplifier_0_1_data_22;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_23 <= amplifier_0_3_data_23;
    end else begin
      amplifier_1_1_data_23 <= amplifier_0_1_data_23;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_24 <= amplifier_0_3_data_24;
    end else begin
      amplifier_1_1_data_24 <= amplifier_0_1_data_24;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_25 <= amplifier_0_3_data_25;
    end else begin
      amplifier_1_1_data_25 <= amplifier_0_1_data_25;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_26 <= amplifier_0_3_data_26;
    end else begin
      amplifier_1_1_data_26 <= amplifier_0_1_data_26;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_27 <= amplifier_0_3_data_27;
    end else begin
      amplifier_1_1_data_27 <= amplifier_0_1_data_27;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_28 <= amplifier_0_3_data_28;
    end else begin
      amplifier_1_1_data_28 <= amplifier_0_1_data_28;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_29 <= amplifier_0_3_data_29;
    end else begin
      amplifier_1_1_data_29 <= amplifier_0_1_data_29;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_30 <= amplifier_0_3_data_30;
    end else begin
      amplifier_1_1_data_30 <= amplifier_0_1_data_30;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_31 <= amplifier_0_3_data_31;
    end else begin
      amplifier_1_1_data_31 <= amplifier_0_1_data_31;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_32 <= amplifier_0_3_data_32;
    end else begin
      amplifier_1_1_data_32 <= amplifier_0_1_data_32;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_33 <= amplifier_0_3_data_33;
    end else begin
      amplifier_1_1_data_33 <= amplifier_0_1_data_33;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_34 <= amplifier_0_3_data_34;
    end else begin
      amplifier_1_1_data_34 <= amplifier_0_1_data_34;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_35 <= amplifier_0_3_data_35;
    end else begin
      amplifier_1_1_data_35 <= amplifier_0_1_data_35;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_36 <= amplifier_0_3_data_36;
    end else begin
      amplifier_1_1_data_36 <= amplifier_0_1_data_36;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_37 <= amplifier_0_3_data_37;
    end else begin
      amplifier_1_1_data_37 <= amplifier_0_1_data_37;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_38 <= amplifier_0_3_data_38;
    end else begin
      amplifier_1_1_data_38 <= amplifier_0_1_data_38;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_39 <= amplifier_0_3_data_39;
    end else begin
      amplifier_1_1_data_39 <= amplifier_0_1_data_39;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_40 <= amplifier_0_3_data_40;
    end else begin
      amplifier_1_1_data_40 <= amplifier_0_1_data_40;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_41 <= amplifier_0_3_data_41;
    end else begin
      amplifier_1_1_data_41 <= amplifier_0_1_data_41;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_42 <= amplifier_0_3_data_42;
    end else begin
      amplifier_1_1_data_42 <= amplifier_0_1_data_42;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_43 <= amplifier_0_3_data_43;
    end else begin
      amplifier_1_1_data_43 <= amplifier_0_1_data_43;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_44 <= amplifier_0_3_data_44;
    end else begin
      amplifier_1_1_data_44 <= amplifier_0_1_data_44;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_45 <= amplifier_0_3_data_45;
    end else begin
      amplifier_1_1_data_45 <= amplifier_0_1_data_45;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_46 <= amplifier_0_3_data_46;
    end else begin
      amplifier_1_1_data_46 <= amplifier_0_1_data_46;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_47 <= amplifier_0_3_data_47;
    end else begin
      amplifier_1_1_data_47 <= amplifier_0_1_data_47;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_48 <= amplifier_0_3_data_48;
    end else begin
      amplifier_1_1_data_48 <= amplifier_0_1_data_48;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_49 <= amplifier_0_3_data_49;
    end else begin
      amplifier_1_1_data_49 <= amplifier_0_1_data_49;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_50 <= amplifier_0_3_data_50;
    end else begin
      amplifier_1_1_data_50 <= amplifier_0_1_data_50;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_51 <= amplifier_0_3_data_51;
    end else begin
      amplifier_1_1_data_51 <= amplifier_0_1_data_51;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_52 <= amplifier_0_3_data_52;
    end else begin
      amplifier_1_1_data_52 <= amplifier_0_1_data_52;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_53 <= amplifier_0_3_data_53;
    end else begin
      amplifier_1_1_data_53 <= amplifier_0_1_data_53;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_54 <= amplifier_0_3_data_54;
    end else begin
      amplifier_1_1_data_54 <= amplifier_0_1_data_54;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_55 <= amplifier_0_3_data_55;
    end else begin
      amplifier_1_1_data_55 <= amplifier_0_1_data_55;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_56 <= amplifier_0_3_data_56;
    end else begin
      amplifier_1_1_data_56 <= amplifier_0_1_data_56;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_57 <= amplifier_0_3_data_57;
    end else begin
      amplifier_1_1_data_57 <= amplifier_0_1_data_57;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_58 <= amplifier_0_3_data_58;
    end else begin
      amplifier_1_1_data_58 <= amplifier_0_1_data_58;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_59 <= amplifier_0_3_data_59;
    end else begin
      amplifier_1_1_data_59 <= amplifier_0_1_data_59;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_60 <= amplifier_0_3_data_60;
    end else begin
      amplifier_1_1_data_60 <= amplifier_0_1_data_60;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_61 <= amplifier_0_3_data_61;
    end else begin
      amplifier_1_1_data_61 <= amplifier_0_1_data_61;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_62 <= amplifier_0_3_data_62;
    end else begin
      amplifier_1_1_data_62 <= amplifier_0_1_data_62;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_63 <= amplifier_0_3_data_63;
    end else begin
      amplifier_1_1_data_63 <= amplifier_0_1_data_63;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_64 <= amplifier_0_3_data_64;
    end else begin
      amplifier_1_1_data_64 <= amplifier_0_1_data_64;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_65 <= amplifier_0_3_data_65;
    end else begin
      amplifier_1_1_data_65 <= amplifier_0_1_data_65;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_66 <= amplifier_0_3_data_66;
    end else begin
      amplifier_1_1_data_66 <= amplifier_0_1_data_66;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_67 <= amplifier_0_3_data_67;
    end else begin
      amplifier_1_1_data_67 <= amplifier_0_1_data_67;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_68 <= amplifier_0_3_data_68;
    end else begin
      amplifier_1_1_data_68 <= amplifier_0_1_data_68;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_69 <= amplifier_0_3_data_69;
    end else begin
      amplifier_1_1_data_69 <= amplifier_0_1_data_69;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_70 <= amplifier_0_3_data_70;
    end else begin
      amplifier_1_1_data_70 <= amplifier_0_1_data_70;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_71 <= amplifier_0_3_data_71;
    end else begin
      amplifier_1_1_data_71 <= amplifier_0_1_data_71;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_72 <= amplifier_0_3_data_72;
    end else begin
      amplifier_1_1_data_72 <= amplifier_0_1_data_72;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_73 <= amplifier_0_3_data_73;
    end else begin
      amplifier_1_1_data_73 <= amplifier_0_1_data_73;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_74 <= amplifier_0_3_data_74;
    end else begin
      amplifier_1_1_data_74 <= amplifier_0_1_data_74;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_75 <= amplifier_0_3_data_75;
    end else begin
      amplifier_1_1_data_75 <= amplifier_0_1_data_75;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_76 <= amplifier_0_3_data_76;
    end else begin
      amplifier_1_1_data_76 <= amplifier_0_1_data_76;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_77 <= amplifier_0_3_data_77;
    end else begin
      amplifier_1_1_data_77 <= amplifier_0_1_data_77;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_78 <= amplifier_0_3_data_78;
    end else begin
      amplifier_1_1_data_78 <= amplifier_0_1_data_78;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_79 <= amplifier_0_3_data_79;
    end else begin
      amplifier_1_1_data_79 <= amplifier_0_1_data_79;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_80 <= amplifier_0_3_data_80;
    end else begin
      amplifier_1_1_data_80 <= amplifier_0_1_data_80;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_81 <= amplifier_0_3_data_81;
    end else begin
      amplifier_1_1_data_81 <= amplifier_0_1_data_81;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_82 <= amplifier_0_3_data_82;
    end else begin
      amplifier_1_1_data_82 <= amplifier_0_1_data_82;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_83 <= amplifier_0_3_data_83;
    end else begin
      amplifier_1_1_data_83 <= amplifier_0_1_data_83;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_84 <= amplifier_0_3_data_84;
    end else begin
      amplifier_1_1_data_84 <= amplifier_0_1_data_84;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_85 <= amplifier_0_3_data_85;
    end else begin
      amplifier_1_1_data_85 <= amplifier_0_1_data_85;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_86 <= amplifier_0_3_data_86;
    end else begin
      amplifier_1_1_data_86 <= amplifier_0_1_data_86;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_87 <= amplifier_0_3_data_87;
    end else begin
      amplifier_1_1_data_87 <= amplifier_0_1_data_87;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_88 <= amplifier_0_3_data_88;
    end else begin
      amplifier_1_1_data_88 <= amplifier_0_1_data_88;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_89 <= amplifier_0_3_data_89;
    end else begin
      amplifier_1_1_data_89 <= amplifier_0_1_data_89;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_90 <= amplifier_0_3_data_90;
    end else begin
      amplifier_1_1_data_90 <= amplifier_0_1_data_90;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_91 <= amplifier_0_3_data_91;
    end else begin
      amplifier_1_1_data_91 <= amplifier_0_1_data_91;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_92 <= amplifier_0_3_data_92;
    end else begin
      amplifier_1_1_data_92 <= amplifier_0_1_data_92;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_93 <= amplifier_0_3_data_93;
    end else begin
      amplifier_1_1_data_93 <= amplifier_0_1_data_93;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_94 <= amplifier_0_3_data_94;
    end else begin
      amplifier_1_1_data_94 <= amplifier_0_1_data_94;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_95 <= amplifier_0_3_data_95;
    end else begin
      amplifier_1_1_data_95 <= amplifier_0_1_data_95;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_96 <= amplifier_0_3_data_96;
    end else begin
      amplifier_1_1_data_96 <= amplifier_0_1_data_96;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_97 <= amplifier_0_3_data_97;
    end else begin
      amplifier_1_1_data_97 <= amplifier_0_1_data_97;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_98 <= amplifier_0_3_data_98;
    end else begin
      amplifier_1_1_data_98 <= amplifier_0_1_data_98;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_99 <= amplifier_0_3_data_99;
    end else begin
      amplifier_1_1_data_99 <= amplifier_0_1_data_99;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_100 <= amplifier_0_3_data_100;
    end else begin
      amplifier_1_1_data_100 <= amplifier_0_1_data_100;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_101 <= amplifier_0_3_data_101;
    end else begin
      amplifier_1_1_data_101 <= amplifier_0_1_data_101;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_102 <= amplifier_0_3_data_102;
    end else begin
      amplifier_1_1_data_102 <= amplifier_0_1_data_102;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_103 <= amplifier_0_3_data_103;
    end else begin
      amplifier_1_1_data_103 <= amplifier_0_1_data_103;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_104 <= amplifier_0_3_data_104;
    end else begin
      amplifier_1_1_data_104 <= amplifier_0_1_data_104;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_105 <= amplifier_0_3_data_105;
    end else begin
      amplifier_1_1_data_105 <= amplifier_0_1_data_105;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_106 <= amplifier_0_3_data_106;
    end else begin
      amplifier_1_1_data_106 <= amplifier_0_1_data_106;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_107 <= amplifier_0_3_data_107;
    end else begin
      amplifier_1_1_data_107 <= amplifier_0_1_data_107;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_108 <= amplifier_0_3_data_108;
    end else begin
      amplifier_1_1_data_108 <= amplifier_0_1_data_108;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_109 <= amplifier_0_3_data_109;
    end else begin
      amplifier_1_1_data_109 <= amplifier_0_1_data_109;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_110 <= amplifier_0_3_data_110;
    end else begin
      amplifier_1_1_data_110 <= amplifier_0_1_data_110;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_111 <= amplifier_0_3_data_111;
    end else begin
      amplifier_1_1_data_111 <= amplifier_0_1_data_111;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_112 <= amplifier_0_3_data_112;
    end else begin
      amplifier_1_1_data_112 <= amplifier_0_1_data_112;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_113 <= amplifier_0_3_data_113;
    end else begin
      amplifier_1_1_data_113 <= amplifier_0_1_data_113;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_114 <= amplifier_0_3_data_114;
    end else begin
      amplifier_1_1_data_114 <= amplifier_0_1_data_114;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_115 <= amplifier_0_3_data_115;
    end else begin
      amplifier_1_1_data_115 <= amplifier_0_1_data_115;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_116 <= amplifier_0_3_data_116;
    end else begin
      amplifier_1_1_data_116 <= amplifier_0_1_data_116;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_117 <= amplifier_0_3_data_117;
    end else begin
      amplifier_1_1_data_117 <= amplifier_0_1_data_117;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_118 <= amplifier_0_3_data_118;
    end else begin
      amplifier_1_1_data_118 <= amplifier_0_1_data_118;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_119 <= amplifier_0_3_data_119;
    end else begin
      amplifier_1_1_data_119 <= amplifier_0_1_data_119;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_120 <= amplifier_0_3_data_120;
    end else begin
      amplifier_1_1_data_120 <= amplifier_0_1_data_120;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_121 <= amplifier_0_3_data_121;
    end else begin
      amplifier_1_1_data_121 <= amplifier_0_1_data_121;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_122 <= amplifier_0_3_data_122;
    end else begin
      amplifier_1_1_data_122 <= amplifier_0_1_data_122;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_123 <= amplifier_0_3_data_123;
    end else begin
      amplifier_1_1_data_123 <= amplifier_0_1_data_123;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_124 <= amplifier_0_3_data_124;
    end else begin
      amplifier_1_1_data_124 <= amplifier_0_1_data_124;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_125 <= amplifier_0_3_data_125;
    end else begin
      amplifier_1_1_data_125 <= amplifier_0_1_data_125;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_126 <= amplifier_0_3_data_126;
    end else begin
      amplifier_1_1_data_126 <= amplifier_0_1_data_126;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_127 <= amplifier_0_3_data_127;
    end else begin
      amplifier_1_1_data_127 <= amplifier_0_1_data_127;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_128 <= amplifier_0_3_data_128;
    end else begin
      amplifier_1_1_data_128 <= amplifier_0_1_data_128;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_129 <= amplifier_0_3_data_129;
    end else begin
      amplifier_1_1_data_129 <= amplifier_0_1_data_129;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_130 <= amplifier_0_3_data_130;
    end else begin
      amplifier_1_1_data_130 <= amplifier_0_1_data_130;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_131 <= amplifier_0_3_data_131;
    end else begin
      amplifier_1_1_data_131 <= amplifier_0_1_data_131;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_132 <= amplifier_0_3_data_132;
    end else begin
      amplifier_1_1_data_132 <= amplifier_0_1_data_132;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_133 <= amplifier_0_3_data_133;
    end else begin
      amplifier_1_1_data_133 <= amplifier_0_1_data_133;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_134 <= amplifier_0_3_data_134;
    end else begin
      amplifier_1_1_data_134 <= amplifier_0_1_data_134;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_135 <= amplifier_0_3_data_135;
    end else begin
      amplifier_1_1_data_135 <= amplifier_0_1_data_135;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_136 <= amplifier_0_3_data_136;
    end else begin
      amplifier_1_1_data_136 <= amplifier_0_1_data_136;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_137 <= amplifier_0_3_data_137;
    end else begin
      amplifier_1_1_data_137 <= amplifier_0_1_data_137;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_138 <= amplifier_0_3_data_138;
    end else begin
      amplifier_1_1_data_138 <= amplifier_0_1_data_138;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_139 <= amplifier_0_3_data_139;
    end else begin
      amplifier_1_1_data_139 <= amplifier_0_1_data_139;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_140 <= amplifier_0_3_data_140;
    end else begin
      amplifier_1_1_data_140 <= amplifier_0_1_data_140;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_141 <= amplifier_0_3_data_141;
    end else begin
      amplifier_1_1_data_141 <= amplifier_0_1_data_141;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_142 <= amplifier_0_3_data_142;
    end else begin
      amplifier_1_1_data_142 <= amplifier_0_1_data_142;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_143 <= amplifier_0_3_data_143;
    end else begin
      amplifier_1_1_data_143 <= amplifier_0_1_data_143;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_144 <= amplifier_0_3_data_144;
    end else begin
      amplifier_1_1_data_144 <= amplifier_0_1_data_144;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_145 <= amplifier_0_3_data_145;
    end else begin
      amplifier_1_1_data_145 <= amplifier_0_1_data_145;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_146 <= amplifier_0_3_data_146;
    end else begin
      amplifier_1_1_data_146 <= amplifier_0_1_data_146;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_147 <= amplifier_0_3_data_147;
    end else begin
      amplifier_1_1_data_147 <= amplifier_0_1_data_147;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_148 <= amplifier_0_3_data_148;
    end else begin
      amplifier_1_1_data_148 <= amplifier_0_1_data_148;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_149 <= amplifier_0_3_data_149;
    end else begin
      amplifier_1_1_data_149 <= amplifier_0_1_data_149;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_150 <= amplifier_0_3_data_150;
    end else begin
      amplifier_1_1_data_150 <= amplifier_0_1_data_150;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_151 <= amplifier_0_3_data_151;
    end else begin
      amplifier_1_1_data_151 <= amplifier_0_1_data_151;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_152 <= amplifier_0_3_data_152;
    end else begin
      amplifier_1_1_data_152 <= amplifier_0_1_data_152;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_153 <= amplifier_0_3_data_153;
    end else begin
      amplifier_1_1_data_153 <= amplifier_0_1_data_153;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_154 <= amplifier_0_3_data_154;
    end else begin
      amplifier_1_1_data_154 <= amplifier_0_1_data_154;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_155 <= amplifier_0_3_data_155;
    end else begin
      amplifier_1_1_data_155 <= amplifier_0_1_data_155;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_156 <= amplifier_0_3_data_156;
    end else begin
      amplifier_1_1_data_156 <= amplifier_0_1_data_156;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_157 <= amplifier_0_3_data_157;
    end else begin
      amplifier_1_1_data_157 <= amplifier_0_1_data_157;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_158 <= amplifier_0_3_data_158;
    end else begin
      amplifier_1_1_data_158 <= amplifier_0_1_data_158;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_159 <= amplifier_0_3_data_159;
    end else begin
      amplifier_1_1_data_159 <= amplifier_0_1_data_159;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_160 <= amplifier_0_3_data_160;
    end else begin
      amplifier_1_1_data_160 <= amplifier_0_1_data_160;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_161 <= amplifier_0_3_data_161;
    end else begin
      amplifier_1_1_data_161 <= amplifier_0_1_data_161;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_162 <= amplifier_0_3_data_162;
    end else begin
      amplifier_1_1_data_162 <= amplifier_0_1_data_162;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_163 <= amplifier_0_3_data_163;
    end else begin
      amplifier_1_1_data_163 <= amplifier_0_1_data_163;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_164 <= amplifier_0_3_data_164;
    end else begin
      amplifier_1_1_data_164 <= amplifier_0_1_data_164;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_165 <= amplifier_0_3_data_165;
    end else begin
      amplifier_1_1_data_165 <= amplifier_0_1_data_165;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_166 <= amplifier_0_3_data_166;
    end else begin
      amplifier_1_1_data_166 <= amplifier_0_1_data_166;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_167 <= amplifier_0_3_data_167;
    end else begin
      amplifier_1_1_data_167 <= amplifier_0_1_data_167;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_168 <= amplifier_0_3_data_168;
    end else begin
      amplifier_1_1_data_168 <= amplifier_0_1_data_168;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_169 <= amplifier_0_3_data_169;
    end else begin
      amplifier_1_1_data_169 <= amplifier_0_1_data_169;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_170 <= amplifier_0_3_data_170;
    end else begin
      amplifier_1_1_data_170 <= amplifier_0_1_data_170;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_171 <= amplifier_0_3_data_171;
    end else begin
      amplifier_1_1_data_171 <= amplifier_0_1_data_171;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_172 <= amplifier_0_3_data_172;
    end else begin
      amplifier_1_1_data_172 <= amplifier_0_1_data_172;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_173 <= amplifier_0_3_data_173;
    end else begin
      amplifier_1_1_data_173 <= amplifier_0_1_data_173;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_174 <= amplifier_0_3_data_174;
    end else begin
      amplifier_1_1_data_174 <= amplifier_0_1_data_174;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_175 <= amplifier_0_3_data_175;
    end else begin
      amplifier_1_1_data_175 <= amplifier_0_1_data_175;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_176 <= amplifier_0_3_data_176;
    end else begin
      amplifier_1_1_data_176 <= amplifier_0_1_data_176;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_177 <= amplifier_0_3_data_177;
    end else begin
      amplifier_1_1_data_177 <= amplifier_0_1_data_177;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_178 <= amplifier_0_3_data_178;
    end else begin
      amplifier_1_1_data_178 <= amplifier_0_1_data_178;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_179 <= amplifier_0_3_data_179;
    end else begin
      amplifier_1_1_data_179 <= amplifier_0_1_data_179;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_180 <= amplifier_0_3_data_180;
    end else begin
      amplifier_1_1_data_180 <= amplifier_0_1_data_180;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_181 <= amplifier_0_3_data_181;
    end else begin
      amplifier_1_1_data_181 <= amplifier_0_1_data_181;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_182 <= amplifier_0_3_data_182;
    end else begin
      amplifier_1_1_data_182 <= amplifier_0_1_data_182;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_183 <= amplifier_0_3_data_183;
    end else begin
      amplifier_1_1_data_183 <= amplifier_0_1_data_183;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_184 <= amplifier_0_3_data_184;
    end else begin
      amplifier_1_1_data_184 <= amplifier_0_1_data_184;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_185 <= amplifier_0_3_data_185;
    end else begin
      amplifier_1_1_data_185 <= amplifier_0_1_data_185;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_186 <= amplifier_0_3_data_186;
    end else begin
      amplifier_1_1_data_186 <= amplifier_0_1_data_186;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_187 <= amplifier_0_3_data_187;
    end else begin
      amplifier_1_1_data_187 <= amplifier_0_1_data_187;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_188 <= amplifier_0_3_data_188;
    end else begin
      amplifier_1_1_data_188 <= amplifier_0_1_data_188;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_189 <= amplifier_0_3_data_189;
    end else begin
      amplifier_1_1_data_189 <= amplifier_0_1_data_189;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_190 <= amplifier_0_3_data_190;
    end else begin
      amplifier_1_1_data_190 <= amplifier_0_1_data_190;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_191 <= amplifier_0_3_data_191;
    end else begin
      amplifier_1_1_data_191 <= amplifier_0_1_data_191;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_192 <= amplifier_0_3_data_192;
    end else begin
      amplifier_1_1_data_192 <= amplifier_0_1_data_192;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_193 <= amplifier_0_3_data_193;
    end else begin
      amplifier_1_1_data_193 <= amplifier_0_1_data_193;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_194 <= amplifier_0_3_data_194;
    end else begin
      amplifier_1_1_data_194 <= amplifier_0_1_data_194;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_195 <= amplifier_0_3_data_195;
    end else begin
      amplifier_1_1_data_195 <= amplifier_0_1_data_195;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_196 <= amplifier_0_3_data_196;
    end else begin
      amplifier_1_1_data_196 <= amplifier_0_1_data_196;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_197 <= amplifier_0_3_data_197;
    end else begin
      amplifier_1_1_data_197 <= amplifier_0_1_data_197;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_198 <= amplifier_0_3_data_198;
    end else begin
      amplifier_1_1_data_198 <= amplifier_0_1_data_198;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_199 <= amplifier_0_3_data_199;
    end else begin
      amplifier_1_1_data_199 <= amplifier_0_1_data_199;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_200 <= amplifier_0_3_data_200;
    end else begin
      amplifier_1_1_data_200 <= amplifier_0_1_data_200;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_201 <= amplifier_0_3_data_201;
    end else begin
      amplifier_1_1_data_201 <= amplifier_0_1_data_201;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_202 <= amplifier_0_3_data_202;
    end else begin
      amplifier_1_1_data_202 <= amplifier_0_1_data_202;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_203 <= amplifier_0_3_data_203;
    end else begin
      amplifier_1_1_data_203 <= amplifier_0_1_data_203;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_204 <= amplifier_0_3_data_204;
    end else begin
      amplifier_1_1_data_204 <= amplifier_0_1_data_204;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_205 <= amplifier_0_3_data_205;
    end else begin
      amplifier_1_1_data_205 <= amplifier_0_1_data_205;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_206 <= amplifier_0_3_data_206;
    end else begin
      amplifier_1_1_data_206 <= amplifier_0_1_data_206;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_207 <= amplifier_0_3_data_207;
    end else begin
      amplifier_1_1_data_207 <= amplifier_0_1_data_207;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_208 <= amplifier_0_3_data_208;
    end else begin
      amplifier_1_1_data_208 <= amplifier_0_1_data_208;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_209 <= amplifier_0_3_data_209;
    end else begin
      amplifier_1_1_data_209 <= amplifier_0_1_data_209;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_210 <= amplifier_0_3_data_210;
    end else begin
      amplifier_1_1_data_210 <= amplifier_0_1_data_210;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_211 <= amplifier_0_3_data_211;
    end else begin
      amplifier_1_1_data_211 <= amplifier_0_1_data_211;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_212 <= amplifier_0_3_data_212;
    end else begin
      amplifier_1_1_data_212 <= amplifier_0_1_data_212;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_213 <= amplifier_0_3_data_213;
    end else begin
      amplifier_1_1_data_213 <= amplifier_0_1_data_213;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_214 <= amplifier_0_3_data_214;
    end else begin
      amplifier_1_1_data_214 <= amplifier_0_1_data_214;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_215 <= amplifier_0_3_data_215;
    end else begin
      amplifier_1_1_data_215 <= amplifier_0_1_data_215;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_216 <= amplifier_0_3_data_216;
    end else begin
      amplifier_1_1_data_216 <= amplifier_0_1_data_216;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_217 <= amplifier_0_3_data_217;
    end else begin
      amplifier_1_1_data_217 <= amplifier_0_1_data_217;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_218 <= amplifier_0_3_data_218;
    end else begin
      amplifier_1_1_data_218 <= amplifier_0_1_data_218;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_219 <= amplifier_0_3_data_219;
    end else begin
      amplifier_1_1_data_219 <= amplifier_0_1_data_219;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_220 <= amplifier_0_3_data_220;
    end else begin
      amplifier_1_1_data_220 <= amplifier_0_1_data_220;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_221 <= amplifier_0_3_data_221;
    end else begin
      amplifier_1_1_data_221 <= amplifier_0_1_data_221;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_222 <= amplifier_0_3_data_222;
    end else begin
      amplifier_1_1_data_222 <= amplifier_0_1_data_222;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_223 <= amplifier_0_3_data_223;
    end else begin
      amplifier_1_1_data_223 <= amplifier_0_1_data_223;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_224 <= amplifier_0_3_data_224;
    end else begin
      amplifier_1_1_data_224 <= amplifier_0_1_data_224;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_225 <= amplifier_0_3_data_225;
    end else begin
      amplifier_1_1_data_225 <= amplifier_0_1_data_225;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_226 <= amplifier_0_3_data_226;
    end else begin
      amplifier_1_1_data_226 <= amplifier_0_1_data_226;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_227 <= amplifier_0_3_data_227;
    end else begin
      amplifier_1_1_data_227 <= amplifier_0_1_data_227;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_228 <= amplifier_0_3_data_228;
    end else begin
      amplifier_1_1_data_228 <= amplifier_0_1_data_228;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_229 <= amplifier_0_3_data_229;
    end else begin
      amplifier_1_1_data_229 <= amplifier_0_1_data_229;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_230 <= amplifier_0_3_data_230;
    end else begin
      amplifier_1_1_data_230 <= amplifier_0_1_data_230;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_231 <= amplifier_0_3_data_231;
    end else begin
      amplifier_1_1_data_231 <= amplifier_0_1_data_231;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_232 <= amplifier_0_3_data_232;
    end else begin
      amplifier_1_1_data_232 <= amplifier_0_1_data_232;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_233 <= amplifier_0_3_data_233;
    end else begin
      amplifier_1_1_data_233 <= amplifier_0_1_data_233;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_234 <= amplifier_0_3_data_234;
    end else begin
      amplifier_1_1_data_234 <= amplifier_0_1_data_234;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_235 <= amplifier_0_3_data_235;
    end else begin
      amplifier_1_1_data_235 <= amplifier_0_1_data_235;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_236 <= amplifier_0_3_data_236;
    end else begin
      amplifier_1_1_data_236 <= amplifier_0_1_data_236;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_237 <= amplifier_0_3_data_237;
    end else begin
      amplifier_1_1_data_237 <= amplifier_0_1_data_237;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_238 <= amplifier_0_3_data_238;
    end else begin
      amplifier_1_1_data_238 <= amplifier_0_1_data_238;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_239 <= amplifier_0_3_data_239;
    end else begin
      amplifier_1_1_data_239 <= amplifier_0_1_data_239;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_240 <= amplifier_0_3_data_240;
    end else begin
      amplifier_1_1_data_240 <= amplifier_0_1_data_240;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_241 <= amplifier_0_3_data_241;
    end else begin
      amplifier_1_1_data_241 <= amplifier_0_1_data_241;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_242 <= amplifier_0_3_data_242;
    end else begin
      amplifier_1_1_data_242 <= amplifier_0_1_data_242;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_243 <= amplifier_0_3_data_243;
    end else begin
      amplifier_1_1_data_243 <= amplifier_0_1_data_243;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_244 <= amplifier_0_3_data_244;
    end else begin
      amplifier_1_1_data_244 <= amplifier_0_1_data_244;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_245 <= amplifier_0_3_data_245;
    end else begin
      amplifier_1_1_data_245 <= amplifier_0_1_data_245;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_246 <= amplifier_0_3_data_246;
    end else begin
      amplifier_1_1_data_246 <= amplifier_0_1_data_246;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_247 <= amplifier_0_3_data_247;
    end else begin
      amplifier_1_1_data_247 <= amplifier_0_1_data_247;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_248 <= amplifier_0_3_data_248;
    end else begin
      amplifier_1_1_data_248 <= amplifier_0_1_data_248;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_249 <= amplifier_0_3_data_249;
    end else begin
      amplifier_1_1_data_249 <= amplifier_0_1_data_249;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_250 <= amplifier_0_3_data_250;
    end else begin
      amplifier_1_1_data_250 <= amplifier_0_1_data_250;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_251 <= amplifier_0_3_data_251;
    end else begin
      amplifier_1_1_data_251 <= amplifier_0_1_data_251;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_252 <= amplifier_0_3_data_252;
    end else begin
      amplifier_1_1_data_252 <= amplifier_0_1_data_252;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_253 <= amplifier_0_3_data_253;
    end else begin
      amplifier_1_1_data_253 <= amplifier_0_1_data_253;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_254 <= amplifier_0_3_data_254;
    end else begin
      amplifier_1_1_data_254 <= amplifier_0_1_data_254;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_data_255 <= amplifier_0_3_data_255;
    end else begin
      amplifier_1_1_data_255 <= amplifier_0_1_data_255;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_header_0 <= amplifier_0_3_header_0;
    end else begin
      amplifier_1_1_header_0 <= amplifier_0_1_header_0;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_header_1 <= amplifier_0_3_header_1;
    end else begin
      amplifier_1_1_header_1 <= amplifier_0_1_header_1;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_header_2 <= amplifier_0_3_header_2;
    end else begin
      amplifier_1_1_header_2 <= amplifier_0_1_header_2;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_header_3 <= amplifier_0_3_header_3;
    end else begin
      amplifier_1_1_header_3 <= amplifier_0_1_header_3;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_header_4 <= amplifier_0_3_header_4;
    end else begin
      amplifier_1_1_header_4 <= amplifier_0_1_header_4;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_header_5 <= amplifier_0_3_header_5;
    end else begin
      amplifier_1_1_header_5 <= amplifier_0_1_header_5;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_header_6 <= amplifier_0_3_header_6;
    end else begin
      amplifier_1_1_header_6 <= amplifier_0_1_header_6;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_header_7 <= amplifier_0_3_header_7;
    end else begin
      amplifier_1_1_header_7 <= amplifier_0_1_header_7;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_header_8 <= amplifier_0_3_header_8;
    end else begin
      amplifier_1_1_header_8 <= amplifier_0_1_header_8;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_header_9 <= amplifier_0_3_header_9;
    end else begin
      amplifier_1_1_header_9 <= amplifier_0_1_header_9;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_header_10 <= amplifier_0_3_header_10;
    end else begin
      amplifier_1_1_header_10 <= amplifier_0_1_header_10;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_header_11 <= amplifier_0_3_header_11;
    end else begin
      amplifier_1_1_header_11 <= amplifier_0_1_header_11;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_header_12 <= amplifier_0_3_header_12;
    end else begin
      amplifier_1_1_header_12 <= amplifier_0_1_header_12;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_header_13 <= amplifier_0_3_header_13;
    end else begin
      amplifier_1_1_header_13 <= amplifier_0_1_header_13;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_header_14 <= amplifier_0_3_header_14;
    end else begin
      amplifier_1_1_header_14 <= amplifier_0_1_header_14;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_header_15 <= amplifier_0_3_header_15;
    end else begin
      amplifier_1_1_header_15 <= amplifier_0_1_header_15;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_parse_current_state <= amplifier_0_3_parse_current_state;
    end else begin
      amplifier_1_1_parse_current_state <= amplifier_0_1_parse_current_state;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_parse_current_offset <= amplifier_0_3_parse_current_offset;
    end else begin
      amplifier_1_1_parse_current_offset <= amplifier_0_1_parse_current_offset;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_parse_transition_field <= amplifier_0_3_parse_transition_field;
    end else begin
      amplifier_1_1_parse_transition_field <= amplifier_0_1_parse_transition_field;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_next_processor_id <= amplifier_0_3_next_processor_id;
    end else begin
      amplifier_1_1_next_processor_id <= amplifier_0_1_next_processor_id;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_next_config_id <= amplifier_0_3_next_config_id;
    end else begin
      amplifier_1_1_next_config_id <= amplifier_0_1_next_config_id;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 135:31]
      amplifier_1_1_is_valid_processor <= amplifier_0_3_is_valid_processor;
    end else begin
      amplifier_1_1_is_valid_processor <= amplifier_0_1_is_valid_processor;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_0 <= amplifier_0_0_data_0;
    end else begin
      amplifier_1_2_data_0 <= amplifier_0_2_data_0;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_1 <= amplifier_0_0_data_1;
    end else begin
      amplifier_1_2_data_1 <= amplifier_0_2_data_1;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_2 <= amplifier_0_0_data_2;
    end else begin
      amplifier_1_2_data_2 <= amplifier_0_2_data_2;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_3 <= amplifier_0_0_data_3;
    end else begin
      amplifier_1_2_data_3 <= amplifier_0_2_data_3;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_4 <= amplifier_0_0_data_4;
    end else begin
      amplifier_1_2_data_4 <= amplifier_0_2_data_4;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_5 <= amplifier_0_0_data_5;
    end else begin
      amplifier_1_2_data_5 <= amplifier_0_2_data_5;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_6 <= amplifier_0_0_data_6;
    end else begin
      amplifier_1_2_data_6 <= amplifier_0_2_data_6;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_7 <= amplifier_0_0_data_7;
    end else begin
      amplifier_1_2_data_7 <= amplifier_0_2_data_7;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_8 <= amplifier_0_0_data_8;
    end else begin
      amplifier_1_2_data_8 <= amplifier_0_2_data_8;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_9 <= amplifier_0_0_data_9;
    end else begin
      amplifier_1_2_data_9 <= amplifier_0_2_data_9;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_10 <= amplifier_0_0_data_10;
    end else begin
      amplifier_1_2_data_10 <= amplifier_0_2_data_10;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_11 <= amplifier_0_0_data_11;
    end else begin
      amplifier_1_2_data_11 <= amplifier_0_2_data_11;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_12 <= amplifier_0_0_data_12;
    end else begin
      amplifier_1_2_data_12 <= amplifier_0_2_data_12;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_13 <= amplifier_0_0_data_13;
    end else begin
      amplifier_1_2_data_13 <= amplifier_0_2_data_13;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_14 <= amplifier_0_0_data_14;
    end else begin
      amplifier_1_2_data_14 <= amplifier_0_2_data_14;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_15 <= amplifier_0_0_data_15;
    end else begin
      amplifier_1_2_data_15 <= amplifier_0_2_data_15;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_16 <= amplifier_0_0_data_16;
    end else begin
      amplifier_1_2_data_16 <= amplifier_0_2_data_16;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_17 <= amplifier_0_0_data_17;
    end else begin
      amplifier_1_2_data_17 <= amplifier_0_2_data_17;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_18 <= amplifier_0_0_data_18;
    end else begin
      amplifier_1_2_data_18 <= amplifier_0_2_data_18;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_19 <= amplifier_0_0_data_19;
    end else begin
      amplifier_1_2_data_19 <= amplifier_0_2_data_19;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_20 <= amplifier_0_0_data_20;
    end else begin
      amplifier_1_2_data_20 <= amplifier_0_2_data_20;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_21 <= amplifier_0_0_data_21;
    end else begin
      amplifier_1_2_data_21 <= amplifier_0_2_data_21;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_22 <= amplifier_0_0_data_22;
    end else begin
      amplifier_1_2_data_22 <= amplifier_0_2_data_22;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_23 <= amplifier_0_0_data_23;
    end else begin
      amplifier_1_2_data_23 <= amplifier_0_2_data_23;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_24 <= amplifier_0_0_data_24;
    end else begin
      amplifier_1_2_data_24 <= amplifier_0_2_data_24;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_25 <= amplifier_0_0_data_25;
    end else begin
      amplifier_1_2_data_25 <= amplifier_0_2_data_25;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_26 <= amplifier_0_0_data_26;
    end else begin
      amplifier_1_2_data_26 <= amplifier_0_2_data_26;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_27 <= amplifier_0_0_data_27;
    end else begin
      amplifier_1_2_data_27 <= amplifier_0_2_data_27;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_28 <= amplifier_0_0_data_28;
    end else begin
      amplifier_1_2_data_28 <= amplifier_0_2_data_28;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_29 <= amplifier_0_0_data_29;
    end else begin
      amplifier_1_2_data_29 <= amplifier_0_2_data_29;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_30 <= amplifier_0_0_data_30;
    end else begin
      amplifier_1_2_data_30 <= amplifier_0_2_data_30;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_31 <= amplifier_0_0_data_31;
    end else begin
      amplifier_1_2_data_31 <= amplifier_0_2_data_31;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_32 <= amplifier_0_0_data_32;
    end else begin
      amplifier_1_2_data_32 <= amplifier_0_2_data_32;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_33 <= amplifier_0_0_data_33;
    end else begin
      amplifier_1_2_data_33 <= amplifier_0_2_data_33;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_34 <= amplifier_0_0_data_34;
    end else begin
      amplifier_1_2_data_34 <= amplifier_0_2_data_34;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_35 <= amplifier_0_0_data_35;
    end else begin
      amplifier_1_2_data_35 <= amplifier_0_2_data_35;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_36 <= amplifier_0_0_data_36;
    end else begin
      amplifier_1_2_data_36 <= amplifier_0_2_data_36;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_37 <= amplifier_0_0_data_37;
    end else begin
      amplifier_1_2_data_37 <= amplifier_0_2_data_37;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_38 <= amplifier_0_0_data_38;
    end else begin
      amplifier_1_2_data_38 <= amplifier_0_2_data_38;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_39 <= amplifier_0_0_data_39;
    end else begin
      amplifier_1_2_data_39 <= amplifier_0_2_data_39;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_40 <= amplifier_0_0_data_40;
    end else begin
      amplifier_1_2_data_40 <= amplifier_0_2_data_40;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_41 <= amplifier_0_0_data_41;
    end else begin
      amplifier_1_2_data_41 <= amplifier_0_2_data_41;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_42 <= amplifier_0_0_data_42;
    end else begin
      amplifier_1_2_data_42 <= amplifier_0_2_data_42;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_43 <= amplifier_0_0_data_43;
    end else begin
      amplifier_1_2_data_43 <= amplifier_0_2_data_43;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_44 <= amplifier_0_0_data_44;
    end else begin
      amplifier_1_2_data_44 <= amplifier_0_2_data_44;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_45 <= amplifier_0_0_data_45;
    end else begin
      amplifier_1_2_data_45 <= amplifier_0_2_data_45;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_46 <= amplifier_0_0_data_46;
    end else begin
      amplifier_1_2_data_46 <= amplifier_0_2_data_46;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_47 <= amplifier_0_0_data_47;
    end else begin
      amplifier_1_2_data_47 <= amplifier_0_2_data_47;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_48 <= amplifier_0_0_data_48;
    end else begin
      amplifier_1_2_data_48 <= amplifier_0_2_data_48;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_49 <= amplifier_0_0_data_49;
    end else begin
      amplifier_1_2_data_49 <= amplifier_0_2_data_49;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_50 <= amplifier_0_0_data_50;
    end else begin
      amplifier_1_2_data_50 <= amplifier_0_2_data_50;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_51 <= amplifier_0_0_data_51;
    end else begin
      amplifier_1_2_data_51 <= amplifier_0_2_data_51;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_52 <= amplifier_0_0_data_52;
    end else begin
      amplifier_1_2_data_52 <= amplifier_0_2_data_52;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_53 <= amplifier_0_0_data_53;
    end else begin
      amplifier_1_2_data_53 <= amplifier_0_2_data_53;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_54 <= amplifier_0_0_data_54;
    end else begin
      amplifier_1_2_data_54 <= amplifier_0_2_data_54;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_55 <= amplifier_0_0_data_55;
    end else begin
      amplifier_1_2_data_55 <= amplifier_0_2_data_55;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_56 <= amplifier_0_0_data_56;
    end else begin
      amplifier_1_2_data_56 <= amplifier_0_2_data_56;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_57 <= amplifier_0_0_data_57;
    end else begin
      amplifier_1_2_data_57 <= amplifier_0_2_data_57;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_58 <= amplifier_0_0_data_58;
    end else begin
      amplifier_1_2_data_58 <= amplifier_0_2_data_58;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_59 <= amplifier_0_0_data_59;
    end else begin
      amplifier_1_2_data_59 <= amplifier_0_2_data_59;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_60 <= amplifier_0_0_data_60;
    end else begin
      amplifier_1_2_data_60 <= amplifier_0_2_data_60;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_61 <= amplifier_0_0_data_61;
    end else begin
      amplifier_1_2_data_61 <= amplifier_0_2_data_61;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_62 <= amplifier_0_0_data_62;
    end else begin
      amplifier_1_2_data_62 <= amplifier_0_2_data_62;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_63 <= amplifier_0_0_data_63;
    end else begin
      amplifier_1_2_data_63 <= amplifier_0_2_data_63;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_64 <= amplifier_0_0_data_64;
    end else begin
      amplifier_1_2_data_64 <= amplifier_0_2_data_64;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_65 <= amplifier_0_0_data_65;
    end else begin
      amplifier_1_2_data_65 <= amplifier_0_2_data_65;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_66 <= amplifier_0_0_data_66;
    end else begin
      amplifier_1_2_data_66 <= amplifier_0_2_data_66;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_67 <= amplifier_0_0_data_67;
    end else begin
      amplifier_1_2_data_67 <= amplifier_0_2_data_67;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_68 <= amplifier_0_0_data_68;
    end else begin
      amplifier_1_2_data_68 <= amplifier_0_2_data_68;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_69 <= amplifier_0_0_data_69;
    end else begin
      amplifier_1_2_data_69 <= amplifier_0_2_data_69;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_70 <= amplifier_0_0_data_70;
    end else begin
      amplifier_1_2_data_70 <= amplifier_0_2_data_70;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_71 <= amplifier_0_0_data_71;
    end else begin
      amplifier_1_2_data_71 <= amplifier_0_2_data_71;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_72 <= amplifier_0_0_data_72;
    end else begin
      amplifier_1_2_data_72 <= amplifier_0_2_data_72;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_73 <= amplifier_0_0_data_73;
    end else begin
      amplifier_1_2_data_73 <= amplifier_0_2_data_73;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_74 <= amplifier_0_0_data_74;
    end else begin
      amplifier_1_2_data_74 <= amplifier_0_2_data_74;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_75 <= amplifier_0_0_data_75;
    end else begin
      amplifier_1_2_data_75 <= amplifier_0_2_data_75;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_76 <= amplifier_0_0_data_76;
    end else begin
      amplifier_1_2_data_76 <= amplifier_0_2_data_76;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_77 <= amplifier_0_0_data_77;
    end else begin
      amplifier_1_2_data_77 <= amplifier_0_2_data_77;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_78 <= amplifier_0_0_data_78;
    end else begin
      amplifier_1_2_data_78 <= amplifier_0_2_data_78;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_79 <= amplifier_0_0_data_79;
    end else begin
      amplifier_1_2_data_79 <= amplifier_0_2_data_79;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_80 <= amplifier_0_0_data_80;
    end else begin
      amplifier_1_2_data_80 <= amplifier_0_2_data_80;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_81 <= amplifier_0_0_data_81;
    end else begin
      amplifier_1_2_data_81 <= amplifier_0_2_data_81;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_82 <= amplifier_0_0_data_82;
    end else begin
      amplifier_1_2_data_82 <= amplifier_0_2_data_82;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_83 <= amplifier_0_0_data_83;
    end else begin
      amplifier_1_2_data_83 <= amplifier_0_2_data_83;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_84 <= amplifier_0_0_data_84;
    end else begin
      amplifier_1_2_data_84 <= amplifier_0_2_data_84;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_85 <= amplifier_0_0_data_85;
    end else begin
      amplifier_1_2_data_85 <= amplifier_0_2_data_85;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_86 <= amplifier_0_0_data_86;
    end else begin
      amplifier_1_2_data_86 <= amplifier_0_2_data_86;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_87 <= amplifier_0_0_data_87;
    end else begin
      amplifier_1_2_data_87 <= amplifier_0_2_data_87;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_88 <= amplifier_0_0_data_88;
    end else begin
      amplifier_1_2_data_88 <= amplifier_0_2_data_88;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_89 <= amplifier_0_0_data_89;
    end else begin
      amplifier_1_2_data_89 <= amplifier_0_2_data_89;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_90 <= amplifier_0_0_data_90;
    end else begin
      amplifier_1_2_data_90 <= amplifier_0_2_data_90;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_91 <= amplifier_0_0_data_91;
    end else begin
      amplifier_1_2_data_91 <= amplifier_0_2_data_91;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_92 <= amplifier_0_0_data_92;
    end else begin
      amplifier_1_2_data_92 <= amplifier_0_2_data_92;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_93 <= amplifier_0_0_data_93;
    end else begin
      amplifier_1_2_data_93 <= amplifier_0_2_data_93;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_94 <= amplifier_0_0_data_94;
    end else begin
      amplifier_1_2_data_94 <= amplifier_0_2_data_94;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_95 <= amplifier_0_0_data_95;
    end else begin
      amplifier_1_2_data_95 <= amplifier_0_2_data_95;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_96 <= amplifier_0_0_data_96;
    end else begin
      amplifier_1_2_data_96 <= amplifier_0_2_data_96;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_97 <= amplifier_0_0_data_97;
    end else begin
      amplifier_1_2_data_97 <= amplifier_0_2_data_97;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_98 <= amplifier_0_0_data_98;
    end else begin
      amplifier_1_2_data_98 <= amplifier_0_2_data_98;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_99 <= amplifier_0_0_data_99;
    end else begin
      amplifier_1_2_data_99 <= amplifier_0_2_data_99;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_100 <= amplifier_0_0_data_100;
    end else begin
      amplifier_1_2_data_100 <= amplifier_0_2_data_100;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_101 <= amplifier_0_0_data_101;
    end else begin
      amplifier_1_2_data_101 <= amplifier_0_2_data_101;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_102 <= amplifier_0_0_data_102;
    end else begin
      amplifier_1_2_data_102 <= amplifier_0_2_data_102;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_103 <= amplifier_0_0_data_103;
    end else begin
      amplifier_1_2_data_103 <= amplifier_0_2_data_103;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_104 <= amplifier_0_0_data_104;
    end else begin
      amplifier_1_2_data_104 <= amplifier_0_2_data_104;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_105 <= amplifier_0_0_data_105;
    end else begin
      amplifier_1_2_data_105 <= amplifier_0_2_data_105;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_106 <= amplifier_0_0_data_106;
    end else begin
      amplifier_1_2_data_106 <= amplifier_0_2_data_106;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_107 <= amplifier_0_0_data_107;
    end else begin
      amplifier_1_2_data_107 <= amplifier_0_2_data_107;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_108 <= amplifier_0_0_data_108;
    end else begin
      amplifier_1_2_data_108 <= amplifier_0_2_data_108;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_109 <= amplifier_0_0_data_109;
    end else begin
      amplifier_1_2_data_109 <= amplifier_0_2_data_109;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_110 <= amplifier_0_0_data_110;
    end else begin
      amplifier_1_2_data_110 <= amplifier_0_2_data_110;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_111 <= amplifier_0_0_data_111;
    end else begin
      amplifier_1_2_data_111 <= amplifier_0_2_data_111;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_112 <= amplifier_0_0_data_112;
    end else begin
      amplifier_1_2_data_112 <= amplifier_0_2_data_112;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_113 <= amplifier_0_0_data_113;
    end else begin
      amplifier_1_2_data_113 <= amplifier_0_2_data_113;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_114 <= amplifier_0_0_data_114;
    end else begin
      amplifier_1_2_data_114 <= amplifier_0_2_data_114;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_115 <= amplifier_0_0_data_115;
    end else begin
      amplifier_1_2_data_115 <= amplifier_0_2_data_115;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_116 <= amplifier_0_0_data_116;
    end else begin
      amplifier_1_2_data_116 <= amplifier_0_2_data_116;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_117 <= amplifier_0_0_data_117;
    end else begin
      amplifier_1_2_data_117 <= amplifier_0_2_data_117;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_118 <= amplifier_0_0_data_118;
    end else begin
      amplifier_1_2_data_118 <= amplifier_0_2_data_118;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_119 <= amplifier_0_0_data_119;
    end else begin
      amplifier_1_2_data_119 <= amplifier_0_2_data_119;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_120 <= amplifier_0_0_data_120;
    end else begin
      amplifier_1_2_data_120 <= amplifier_0_2_data_120;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_121 <= amplifier_0_0_data_121;
    end else begin
      amplifier_1_2_data_121 <= amplifier_0_2_data_121;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_122 <= amplifier_0_0_data_122;
    end else begin
      amplifier_1_2_data_122 <= amplifier_0_2_data_122;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_123 <= amplifier_0_0_data_123;
    end else begin
      amplifier_1_2_data_123 <= amplifier_0_2_data_123;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_124 <= amplifier_0_0_data_124;
    end else begin
      amplifier_1_2_data_124 <= amplifier_0_2_data_124;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_125 <= amplifier_0_0_data_125;
    end else begin
      amplifier_1_2_data_125 <= amplifier_0_2_data_125;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_126 <= amplifier_0_0_data_126;
    end else begin
      amplifier_1_2_data_126 <= amplifier_0_2_data_126;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_127 <= amplifier_0_0_data_127;
    end else begin
      amplifier_1_2_data_127 <= amplifier_0_2_data_127;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_128 <= amplifier_0_0_data_128;
    end else begin
      amplifier_1_2_data_128 <= amplifier_0_2_data_128;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_129 <= amplifier_0_0_data_129;
    end else begin
      amplifier_1_2_data_129 <= amplifier_0_2_data_129;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_130 <= amplifier_0_0_data_130;
    end else begin
      amplifier_1_2_data_130 <= amplifier_0_2_data_130;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_131 <= amplifier_0_0_data_131;
    end else begin
      amplifier_1_2_data_131 <= amplifier_0_2_data_131;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_132 <= amplifier_0_0_data_132;
    end else begin
      amplifier_1_2_data_132 <= amplifier_0_2_data_132;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_133 <= amplifier_0_0_data_133;
    end else begin
      amplifier_1_2_data_133 <= amplifier_0_2_data_133;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_134 <= amplifier_0_0_data_134;
    end else begin
      amplifier_1_2_data_134 <= amplifier_0_2_data_134;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_135 <= amplifier_0_0_data_135;
    end else begin
      amplifier_1_2_data_135 <= amplifier_0_2_data_135;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_136 <= amplifier_0_0_data_136;
    end else begin
      amplifier_1_2_data_136 <= amplifier_0_2_data_136;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_137 <= amplifier_0_0_data_137;
    end else begin
      amplifier_1_2_data_137 <= amplifier_0_2_data_137;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_138 <= amplifier_0_0_data_138;
    end else begin
      amplifier_1_2_data_138 <= amplifier_0_2_data_138;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_139 <= amplifier_0_0_data_139;
    end else begin
      amplifier_1_2_data_139 <= amplifier_0_2_data_139;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_140 <= amplifier_0_0_data_140;
    end else begin
      amplifier_1_2_data_140 <= amplifier_0_2_data_140;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_141 <= amplifier_0_0_data_141;
    end else begin
      amplifier_1_2_data_141 <= amplifier_0_2_data_141;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_142 <= amplifier_0_0_data_142;
    end else begin
      amplifier_1_2_data_142 <= amplifier_0_2_data_142;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_143 <= amplifier_0_0_data_143;
    end else begin
      amplifier_1_2_data_143 <= amplifier_0_2_data_143;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_144 <= amplifier_0_0_data_144;
    end else begin
      amplifier_1_2_data_144 <= amplifier_0_2_data_144;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_145 <= amplifier_0_0_data_145;
    end else begin
      amplifier_1_2_data_145 <= amplifier_0_2_data_145;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_146 <= amplifier_0_0_data_146;
    end else begin
      amplifier_1_2_data_146 <= amplifier_0_2_data_146;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_147 <= amplifier_0_0_data_147;
    end else begin
      amplifier_1_2_data_147 <= amplifier_0_2_data_147;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_148 <= amplifier_0_0_data_148;
    end else begin
      amplifier_1_2_data_148 <= amplifier_0_2_data_148;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_149 <= amplifier_0_0_data_149;
    end else begin
      amplifier_1_2_data_149 <= amplifier_0_2_data_149;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_150 <= amplifier_0_0_data_150;
    end else begin
      amplifier_1_2_data_150 <= amplifier_0_2_data_150;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_151 <= amplifier_0_0_data_151;
    end else begin
      amplifier_1_2_data_151 <= amplifier_0_2_data_151;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_152 <= amplifier_0_0_data_152;
    end else begin
      amplifier_1_2_data_152 <= amplifier_0_2_data_152;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_153 <= amplifier_0_0_data_153;
    end else begin
      amplifier_1_2_data_153 <= amplifier_0_2_data_153;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_154 <= amplifier_0_0_data_154;
    end else begin
      amplifier_1_2_data_154 <= amplifier_0_2_data_154;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_155 <= amplifier_0_0_data_155;
    end else begin
      amplifier_1_2_data_155 <= amplifier_0_2_data_155;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_156 <= amplifier_0_0_data_156;
    end else begin
      amplifier_1_2_data_156 <= amplifier_0_2_data_156;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_157 <= amplifier_0_0_data_157;
    end else begin
      amplifier_1_2_data_157 <= amplifier_0_2_data_157;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_158 <= amplifier_0_0_data_158;
    end else begin
      amplifier_1_2_data_158 <= amplifier_0_2_data_158;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_159 <= amplifier_0_0_data_159;
    end else begin
      amplifier_1_2_data_159 <= amplifier_0_2_data_159;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_160 <= amplifier_0_0_data_160;
    end else begin
      amplifier_1_2_data_160 <= amplifier_0_2_data_160;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_161 <= amplifier_0_0_data_161;
    end else begin
      amplifier_1_2_data_161 <= amplifier_0_2_data_161;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_162 <= amplifier_0_0_data_162;
    end else begin
      amplifier_1_2_data_162 <= amplifier_0_2_data_162;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_163 <= amplifier_0_0_data_163;
    end else begin
      amplifier_1_2_data_163 <= amplifier_0_2_data_163;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_164 <= amplifier_0_0_data_164;
    end else begin
      amplifier_1_2_data_164 <= amplifier_0_2_data_164;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_165 <= amplifier_0_0_data_165;
    end else begin
      amplifier_1_2_data_165 <= amplifier_0_2_data_165;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_166 <= amplifier_0_0_data_166;
    end else begin
      amplifier_1_2_data_166 <= amplifier_0_2_data_166;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_167 <= amplifier_0_0_data_167;
    end else begin
      amplifier_1_2_data_167 <= amplifier_0_2_data_167;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_168 <= amplifier_0_0_data_168;
    end else begin
      amplifier_1_2_data_168 <= amplifier_0_2_data_168;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_169 <= amplifier_0_0_data_169;
    end else begin
      amplifier_1_2_data_169 <= amplifier_0_2_data_169;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_170 <= amplifier_0_0_data_170;
    end else begin
      amplifier_1_2_data_170 <= amplifier_0_2_data_170;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_171 <= amplifier_0_0_data_171;
    end else begin
      amplifier_1_2_data_171 <= amplifier_0_2_data_171;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_172 <= amplifier_0_0_data_172;
    end else begin
      amplifier_1_2_data_172 <= amplifier_0_2_data_172;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_173 <= amplifier_0_0_data_173;
    end else begin
      amplifier_1_2_data_173 <= amplifier_0_2_data_173;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_174 <= amplifier_0_0_data_174;
    end else begin
      amplifier_1_2_data_174 <= amplifier_0_2_data_174;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_175 <= amplifier_0_0_data_175;
    end else begin
      amplifier_1_2_data_175 <= amplifier_0_2_data_175;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_176 <= amplifier_0_0_data_176;
    end else begin
      amplifier_1_2_data_176 <= amplifier_0_2_data_176;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_177 <= amplifier_0_0_data_177;
    end else begin
      amplifier_1_2_data_177 <= amplifier_0_2_data_177;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_178 <= amplifier_0_0_data_178;
    end else begin
      amplifier_1_2_data_178 <= amplifier_0_2_data_178;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_179 <= amplifier_0_0_data_179;
    end else begin
      amplifier_1_2_data_179 <= amplifier_0_2_data_179;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_180 <= amplifier_0_0_data_180;
    end else begin
      amplifier_1_2_data_180 <= amplifier_0_2_data_180;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_181 <= amplifier_0_0_data_181;
    end else begin
      amplifier_1_2_data_181 <= amplifier_0_2_data_181;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_182 <= amplifier_0_0_data_182;
    end else begin
      amplifier_1_2_data_182 <= amplifier_0_2_data_182;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_183 <= amplifier_0_0_data_183;
    end else begin
      amplifier_1_2_data_183 <= amplifier_0_2_data_183;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_184 <= amplifier_0_0_data_184;
    end else begin
      amplifier_1_2_data_184 <= amplifier_0_2_data_184;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_185 <= amplifier_0_0_data_185;
    end else begin
      amplifier_1_2_data_185 <= amplifier_0_2_data_185;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_186 <= amplifier_0_0_data_186;
    end else begin
      amplifier_1_2_data_186 <= amplifier_0_2_data_186;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_187 <= amplifier_0_0_data_187;
    end else begin
      amplifier_1_2_data_187 <= amplifier_0_2_data_187;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_188 <= amplifier_0_0_data_188;
    end else begin
      amplifier_1_2_data_188 <= amplifier_0_2_data_188;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_189 <= amplifier_0_0_data_189;
    end else begin
      amplifier_1_2_data_189 <= amplifier_0_2_data_189;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_190 <= amplifier_0_0_data_190;
    end else begin
      amplifier_1_2_data_190 <= amplifier_0_2_data_190;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_191 <= amplifier_0_0_data_191;
    end else begin
      amplifier_1_2_data_191 <= amplifier_0_2_data_191;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_192 <= amplifier_0_0_data_192;
    end else begin
      amplifier_1_2_data_192 <= amplifier_0_2_data_192;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_193 <= amplifier_0_0_data_193;
    end else begin
      amplifier_1_2_data_193 <= amplifier_0_2_data_193;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_194 <= amplifier_0_0_data_194;
    end else begin
      amplifier_1_2_data_194 <= amplifier_0_2_data_194;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_195 <= amplifier_0_0_data_195;
    end else begin
      amplifier_1_2_data_195 <= amplifier_0_2_data_195;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_196 <= amplifier_0_0_data_196;
    end else begin
      amplifier_1_2_data_196 <= amplifier_0_2_data_196;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_197 <= amplifier_0_0_data_197;
    end else begin
      amplifier_1_2_data_197 <= amplifier_0_2_data_197;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_198 <= amplifier_0_0_data_198;
    end else begin
      amplifier_1_2_data_198 <= amplifier_0_2_data_198;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_199 <= amplifier_0_0_data_199;
    end else begin
      amplifier_1_2_data_199 <= amplifier_0_2_data_199;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_200 <= amplifier_0_0_data_200;
    end else begin
      amplifier_1_2_data_200 <= amplifier_0_2_data_200;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_201 <= amplifier_0_0_data_201;
    end else begin
      amplifier_1_2_data_201 <= amplifier_0_2_data_201;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_202 <= amplifier_0_0_data_202;
    end else begin
      amplifier_1_2_data_202 <= amplifier_0_2_data_202;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_203 <= amplifier_0_0_data_203;
    end else begin
      amplifier_1_2_data_203 <= amplifier_0_2_data_203;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_204 <= amplifier_0_0_data_204;
    end else begin
      amplifier_1_2_data_204 <= amplifier_0_2_data_204;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_205 <= amplifier_0_0_data_205;
    end else begin
      amplifier_1_2_data_205 <= amplifier_0_2_data_205;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_206 <= amplifier_0_0_data_206;
    end else begin
      amplifier_1_2_data_206 <= amplifier_0_2_data_206;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_207 <= amplifier_0_0_data_207;
    end else begin
      amplifier_1_2_data_207 <= amplifier_0_2_data_207;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_208 <= amplifier_0_0_data_208;
    end else begin
      amplifier_1_2_data_208 <= amplifier_0_2_data_208;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_209 <= amplifier_0_0_data_209;
    end else begin
      amplifier_1_2_data_209 <= amplifier_0_2_data_209;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_210 <= amplifier_0_0_data_210;
    end else begin
      amplifier_1_2_data_210 <= amplifier_0_2_data_210;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_211 <= amplifier_0_0_data_211;
    end else begin
      amplifier_1_2_data_211 <= amplifier_0_2_data_211;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_212 <= amplifier_0_0_data_212;
    end else begin
      amplifier_1_2_data_212 <= amplifier_0_2_data_212;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_213 <= amplifier_0_0_data_213;
    end else begin
      amplifier_1_2_data_213 <= amplifier_0_2_data_213;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_214 <= amplifier_0_0_data_214;
    end else begin
      amplifier_1_2_data_214 <= amplifier_0_2_data_214;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_215 <= amplifier_0_0_data_215;
    end else begin
      amplifier_1_2_data_215 <= amplifier_0_2_data_215;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_216 <= amplifier_0_0_data_216;
    end else begin
      amplifier_1_2_data_216 <= amplifier_0_2_data_216;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_217 <= amplifier_0_0_data_217;
    end else begin
      amplifier_1_2_data_217 <= amplifier_0_2_data_217;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_218 <= amplifier_0_0_data_218;
    end else begin
      amplifier_1_2_data_218 <= amplifier_0_2_data_218;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_219 <= amplifier_0_0_data_219;
    end else begin
      amplifier_1_2_data_219 <= amplifier_0_2_data_219;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_220 <= amplifier_0_0_data_220;
    end else begin
      amplifier_1_2_data_220 <= amplifier_0_2_data_220;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_221 <= amplifier_0_0_data_221;
    end else begin
      amplifier_1_2_data_221 <= amplifier_0_2_data_221;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_222 <= amplifier_0_0_data_222;
    end else begin
      amplifier_1_2_data_222 <= amplifier_0_2_data_222;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_223 <= amplifier_0_0_data_223;
    end else begin
      amplifier_1_2_data_223 <= amplifier_0_2_data_223;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_224 <= amplifier_0_0_data_224;
    end else begin
      amplifier_1_2_data_224 <= amplifier_0_2_data_224;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_225 <= amplifier_0_0_data_225;
    end else begin
      amplifier_1_2_data_225 <= amplifier_0_2_data_225;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_226 <= amplifier_0_0_data_226;
    end else begin
      amplifier_1_2_data_226 <= amplifier_0_2_data_226;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_227 <= amplifier_0_0_data_227;
    end else begin
      amplifier_1_2_data_227 <= amplifier_0_2_data_227;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_228 <= amplifier_0_0_data_228;
    end else begin
      amplifier_1_2_data_228 <= amplifier_0_2_data_228;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_229 <= amplifier_0_0_data_229;
    end else begin
      amplifier_1_2_data_229 <= amplifier_0_2_data_229;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_230 <= amplifier_0_0_data_230;
    end else begin
      amplifier_1_2_data_230 <= amplifier_0_2_data_230;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_231 <= amplifier_0_0_data_231;
    end else begin
      amplifier_1_2_data_231 <= amplifier_0_2_data_231;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_232 <= amplifier_0_0_data_232;
    end else begin
      amplifier_1_2_data_232 <= amplifier_0_2_data_232;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_233 <= amplifier_0_0_data_233;
    end else begin
      amplifier_1_2_data_233 <= amplifier_0_2_data_233;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_234 <= amplifier_0_0_data_234;
    end else begin
      amplifier_1_2_data_234 <= amplifier_0_2_data_234;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_235 <= amplifier_0_0_data_235;
    end else begin
      amplifier_1_2_data_235 <= amplifier_0_2_data_235;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_236 <= amplifier_0_0_data_236;
    end else begin
      amplifier_1_2_data_236 <= amplifier_0_2_data_236;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_237 <= amplifier_0_0_data_237;
    end else begin
      amplifier_1_2_data_237 <= amplifier_0_2_data_237;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_238 <= amplifier_0_0_data_238;
    end else begin
      amplifier_1_2_data_238 <= amplifier_0_2_data_238;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_239 <= amplifier_0_0_data_239;
    end else begin
      amplifier_1_2_data_239 <= amplifier_0_2_data_239;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_240 <= amplifier_0_0_data_240;
    end else begin
      amplifier_1_2_data_240 <= amplifier_0_2_data_240;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_241 <= amplifier_0_0_data_241;
    end else begin
      amplifier_1_2_data_241 <= amplifier_0_2_data_241;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_242 <= amplifier_0_0_data_242;
    end else begin
      amplifier_1_2_data_242 <= amplifier_0_2_data_242;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_243 <= amplifier_0_0_data_243;
    end else begin
      amplifier_1_2_data_243 <= amplifier_0_2_data_243;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_244 <= amplifier_0_0_data_244;
    end else begin
      amplifier_1_2_data_244 <= amplifier_0_2_data_244;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_245 <= amplifier_0_0_data_245;
    end else begin
      amplifier_1_2_data_245 <= amplifier_0_2_data_245;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_246 <= amplifier_0_0_data_246;
    end else begin
      amplifier_1_2_data_246 <= amplifier_0_2_data_246;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_247 <= amplifier_0_0_data_247;
    end else begin
      amplifier_1_2_data_247 <= amplifier_0_2_data_247;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_248 <= amplifier_0_0_data_248;
    end else begin
      amplifier_1_2_data_248 <= amplifier_0_2_data_248;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_249 <= amplifier_0_0_data_249;
    end else begin
      amplifier_1_2_data_249 <= amplifier_0_2_data_249;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_250 <= amplifier_0_0_data_250;
    end else begin
      amplifier_1_2_data_250 <= amplifier_0_2_data_250;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_251 <= amplifier_0_0_data_251;
    end else begin
      amplifier_1_2_data_251 <= amplifier_0_2_data_251;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_252 <= amplifier_0_0_data_252;
    end else begin
      amplifier_1_2_data_252 <= amplifier_0_2_data_252;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_253 <= amplifier_0_0_data_253;
    end else begin
      amplifier_1_2_data_253 <= amplifier_0_2_data_253;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_254 <= amplifier_0_0_data_254;
    end else begin
      amplifier_1_2_data_254 <= amplifier_0_2_data_254;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_data_255 <= amplifier_0_0_data_255;
    end else begin
      amplifier_1_2_data_255 <= amplifier_0_2_data_255;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_header_0 <= amplifier_0_0_header_0;
    end else begin
      amplifier_1_2_header_0 <= amplifier_0_2_header_0;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_header_1 <= amplifier_0_0_header_1;
    end else begin
      amplifier_1_2_header_1 <= amplifier_0_2_header_1;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_header_2 <= amplifier_0_0_header_2;
    end else begin
      amplifier_1_2_header_2 <= amplifier_0_2_header_2;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_header_3 <= amplifier_0_0_header_3;
    end else begin
      amplifier_1_2_header_3 <= amplifier_0_2_header_3;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_header_4 <= amplifier_0_0_header_4;
    end else begin
      amplifier_1_2_header_4 <= amplifier_0_2_header_4;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_header_5 <= amplifier_0_0_header_5;
    end else begin
      amplifier_1_2_header_5 <= amplifier_0_2_header_5;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_header_6 <= amplifier_0_0_header_6;
    end else begin
      amplifier_1_2_header_6 <= amplifier_0_2_header_6;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_header_7 <= amplifier_0_0_header_7;
    end else begin
      amplifier_1_2_header_7 <= amplifier_0_2_header_7;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_header_8 <= amplifier_0_0_header_8;
    end else begin
      amplifier_1_2_header_8 <= amplifier_0_2_header_8;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_header_9 <= amplifier_0_0_header_9;
    end else begin
      amplifier_1_2_header_9 <= amplifier_0_2_header_9;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_header_10 <= amplifier_0_0_header_10;
    end else begin
      amplifier_1_2_header_10 <= amplifier_0_2_header_10;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_header_11 <= amplifier_0_0_header_11;
    end else begin
      amplifier_1_2_header_11 <= amplifier_0_2_header_11;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_header_12 <= amplifier_0_0_header_12;
    end else begin
      amplifier_1_2_header_12 <= amplifier_0_2_header_12;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_header_13 <= amplifier_0_0_header_13;
    end else begin
      amplifier_1_2_header_13 <= amplifier_0_2_header_13;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_header_14 <= amplifier_0_0_header_14;
    end else begin
      amplifier_1_2_header_14 <= amplifier_0_2_header_14;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_header_15 <= amplifier_0_0_header_15;
    end else begin
      amplifier_1_2_header_15 <= amplifier_0_2_header_15;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_parse_current_state <= amplifier_0_0_parse_current_state;
    end else begin
      amplifier_1_2_parse_current_state <= amplifier_0_2_parse_current_state;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_parse_current_offset <= amplifier_0_0_parse_current_offset;
    end else begin
      amplifier_1_2_parse_current_offset <= amplifier_0_2_parse_current_offset;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_parse_transition_field <= amplifier_0_0_parse_transition_field;
    end else begin
      amplifier_1_2_parse_transition_field <= amplifier_0_2_parse_transition_field;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_next_processor_id <= amplifier_0_0_next_processor_id;
    end else begin
      amplifier_1_2_next_processor_id <= amplifier_0_2_next_processor_id;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_next_config_id <= amplifier_0_0_next_config_id;
    end else begin
      amplifier_1_2_next_config_id <= amplifier_0_2_next_config_id;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 141:31]
      amplifier_1_2_is_valid_processor <= amplifier_0_0_is_valid_processor;
    end else begin
      amplifier_1_2_is_valid_processor <= amplifier_0_2_is_valid_processor;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_0 <= amplifier_0_1_data_0;
    end else begin
      amplifier_1_3_data_0 <= amplifier_0_3_data_0;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_1 <= amplifier_0_1_data_1;
    end else begin
      amplifier_1_3_data_1 <= amplifier_0_3_data_1;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_2 <= amplifier_0_1_data_2;
    end else begin
      amplifier_1_3_data_2 <= amplifier_0_3_data_2;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_3 <= amplifier_0_1_data_3;
    end else begin
      amplifier_1_3_data_3 <= amplifier_0_3_data_3;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_4 <= amplifier_0_1_data_4;
    end else begin
      amplifier_1_3_data_4 <= amplifier_0_3_data_4;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_5 <= amplifier_0_1_data_5;
    end else begin
      amplifier_1_3_data_5 <= amplifier_0_3_data_5;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_6 <= amplifier_0_1_data_6;
    end else begin
      amplifier_1_3_data_6 <= amplifier_0_3_data_6;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_7 <= amplifier_0_1_data_7;
    end else begin
      amplifier_1_3_data_7 <= amplifier_0_3_data_7;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_8 <= amplifier_0_1_data_8;
    end else begin
      amplifier_1_3_data_8 <= amplifier_0_3_data_8;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_9 <= amplifier_0_1_data_9;
    end else begin
      amplifier_1_3_data_9 <= amplifier_0_3_data_9;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_10 <= amplifier_0_1_data_10;
    end else begin
      amplifier_1_3_data_10 <= amplifier_0_3_data_10;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_11 <= amplifier_0_1_data_11;
    end else begin
      amplifier_1_3_data_11 <= amplifier_0_3_data_11;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_12 <= amplifier_0_1_data_12;
    end else begin
      amplifier_1_3_data_12 <= amplifier_0_3_data_12;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_13 <= amplifier_0_1_data_13;
    end else begin
      amplifier_1_3_data_13 <= amplifier_0_3_data_13;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_14 <= amplifier_0_1_data_14;
    end else begin
      amplifier_1_3_data_14 <= amplifier_0_3_data_14;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_15 <= amplifier_0_1_data_15;
    end else begin
      amplifier_1_3_data_15 <= amplifier_0_3_data_15;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_16 <= amplifier_0_1_data_16;
    end else begin
      amplifier_1_3_data_16 <= amplifier_0_3_data_16;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_17 <= amplifier_0_1_data_17;
    end else begin
      amplifier_1_3_data_17 <= amplifier_0_3_data_17;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_18 <= amplifier_0_1_data_18;
    end else begin
      amplifier_1_3_data_18 <= amplifier_0_3_data_18;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_19 <= amplifier_0_1_data_19;
    end else begin
      amplifier_1_3_data_19 <= amplifier_0_3_data_19;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_20 <= amplifier_0_1_data_20;
    end else begin
      amplifier_1_3_data_20 <= amplifier_0_3_data_20;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_21 <= amplifier_0_1_data_21;
    end else begin
      amplifier_1_3_data_21 <= amplifier_0_3_data_21;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_22 <= amplifier_0_1_data_22;
    end else begin
      amplifier_1_3_data_22 <= amplifier_0_3_data_22;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_23 <= amplifier_0_1_data_23;
    end else begin
      amplifier_1_3_data_23 <= amplifier_0_3_data_23;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_24 <= amplifier_0_1_data_24;
    end else begin
      amplifier_1_3_data_24 <= amplifier_0_3_data_24;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_25 <= amplifier_0_1_data_25;
    end else begin
      amplifier_1_3_data_25 <= amplifier_0_3_data_25;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_26 <= amplifier_0_1_data_26;
    end else begin
      amplifier_1_3_data_26 <= amplifier_0_3_data_26;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_27 <= amplifier_0_1_data_27;
    end else begin
      amplifier_1_3_data_27 <= amplifier_0_3_data_27;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_28 <= amplifier_0_1_data_28;
    end else begin
      amplifier_1_3_data_28 <= amplifier_0_3_data_28;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_29 <= amplifier_0_1_data_29;
    end else begin
      amplifier_1_3_data_29 <= amplifier_0_3_data_29;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_30 <= amplifier_0_1_data_30;
    end else begin
      amplifier_1_3_data_30 <= amplifier_0_3_data_30;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_31 <= amplifier_0_1_data_31;
    end else begin
      amplifier_1_3_data_31 <= amplifier_0_3_data_31;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_32 <= amplifier_0_1_data_32;
    end else begin
      amplifier_1_3_data_32 <= amplifier_0_3_data_32;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_33 <= amplifier_0_1_data_33;
    end else begin
      amplifier_1_3_data_33 <= amplifier_0_3_data_33;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_34 <= amplifier_0_1_data_34;
    end else begin
      amplifier_1_3_data_34 <= amplifier_0_3_data_34;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_35 <= amplifier_0_1_data_35;
    end else begin
      amplifier_1_3_data_35 <= amplifier_0_3_data_35;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_36 <= amplifier_0_1_data_36;
    end else begin
      amplifier_1_3_data_36 <= amplifier_0_3_data_36;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_37 <= amplifier_0_1_data_37;
    end else begin
      amplifier_1_3_data_37 <= amplifier_0_3_data_37;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_38 <= amplifier_0_1_data_38;
    end else begin
      amplifier_1_3_data_38 <= amplifier_0_3_data_38;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_39 <= amplifier_0_1_data_39;
    end else begin
      amplifier_1_3_data_39 <= amplifier_0_3_data_39;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_40 <= amplifier_0_1_data_40;
    end else begin
      amplifier_1_3_data_40 <= amplifier_0_3_data_40;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_41 <= amplifier_0_1_data_41;
    end else begin
      amplifier_1_3_data_41 <= amplifier_0_3_data_41;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_42 <= amplifier_0_1_data_42;
    end else begin
      amplifier_1_3_data_42 <= amplifier_0_3_data_42;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_43 <= amplifier_0_1_data_43;
    end else begin
      amplifier_1_3_data_43 <= amplifier_0_3_data_43;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_44 <= amplifier_0_1_data_44;
    end else begin
      amplifier_1_3_data_44 <= amplifier_0_3_data_44;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_45 <= amplifier_0_1_data_45;
    end else begin
      amplifier_1_3_data_45 <= amplifier_0_3_data_45;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_46 <= amplifier_0_1_data_46;
    end else begin
      amplifier_1_3_data_46 <= amplifier_0_3_data_46;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_47 <= amplifier_0_1_data_47;
    end else begin
      amplifier_1_3_data_47 <= amplifier_0_3_data_47;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_48 <= amplifier_0_1_data_48;
    end else begin
      amplifier_1_3_data_48 <= amplifier_0_3_data_48;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_49 <= amplifier_0_1_data_49;
    end else begin
      amplifier_1_3_data_49 <= amplifier_0_3_data_49;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_50 <= amplifier_0_1_data_50;
    end else begin
      amplifier_1_3_data_50 <= amplifier_0_3_data_50;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_51 <= amplifier_0_1_data_51;
    end else begin
      amplifier_1_3_data_51 <= amplifier_0_3_data_51;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_52 <= amplifier_0_1_data_52;
    end else begin
      amplifier_1_3_data_52 <= amplifier_0_3_data_52;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_53 <= amplifier_0_1_data_53;
    end else begin
      amplifier_1_3_data_53 <= amplifier_0_3_data_53;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_54 <= amplifier_0_1_data_54;
    end else begin
      amplifier_1_3_data_54 <= amplifier_0_3_data_54;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_55 <= amplifier_0_1_data_55;
    end else begin
      amplifier_1_3_data_55 <= amplifier_0_3_data_55;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_56 <= amplifier_0_1_data_56;
    end else begin
      amplifier_1_3_data_56 <= amplifier_0_3_data_56;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_57 <= amplifier_0_1_data_57;
    end else begin
      amplifier_1_3_data_57 <= amplifier_0_3_data_57;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_58 <= amplifier_0_1_data_58;
    end else begin
      amplifier_1_3_data_58 <= amplifier_0_3_data_58;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_59 <= amplifier_0_1_data_59;
    end else begin
      amplifier_1_3_data_59 <= amplifier_0_3_data_59;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_60 <= amplifier_0_1_data_60;
    end else begin
      amplifier_1_3_data_60 <= amplifier_0_3_data_60;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_61 <= amplifier_0_1_data_61;
    end else begin
      amplifier_1_3_data_61 <= amplifier_0_3_data_61;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_62 <= amplifier_0_1_data_62;
    end else begin
      amplifier_1_3_data_62 <= amplifier_0_3_data_62;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_63 <= amplifier_0_1_data_63;
    end else begin
      amplifier_1_3_data_63 <= amplifier_0_3_data_63;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_64 <= amplifier_0_1_data_64;
    end else begin
      amplifier_1_3_data_64 <= amplifier_0_3_data_64;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_65 <= amplifier_0_1_data_65;
    end else begin
      amplifier_1_3_data_65 <= amplifier_0_3_data_65;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_66 <= amplifier_0_1_data_66;
    end else begin
      amplifier_1_3_data_66 <= amplifier_0_3_data_66;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_67 <= amplifier_0_1_data_67;
    end else begin
      amplifier_1_3_data_67 <= amplifier_0_3_data_67;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_68 <= amplifier_0_1_data_68;
    end else begin
      amplifier_1_3_data_68 <= amplifier_0_3_data_68;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_69 <= amplifier_0_1_data_69;
    end else begin
      amplifier_1_3_data_69 <= amplifier_0_3_data_69;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_70 <= amplifier_0_1_data_70;
    end else begin
      amplifier_1_3_data_70 <= amplifier_0_3_data_70;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_71 <= amplifier_0_1_data_71;
    end else begin
      amplifier_1_3_data_71 <= amplifier_0_3_data_71;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_72 <= amplifier_0_1_data_72;
    end else begin
      amplifier_1_3_data_72 <= amplifier_0_3_data_72;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_73 <= amplifier_0_1_data_73;
    end else begin
      amplifier_1_3_data_73 <= amplifier_0_3_data_73;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_74 <= amplifier_0_1_data_74;
    end else begin
      amplifier_1_3_data_74 <= amplifier_0_3_data_74;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_75 <= amplifier_0_1_data_75;
    end else begin
      amplifier_1_3_data_75 <= amplifier_0_3_data_75;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_76 <= amplifier_0_1_data_76;
    end else begin
      amplifier_1_3_data_76 <= amplifier_0_3_data_76;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_77 <= amplifier_0_1_data_77;
    end else begin
      amplifier_1_3_data_77 <= amplifier_0_3_data_77;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_78 <= amplifier_0_1_data_78;
    end else begin
      amplifier_1_3_data_78 <= amplifier_0_3_data_78;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_79 <= amplifier_0_1_data_79;
    end else begin
      amplifier_1_3_data_79 <= amplifier_0_3_data_79;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_80 <= amplifier_0_1_data_80;
    end else begin
      amplifier_1_3_data_80 <= amplifier_0_3_data_80;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_81 <= amplifier_0_1_data_81;
    end else begin
      amplifier_1_3_data_81 <= amplifier_0_3_data_81;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_82 <= amplifier_0_1_data_82;
    end else begin
      amplifier_1_3_data_82 <= amplifier_0_3_data_82;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_83 <= amplifier_0_1_data_83;
    end else begin
      amplifier_1_3_data_83 <= amplifier_0_3_data_83;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_84 <= amplifier_0_1_data_84;
    end else begin
      amplifier_1_3_data_84 <= amplifier_0_3_data_84;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_85 <= amplifier_0_1_data_85;
    end else begin
      amplifier_1_3_data_85 <= amplifier_0_3_data_85;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_86 <= amplifier_0_1_data_86;
    end else begin
      amplifier_1_3_data_86 <= amplifier_0_3_data_86;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_87 <= amplifier_0_1_data_87;
    end else begin
      amplifier_1_3_data_87 <= amplifier_0_3_data_87;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_88 <= amplifier_0_1_data_88;
    end else begin
      amplifier_1_3_data_88 <= amplifier_0_3_data_88;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_89 <= amplifier_0_1_data_89;
    end else begin
      amplifier_1_3_data_89 <= amplifier_0_3_data_89;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_90 <= amplifier_0_1_data_90;
    end else begin
      amplifier_1_3_data_90 <= amplifier_0_3_data_90;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_91 <= amplifier_0_1_data_91;
    end else begin
      amplifier_1_3_data_91 <= amplifier_0_3_data_91;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_92 <= amplifier_0_1_data_92;
    end else begin
      amplifier_1_3_data_92 <= amplifier_0_3_data_92;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_93 <= amplifier_0_1_data_93;
    end else begin
      amplifier_1_3_data_93 <= amplifier_0_3_data_93;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_94 <= amplifier_0_1_data_94;
    end else begin
      amplifier_1_3_data_94 <= amplifier_0_3_data_94;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_95 <= amplifier_0_1_data_95;
    end else begin
      amplifier_1_3_data_95 <= amplifier_0_3_data_95;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_96 <= amplifier_0_1_data_96;
    end else begin
      amplifier_1_3_data_96 <= amplifier_0_3_data_96;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_97 <= amplifier_0_1_data_97;
    end else begin
      amplifier_1_3_data_97 <= amplifier_0_3_data_97;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_98 <= amplifier_0_1_data_98;
    end else begin
      amplifier_1_3_data_98 <= amplifier_0_3_data_98;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_99 <= amplifier_0_1_data_99;
    end else begin
      amplifier_1_3_data_99 <= amplifier_0_3_data_99;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_100 <= amplifier_0_1_data_100;
    end else begin
      amplifier_1_3_data_100 <= amplifier_0_3_data_100;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_101 <= amplifier_0_1_data_101;
    end else begin
      amplifier_1_3_data_101 <= amplifier_0_3_data_101;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_102 <= amplifier_0_1_data_102;
    end else begin
      amplifier_1_3_data_102 <= amplifier_0_3_data_102;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_103 <= amplifier_0_1_data_103;
    end else begin
      amplifier_1_3_data_103 <= amplifier_0_3_data_103;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_104 <= amplifier_0_1_data_104;
    end else begin
      amplifier_1_3_data_104 <= amplifier_0_3_data_104;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_105 <= amplifier_0_1_data_105;
    end else begin
      amplifier_1_3_data_105 <= amplifier_0_3_data_105;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_106 <= amplifier_0_1_data_106;
    end else begin
      amplifier_1_3_data_106 <= amplifier_0_3_data_106;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_107 <= amplifier_0_1_data_107;
    end else begin
      amplifier_1_3_data_107 <= amplifier_0_3_data_107;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_108 <= amplifier_0_1_data_108;
    end else begin
      amplifier_1_3_data_108 <= amplifier_0_3_data_108;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_109 <= amplifier_0_1_data_109;
    end else begin
      amplifier_1_3_data_109 <= amplifier_0_3_data_109;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_110 <= amplifier_0_1_data_110;
    end else begin
      amplifier_1_3_data_110 <= amplifier_0_3_data_110;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_111 <= amplifier_0_1_data_111;
    end else begin
      amplifier_1_3_data_111 <= amplifier_0_3_data_111;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_112 <= amplifier_0_1_data_112;
    end else begin
      amplifier_1_3_data_112 <= amplifier_0_3_data_112;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_113 <= amplifier_0_1_data_113;
    end else begin
      amplifier_1_3_data_113 <= amplifier_0_3_data_113;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_114 <= amplifier_0_1_data_114;
    end else begin
      amplifier_1_3_data_114 <= amplifier_0_3_data_114;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_115 <= amplifier_0_1_data_115;
    end else begin
      amplifier_1_3_data_115 <= amplifier_0_3_data_115;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_116 <= amplifier_0_1_data_116;
    end else begin
      amplifier_1_3_data_116 <= amplifier_0_3_data_116;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_117 <= amplifier_0_1_data_117;
    end else begin
      amplifier_1_3_data_117 <= amplifier_0_3_data_117;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_118 <= amplifier_0_1_data_118;
    end else begin
      amplifier_1_3_data_118 <= amplifier_0_3_data_118;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_119 <= amplifier_0_1_data_119;
    end else begin
      amplifier_1_3_data_119 <= amplifier_0_3_data_119;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_120 <= amplifier_0_1_data_120;
    end else begin
      amplifier_1_3_data_120 <= amplifier_0_3_data_120;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_121 <= amplifier_0_1_data_121;
    end else begin
      amplifier_1_3_data_121 <= amplifier_0_3_data_121;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_122 <= amplifier_0_1_data_122;
    end else begin
      amplifier_1_3_data_122 <= amplifier_0_3_data_122;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_123 <= amplifier_0_1_data_123;
    end else begin
      amplifier_1_3_data_123 <= amplifier_0_3_data_123;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_124 <= amplifier_0_1_data_124;
    end else begin
      amplifier_1_3_data_124 <= amplifier_0_3_data_124;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_125 <= amplifier_0_1_data_125;
    end else begin
      amplifier_1_3_data_125 <= amplifier_0_3_data_125;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_126 <= amplifier_0_1_data_126;
    end else begin
      amplifier_1_3_data_126 <= amplifier_0_3_data_126;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_127 <= amplifier_0_1_data_127;
    end else begin
      amplifier_1_3_data_127 <= amplifier_0_3_data_127;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_128 <= amplifier_0_1_data_128;
    end else begin
      amplifier_1_3_data_128 <= amplifier_0_3_data_128;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_129 <= amplifier_0_1_data_129;
    end else begin
      amplifier_1_3_data_129 <= amplifier_0_3_data_129;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_130 <= amplifier_0_1_data_130;
    end else begin
      amplifier_1_3_data_130 <= amplifier_0_3_data_130;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_131 <= amplifier_0_1_data_131;
    end else begin
      amplifier_1_3_data_131 <= amplifier_0_3_data_131;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_132 <= amplifier_0_1_data_132;
    end else begin
      amplifier_1_3_data_132 <= amplifier_0_3_data_132;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_133 <= amplifier_0_1_data_133;
    end else begin
      amplifier_1_3_data_133 <= amplifier_0_3_data_133;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_134 <= amplifier_0_1_data_134;
    end else begin
      amplifier_1_3_data_134 <= amplifier_0_3_data_134;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_135 <= amplifier_0_1_data_135;
    end else begin
      amplifier_1_3_data_135 <= amplifier_0_3_data_135;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_136 <= amplifier_0_1_data_136;
    end else begin
      amplifier_1_3_data_136 <= amplifier_0_3_data_136;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_137 <= amplifier_0_1_data_137;
    end else begin
      amplifier_1_3_data_137 <= amplifier_0_3_data_137;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_138 <= amplifier_0_1_data_138;
    end else begin
      amplifier_1_3_data_138 <= amplifier_0_3_data_138;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_139 <= amplifier_0_1_data_139;
    end else begin
      amplifier_1_3_data_139 <= amplifier_0_3_data_139;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_140 <= amplifier_0_1_data_140;
    end else begin
      amplifier_1_3_data_140 <= amplifier_0_3_data_140;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_141 <= amplifier_0_1_data_141;
    end else begin
      amplifier_1_3_data_141 <= amplifier_0_3_data_141;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_142 <= amplifier_0_1_data_142;
    end else begin
      amplifier_1_3_data_142 <= amplifier_0_3_data_142;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_143 <= amplifier_0_1_data_143;
    end else begin
      amplifier_1_3_data_143 <= amplifier_0_3_data_143;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_144 <= amplifier_0_1_data_144;
    end else begin
      amplifier_1_3_data_144 <= amplifier_0_3_data_144;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_145 <= amplifier_0_1_data_145;
    end else begin
      amplifier_1_3_data_145 <= amplifier_0_3_data_145;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_146 <= amplifier_0_1_data_146;
    end else begin
      amplifier_1_3_data_146 <= amplifier_0_3_data_146;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_147 <= amplifier_0_1_data_147;
    end else begin
      amplifier_1_3_data_147 <= amplifier_0_3_data_147;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_148 <= amplifier_0_1_data_148;
    end else begin
      amplifier_1_3_data_148 <= amplifier_0_3_data_148;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_149 <= amplifier_0_1_data_149;
    end else begin
      amplifier_1_3_data_149 <= amplifier_0_3_data_149;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_150 <= amplifier_0_1_data_150;
    end else begin
      amplifier_1_3_data_150 <= amplifier_0_3_data_150;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_151 <= amplifier_0_1_data_151;
    end else begin
      amplifier_1_3_data_151 <= amplifier_0_3_data_151;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_152 <= amplifier_0_1_data_152;
    end else begin
      amplifier_1_3_data_152 <= amplifier_0_3_data_152;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_153 <= amplifier_0_1_data_153;
    end else begin
      amplifier_1_3_data_153 <= amplifier_0_3_data_153;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_154 <= amplifier_0_1_data_154;
    end else begin
      amplifier_1_3_data_154 <= amplifier_0_3_data_154;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_155 <= amplifier_0_1_data_155;
    end else begin
      amplifier_1_3_data_155 <= amplifier_0_3_data_155;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_156 <= amplifier_0_1_data_156;
    end else begin
      amplifier_1_3_data_156 <= amplifier_0_3_data_156;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_157 <= amplifier_0_1_data_157;
    end else begin
      amplifier_1_3_data_157 <= amplifier_0_3_data_157;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_158 <= amplifier_0_1_data_158;
    end else begin
      amplifier_1_3_data_158 <= amplifier_0_3_data_158;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_159 <= amplifier_0_1_data_159;
    end else begin
      amplifier_1_3_data_159 <= amplifier_0_3_data_159;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_160 <= amplifier_0_1_data_160;
    end else begin
      amplifier_1_3_data_160 <= amplifier_0_3_data_160;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_161 <= amplifier_0_1_data_161;
    end else begin
      amplifier_1_3_data_161 <= amplifier_0_3_data_161;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_162 <= amplifier_0_1_data_162;
    end else begin
      amplifier_1_3_data_162 <= amplifier_0_3_data_162;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_163 <= amplifier_0_1_data_163;
    end else begin
      amplifier_1_3_data_163 <= amplifier_0_3_data_163;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_164 <= amplifier_0_1_data_164;
    end else begin
      amplifier_1_3_data_164 <= amplifier_0_3_data_164;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_165 <= amplifier_0_1_data_165;
    end else begin
      amplifier_1_3_data_165 <= amplifier_0_3_data_165;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_166 <= amplifier_0_1_data_166;
    end else begin
      amplifier_1_3_data_166 <= amplifier_0_3_data_166;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_167 <= amplifier_0_1_data_167;
    end else begin
      amplifier_1_3_data_167 <= amplifier_0_3_data_167;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_168 <= amplifier_0_1_data_168;
    end else begin
      amplifier_1_3_data_168 <= amplifier_0_3_data_168;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_169 <= amplifier_0_1_data_169;
    end else begin
      amplifier_1_3_data_169 <= amplifier_0_3_data_169;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_170 <= amplifier_0_1_data_170;
    end else begin
      amplifier_1_3_data_170 <= amplifier_0_3_data_170;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_171 <= amplifier_0_1_data_171;
    end else begin
      amplifier_1_3_data_171 <= amplifier_0_3_data_171;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_172 <= amplifier_0_1_data_172;
    end else begin
      amplifier_1_3_data_172 <= amplifier_0_3_data_172;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_173 <= amplifier_0_1_data_173;
    end else begin
      amplifier_1_3_data_173 <= amplifier_0_3_data_173;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_174 <= amplifier_0_1_data_174;
    end else begin
      amplifier_1_3_data_174 <= amplifier_0_3_data_174;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_175 <= amplifier_0_1_data_175;
    end else begin
      amplifier_1_3_data_175 <= amplifier_0_3_data_175;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_176 <= amplifier_0_1_data_176;
    end else begin
      amplifier_1_3_data_176 <= amplifier_0_3_data_176;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_177 <= amplifier_0_1_data_177;
    end else begin
      amplifier_1_3_data_177 <= amplifier_0_3_data_177;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_178 <= amplifier_0_1_data_178;
    end else begin
      amplifier_1_3_data_178 <= amplifier_0_3_data_178;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_179 <= amplifier_0_1_data_179;
    end else begin
      amplifier_1_3_data_179 <= amplifier_0_3_data_179;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_180 <= amplifier_0_1_data_180;
    end else begin
      amplifier_1_3_data_180 <= amplifier_0_3_data_180;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_181 <= amplifier_0_1_data_181;
    end else begin
      amplifier_1_3_data_181 <= amplifier_0_3_data_181;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_182 <= amplifier_0_1_data_182;
    end else begin
      amplifier_1_3_data_182 <= amplifier_0_3_data_182;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_183 <= amplifier_0_1_data_183;
    end else begin
      amplifier_1_3_data_183 <= amplifier_0_3_data_183;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_184 <= amplifier_0_1_data_184;
    end else begin
      amplifier_1_3_data_184 <= amplifier_0_3_data_184;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_185 <= amplifier_0_1_data_185;
    end else begin
      amplifier_1_3_data_185 <= amplifier_0_3_data_185;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_186 <= amplifier_0_1_data_186;
    end else begin
      amplifier_1_3_data_186 <= amplifier_0_3_data_186;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_187 <= amplifier_0_1_data_187;
    end else begin
      amplifier_1_3_data_187 <= amplifier_0_3_data_187;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_188 <= amplifier_0_1_data_188;
    end else begin
      amplifier_1_3_data_188 <= amplifier_0_3_data_188;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_189 <= amplifier_0_1_data_189;
    end else begin
      amplifier_1_3_data_189 <= amplifier_0_3_data_189;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_190 <= amplifier_0_1_data_190;
    end else begin
      amplifier_1_3_data_190 <= amplifier_0_3_data_190;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_191 <= amplifier_0_1_data_191;
    end else begin
      amplifier_1_3_data_191 <= amplifier_0_3_data_191;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_192 <= amplifier_0_1_data_192;
    end else begin
      amplifier_1_3_data_192 <= amplifier_0_3_data_192;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_193 <= amplifier_0_1_data_193;
    end else begin
      amplifier_1_3_data_193 <= amplifier_0_3_data_193;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_194 <= amplifier_0_1_data_194;
    end else begin
      amplifier_1_3_data_194 <= amplifier_0_3_data_194;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_195 <= amplifier_0_1_data_195;
    end else begin
      amplifier_1_3_data_195 <= amplifier_0_3_data_195;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_196 <= amplifier_0_1_data_196;
    end else begin
      amplifier_1_3_data_196 <= amplifier_0_3_data_196;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_197 <= amplifier_0_1_data_197;
    end else begin
      amplifier_1_3_data_197 <= amplifier_0_3_data_197;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_198 <= amplifier_0_1_data_198;
    end else begin
      amplifier_1_3_data_198 <= amplifier_0_3_data_198;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_199 <= amplifier_0_1_data_199;
    end else begin
      amplifier_1_3_data_199 <= amplifier_0_3_data_199;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_200 <= amplifier_0_1_data_200;
    end else begin
      amplifier_1_3_data_200 <= amplifier_0_3_data_200;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_201 <= amplifier_0_1_data_201;
    end else begin
      amplifier_1_3_data_201 <= amplifier_0_3_data_201;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_202 <= amplifier_0_1_data_202;
    end else begin
      amplifier_1_3_data_202 <= amplifier_0_3_data_202;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_203 <= amplifier_0_1_data_203;
    end else begin
      amplifier_1_3_data_203 <= amplifier_0_3_data_203;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_204 <= amplifier_0_1_data_204;
    end else begin
      amplifier_1_3_data_204 <= amplifier_0_3_data_204;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_205 <= amplifier_0_1_data_205;
    end else begin
      amplifier_1_3_data_205 <= amplifier_0_3_data_205;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_206 <= amplifier_0_1_data_206;
    end else begin
      amplifier_1_3_data_206 <= amplifier_0_3_data_206;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_207 <= amplifier_0_1_data_207;
    end else begin
      amplifier_1_3_data_207 <= amplifier_0_3_data_207;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_208 <= amplifier_0_1_data_208;
    end else begin
      amplifier_1_3_data_208 <= amplifier_0_3_data_208;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_209 <= amplifier_0_1_data_209;
    end else begin
      amplifier_1_3_data_209 <= amplifier_0_3_data_209;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_210 <= amplifier_0_1_data_210;
    end else begin
      amplifier_1_3_data_210 <= amplifier_0_3_data_210;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_211 <= amplifier_0_1_data_211;
    end else begin
      amplifier_1_3_data_211 <= amplifier_0_3_data_211;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_212 <= amplifier_0_1_data_212;
    end else begin
      amplifier_1_3_data_212 <= amplifier_0_3_data_212;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_213 <= amplifier_0_1_data_213;
    end else begin
      amplifier_1_3_data_213 <= amplifier_0_3_data_213;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_214 <= amplifier_0_1_data_214;
    end else begin
      amplifier_1_3_data_214 <= amplifier_0_3_data_214;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_215 <= amplifier_0_1_data_215;
    end else begin
      amplifier_1_3_data_215 <= amplifier_0_3_data_215;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_216 <= amplifier_0_1_data_216;
    end else begin
      amplifier_1_3_data_216 <= amplifier_0_3_data_216;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_217 <= amplifier_0_1_data_217;
    end else begin
      amplifier_1_3_data_217 <= amplifier_0_3_data_217;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_218 <= amplifier_0_1_data_218;
    end else begin
      amplifier_1_3_data_218 <= amplifier_0_3_data_218;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_219 <= amplifier_0_1_data_219;
    end else begin
      amplifier_1_3_data_219 <= amplifier_0_3_data_219;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_220 <= amplifier_0_1_data_220;
    end else begin
      amplifier_1_3_data_220 <= amplifier_0_3_data_220;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_221 <= amplifier_0_1_data_221;
    end else begin
      amplifier_1_3_data_221 <= amplifier_0_3_data_221;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_222 <= amplifier_0_1_data_222;
    end else begin
      amplifier_1_3_data_222 <= amplifier_0_3_data_222;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_223 <= amplifier_0_1_data_223;
    end else begin
      amplifier_1_3_data_223 <= amplifier_0_3_data_223;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_224 <= amplifier_0_1_data_224;
    end else begin
      amplifier_1_3_data_224 <= amplifier_0_3_data_224;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_225 <= amplifier_0_1_data_225;
    end else begin
      amplifier_1_3_data_225 <= amplifier_0_3_data_225;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_226 <= amplifier_0_1_data_226;
    end else begin
      amplifier_1_3_data_226 <= amplifier_0_3_data_226;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_227 <= amplifier_0_1_data_227;
    end else begin
      amplifier_1_3_data_227 <= amplifier_0_3_data_227;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_228 <= amplifier_0_1_data_228;
    end else begin
      amplifier_1_3_data_228 <= amplifier_0_3_data_228;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_229 <= amplifier_0_1_data_229;
    end else begin
      amplifier_1_3_data_229 <= amplifier_0_3_data_229;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_230 <= amplifier_0_1_data_230;
    end else begin
      amplifier_1_3_data_230 <= amplifier_0_3_data_230;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_231 <= amplifier_0_1_data_231;
    end else begin
      amplifier_1_3_data_231 <= amplifier_0_3_data_231;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_232 <= amplifier_0_1_data_232;
    end else begin
      amplifier_1_3_data_232 <= amplifier_0_3_data_232;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_233 <= amplifier_0_1_data_233;
    end else begin
      amplifier_1_3_data_233 <= amplifier_0_3_data_233;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_234 <= amplifier_0_1_data_234;
    end else begin
      amplifier_1_3_data_234 <= amplifier_0_3_data_234;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_235 <= amplifier_0_1_data_235;
    end else begin
      amplifier_1_3_data_235 <= amplifier_0_3_data_235;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_236 <= amplifier_0_1_data_236;
    end else begin
      amplifier_1_3_data_236 <= amplifier_0_3_data_236;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_237 <= amplifier_0_1_data_237;
    end else begin
      amplifier_1_3_data_237 <= amplifier_0_3_data_237;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_238 <= amplifier_0_1_data_238;
    end else begin
      amplifier_1_3_data_238 <= amplifier_0_3_data_238;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_239 <= amplifier_0_1_data_239;
    end else begin
      amplifier_1_3_data_239 <= amplifier_0_3_data_239;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_240 <= amplifier_0_1_data_240;
    end else begin
      amplifier_1_3_data_240 <= amplifier_0_3_data_240;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_241 <= amplifier_0_1_data_241;
    end else begin
      amplifier_1_3_data_241 <= amplifier_0_3_data_241;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_242 <= amplifier_0_1_data_242;
    end else begin
      amplifier_1_3_data_242 <= amplifier_0_3_data_242;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_243 <= amplifier_0_1_data_243;
    end else begin
      amplifier_1_3_data_243 <= amplifier_0_3_data_243;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_244 <= amplifier_0_1_data_244;
    end else begin
      amplifier_1_3_data_244 <= amplifier_0_3_data_244;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_245 <= amplifier_0_1_data_245;
    end else begin
      amplifier_1_3_data_245 <= amplifier_0_3_data_245;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_246 <= amplifier_0_1_data_246;
    end else begin
      amplifier_1_3_data_246 <= amplifier_0_3_data_246;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_247 <= amplifier_0_1_data_247;
    end else begin
      amplifier_1_3_data_247 <= amplifier_0_3_data_247;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_248 <= amplifier_0_1_data_248;
    end else begin
      amplifier_1_3_data_248 <= amplifier_0_3_data_248;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_249 <= amplifier_0_1_data_249;
    end else begin
      amplifier_1_3_data_249 <= amplifier_0_3_data_249;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_250 <= amplifier_0_1_data_250;
    end else begin
      amplifier_1_3_data_250 <= amplifier_0_3_data_250;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_251 <= amplifier_0_1_data_251;
    end else begin
      amplifier_1_3_data_251 <= amplifier_0_3_data_251;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_252 <= amplifier_0_1_data_252;
    end else begin
      amplifier_1_3_data_252 <= amplifier_0_3_data_252;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_253 <= amplifier_0_1_data_253;
    end else begin
      amplifier_1_3_data_253 <= amplifier_0_3_data_253;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_254 <= amplifier_0_1_data_254;
    end else begin
      amplifier_1_3_data_254 <= amplifier_0_3_data_254;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_data_255 <= amplifier_0_1_data_255;
    end else begin
      amplifier_1_3_data_255 <= amplifier_0_3_data_255;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_header_0 <= amplifier_0_1_header_0;
    end else begin
      amplifier_1_3_header_0 <= amplifier_0_3_header_0;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_header_1 <= amplifier_0_1_header_1;
    end else begin
      amplifier_1_3_header_1 <= amplifier_0_3_header_1;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_header_2 <= amplifier_0_1_header_2;
    end else begin
      amplifier_1_3_header_2 <= amplifier_0_3_header_2;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_header_3 <= amplifier_0_1_header_3;
    end else begin
      amplifier_1_3_header_3 <= amplifier_0_3_header_3;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_header_4 <= amplifier_0_1_header_4;
    end else begin
      amplifier_1_3_header_4 <= amplifier_0_3_header_4;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_header_5 <= amplifier_0_1_header_5;
    end else begin
      amplifier_1_3_header_5 <= amplifier_0_3_header_5;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_header_6 <= amplifier_0_1_header_6;
    end else begin
      amplifier_1_3_header_6 <= amplifier_0_3_header_6;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_header_7 <= amplifier_0_1_header_7;
    end else begin
      amplifier_1_3_header_7 <= amplifier_0_3_header_7;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_header_8 <= amplifier_0_1_header_8;
    end else begin
      amplifier_1_3_header_8 <= amplifier_0_3_header_8;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_header_9 <= amplifier_0_1_header_9;
    end else begin
      amplifier_1_3_header_9 <= amplifier_0_3_header_9;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_header_10 <= amplifier_0_1_header_10;
    end else begin
      amplifier_1_3_header_10 <= amplifier_0_3_header_10;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_header_11 <= amplifier_0_1_header_11;
    end else begin
      amplifier_1_3_header_11 <= amplifier_0_3_header_11;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_header_12 <= amplifier_0_1_header_12;
    end else begin
      amplifier_1_3_header_12 <= amplifier_0_3_header_12;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_header_13 <= amplifier_0_1_header_13;
    end else begin
      amplifier_1_3_header_13 <= amplifier_0_3_header_13;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_header_14 <= amplifier_0_1_header_14;
    end else begin
      amplifier_1_3_header_14 <= amplifier_0_3_header_14;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_header_15 <= amplifier_0_1_header_15;
    end else begin
      amplifier_1_3_header_15 <= amplifier_0_3_header_15;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_parse_current_state <= amplifier_0_1_parse_current_state;
    end else begin
      amplifier_1_3_parse_current_state <= amplifier_0_3_parse_current_state;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_parse_current_offset <= amplifier_0_1_parse_current_offset;
    end else begin
      amplifier_1_3_parse_current_offset <= amplifier_0_3_parse_current_offset;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_parse_transition_field <= amplifier_0_1_parse_transition_field;
    end else begin
      amplifier_1_3_parse_transition_field <= amplifier_0_3_parse_transition_field;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_next_processor_id <= amplifier_0_1_next_processor_id;
    end else begin
      amplifier_1_3_next_processor_id <= amplifier_0_3_next_processor_id;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_next_config_id <= amplifier_0_1_next_config_id;
    end else begin
      amplifier_1_3_next_config_id <= amplifier_0_3_next_config_id;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 141:31]
      amplifier_1_3_is_valid_processor <= amplifier_0_1_is_valid_processor;
    end else begin
      amplifier_1_3_is_valid_processor <= amplifier_0_3_is_valid_processor;
    end
    if (first_proc_id == 2'h0) begin // @[ipsa.scala 126:38]
      next_proc_id_buf_0_0 <= 2'h0; // @[ipsa.scala 128:36]
    end else if (_amplifier_0_0_T) begin // @[ipsa.scala 113:38]
      next_proc_id_buf_0_0 <= 2'h0;
    end else begin
      next_proc_id_buf_0_0 <= trans_0_io_next_proc_id_out;
    end
    if (first_proc_id == 2'h1) begin // @[ipsa.scala 126:38]
      next_proc_id_buf_0_1 <= 2'h1; // @[ipsa.scala 128:36]
    end else if (_amplifier_0_1_T) begin // @[ipsa.scala 120:38]
      next_proc_id_buf_0_1 <= 2'h1;
    end else begin
      next_proc_id_buf_0_1 <= trans_1_io_next_proc_id_out;
    end
    if (first_proc_id == 2'h2) begin // @[ipsa.scala 126:38]
      next_proc_id_buf_0_2 <= 2'h2; // @[ipsa.scala 128:36]
    end else if (_amplifier_0_2_T) begin // @[ipsa.scala 113:38]
      next_proc_id_buf_0_2 <= 2'h2;
    end else begin
      next_proc_id_buf_0_2 <= trans_2_io_next_proc_id_out;
    end
    if (first_proc_id == 2'h3) begin // @[ipsa.scala 126:38]
      next_proc_id_buf_0_3 <= 2'h3; // @[ipsa.scala 128:36]
    end else if (_amplifier_0_3_T) begin // @[ipsa.scala 120:38]
      next_proc_id_buf_0_3 <= 2'h3;
    end else begin
      next_proc_id_buf_0_3 <= trans_3_io_next_proc_id_out;
    end
    if (_amplifier_1_0_T) begin // @[ipsa.scala 138:38]
      next_proc_id_buf_1_0 <= 2'h0;
    end else begin
      next_proc_id_buf_1_0 <= next_proc_id_buf_0_0;
    end
    if (_amplifier_1_1_T) begin // @[ipsa.scala 138:38]
      next_proc_id_buf_1_1 <= 2'h1;
    end else begin
      next_proc_id_buf_1_1 <= next_proc_id_buf_0_1;
    end
    if (_amplifier_1_2_T) begin // @[ipsa.scala 144:38]
      next_proc_id_buf_1_2 <= 2'h2;
    end else begin
      next_proc_id_buf_1_2 <= next_proc_id_buf_0_2;
    end
    if (_amplifier_1_3_T) begin // @[ipsa.scala 144:38]
      next_proc_id_buf_1_3 <= 2'h3;
    end else begin
      next_proc_id_buf_1_3 <= next_proc_id_buf_0_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  first_proc_id = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  last_proc_id = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  next_proc_id_0 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  next_proc_id_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  next_proc_id_2 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  next_proc_id_3 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  recv_0_data_0 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  recv_0_data_1 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  recv_0_data_2 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  recv_0_data_3 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  recv_0_data_4 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  recv_0_data_5 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  recv_0_data_6 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  recv_0_data_7 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  recv_0_data_8 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  recv_0_data_9 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  recv_0_data_10 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  recv_0_data_11 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  recv_0_data_12 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  recv_0_data_13 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  recv_0_data_14 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  recv_0_data_15 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  recv_0_data_16 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  recv_0_data_17 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  recv_0_data_18 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  recv_0_data_19 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  recv_0_data_20 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  recv_0_data_21 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  recv_0_data_22 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  recv_0_data_23 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  recv_0_data_24 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  recv_0_data_25 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  recv_0_data_26 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  recv_0_data_27 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  recv_0_data_28 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  recv_0_data_29 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  recv_0_data_30 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  recv_0_data_31 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  recv_0_data_32 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  recv_0_data_33 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  recv_0_data_34 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  recv_0_data_35 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  recv_0_data_36 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  recv_0_data_37 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  recv_0_data_38 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  recv_0_data_39 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  recv_0_data_40 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  recv_0_data_41 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  recv_0_data_42 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  recv_0_data_43 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  recv_0_data_44 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  recv_0_data_45 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  recv_0_data_46 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  recv_0_data_47 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  recv_0_data_48 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  recv_0_data_49 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  recv_0_data_50 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  recv_0_data_51 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  recv_0_data_52 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  recv_0_data_53 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  recv_0_data_54 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  recv_0_data_55 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  recv_0_data_56 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  recv_0_data_57 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  recv_0_data_58 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  recv_0_data_59 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  recv_0_data_60 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  recv_0_data_61 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  recv_0_data_62 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  recv_0_data_63 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  recv_0_data_64 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  recv_0_data_65 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  recv_0_data_66 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  recv_0_data_67 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  recv_0_data_68 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  recv_0_data_69 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  recv_0_data_70 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  recv_0_data_71 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  recv_0_data_72 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  recv_0_data_73 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  recv_0_data_74 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  recv_0_data_75 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  recv_0_data_76 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  recv_0_data_77 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  recv_0_data_78 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  recv_0_data_79 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  recv_0_data_80 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  recv_0_data_81 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  recv_0_data_82 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  recv_0_data_83 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  recv_0_data_84 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  recv_0_data_85 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  recv_0_data_86 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  recv_0_data_87 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  recv_0_data_88 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  recv_0_data_89 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  recv_0_data_90 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  recv_0_data_91 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  recv_0_data_92 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  recv_0_data_93 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  recv_0_data_94 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  recv_0_data_95 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  recv_0_data_96 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  recv_0_data_97 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  recv_0_data_98 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  recv_0_data_99 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  recv_0_data_100 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  recv_0_data_101 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  recv_0_data_102 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  recv_0_data_103 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  recv_0_data_104 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  recv_0_data_105 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  recv_0_data_106 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  recv_0_data_107 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  recv_0_data_108 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  recv_0_data_109 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  recv_0_data_110 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  recv_0_data_111 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  recv_0_data_112 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  recv_0_data_113 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  recv_0_data_114 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  recv_0_data_115 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  recv_0_data_116 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  recv_0_data_117 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  recv_0_data_118 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  recv_0_data_119 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  recv_0_data_120 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  recv_0_data_121 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  recv_0_data_122 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  recv_0_data_123 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  recv_0_data_124 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  recv_0_data_125 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  recv_0_data_126 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  recv_0_data_127 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  recv_0_data_128 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  recv_0_data_129 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  recv_0_data_130 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  recv_0_data_131 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  recv_0_data_132 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  recv_0_data_133 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  recv_0_data_134 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  recv_0_data_135 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  recv_0_data_136 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  recv_0_data_137 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  recv_0_data_138 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  recv_0_data_139 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  recv_0_data_140 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  recv_0_data_141 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  recv_0_data_142 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  recv_0_data_143 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  recv_0_data_144 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  recv_0_data_145 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  recv_0_data_146 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  recv_0_data_147 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  recv_0_data_148 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  recv_0_data_149 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  recv_0_data_150 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  recv_0_data_151 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  recv_0_data_152 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  recv_0_data_153 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  recv_0_data_154 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  recv_0_data_155 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  recv_0_data_156 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  recv_0_data_157 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  recv_0_data_158 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  recv_0_data_159 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  recv_0_data_160 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  recv_0_data_161 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  recv_0_data_162 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  recv_0_data_163 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  recv_0_data_164 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  recv_0_data_165 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  recv_0_data_166 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  recv_0_data_167 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  recv_0_data_168 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  recv_0_data_169 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  recv_0_data_170 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  recv_0_data_171 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  recv_0_data_172 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  recv_0_data_173 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  recv_0_data_174 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  recv_0_data_175 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  recv_0_data_176 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  recv_0_data_177 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  recv_0_data_178 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  recv_0_data_179 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  recv_0_data_180 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  recv_0_data_181 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  recv_0_data_182 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  recv_0_data_183 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  recv_0_data_184 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  recv_0_data_185 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  recv_0_data_186 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  recv_0_data_187 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  recv_0_data_188 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  recv_0_data_189 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  recv_0_data_190 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  recv_0_data_191 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  recv_0_data_192 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  recv_0_data_193 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  recv_0_data_194 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  recv_0_data_195 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  recv_0_data_196 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  recv_0_data_197 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  recv_0_data_198 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  recv_0_data_199 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  recv_0_data_200 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  recv_0_data_201 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  recv_0_data_202 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  recv_0_data_203 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  recv_0_data_204 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  recv_0_data_205 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  recv_0_data_206 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  recv_0_data_207 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  recv_0_data_208 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  recv_0_data_209 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  recv_0_data_210 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  recv_0_data_211 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  recv_0_data_212 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  recv_0_data_213 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  recv_0_data_214 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  recv_0_data_215 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  recv_0_data_216 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  recv_0_data_217 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  recv_0_data_218 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  recv_0_data_219 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  recv_0_data_220 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  recv_0_data_221 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  recv_0_data_222 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  recv_0_data_223 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  recv_0_data_224 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  recv_0_data_225 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  recv_0_data_226 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  recv_0_data_227 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  recv_0_data_228 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  recv_0_data_229 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  recv_0_data_230 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  recv_0_data_231 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  recv_0_data_232 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  recv_0_data_233 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  recv_0_data_234 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  recv_0_data_235 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  recv_0_data_236 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  recv_0_data_237 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  recv_0_data_238 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  recv_0_data_239 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  recv_0_data_240 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  recv_0_data_241 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  recv_0_data_242 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  recv_0_data_243 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  recv_0_data_244 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  recv_0_data_245 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  recv_0_data_246 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  recv_0_data_247 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  recv_0_data_248 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  recv_0_data_249 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  recv_0_data_250 = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  recv_0_data_251 = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  recv_0_data_252 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  recv_0_data_253 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  recv_0_data_254 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  recv_0_data_255 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  recv_0_header_0 = _RAND_262[15:0];
  _RAND_263 = {1{`RANDOM}};
  recv_0_header_1 = _RAND_263[15:0];
  _RAND_264 = {1{`RANDOM}};
  recv_0_header_2 = _RAND_264[15:0];
  _RAND_265 = {1{`RANDOM}};
  recv_0_header_3 = _RAND_265[15:0];
  _RAND_266 = {1{`RANDOM}};
  recv_0_header_4 = _RAND_266[15:0];
  _RAND_267 = {1{`RANDOM}};
  recv_0_header_5 = _RAND_267[15:0];
  _RAND_268 = {1{`RANDOM}};
  recv_0_header_6 = _RAND_268[15:0];
  _RAND_269 = {1{`RANDOM}};
  recv_0_header_7 = _RAND_269[15:0];
  _RAND_270 = {1{`RANDOM}};
  recv_0_header_8 = _RAND_270[15:0];
  _RAND_271 = {1{`RANDOM}};
  recv_0_header_9 = _RAND_271[15:0];
  _RAND_272 = {1{`RANDOM}};
  recv_0_header_10 = _RAND_272[15:0];
  _RAND_273 = {1{`RANDOM}};
  recv_0_header_11 = _RAND_273[15:0];
  _RAND_274 = {1{`RANDOM}};
  recv_0_header_12 = _RAND_274[15:0];
  _RAND_275 = {1{`RANDOM}};
  recv_0_header_13 = _RAND_275[15:0];
  _RAND_276 = {1{`RANDOM}};
  recv_0_header_14 = _RAND_276[15:0];
  _RAND_277 = {1{`RANDOM}};
  recv_0_header_15 = _RAND_277[15:0];
  _RAND_278 = {1{`RANDOM}};
  recv_0_parse_current_state = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  recv_0_parse_current_offset = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  recv_0_parse_transition_field = _RAND_280[15:0];
  _RAND_281 = {1{`RANDOM}};
  recv_0_next_processor_id = _RAND_281[1:0];
  _RAND_282 = {1{`RANDOM}};
  recv_0_next_config_id = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  recv_0_is_valid_processor = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  recv_1_data_0 = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  recv_1_data_1 = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  recv_1_data_2 = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  recv_1_data_3 = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  recv_1_data_4 = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  recv_1_data_5 = _RAND_289[7:0];
  _RAND_290 = {1{`RANDOM}};
  recv_1_data_6 = _RAND_290[7:0];
  _RAND_291 = {1{`RANDOM}};
  recv_1_data_7 = _RAND_291[7:0];
  _RAND_292 = {1{`RANDOM}};
  recv_1_data_8 = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  recv_1_data_9 = _RAND_293[7:0];
  _RAND_294 = {1{`RANDOM}};
  recv_1_data_10 = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  recv_1_data_11 = _RAND_295[7:0];
  _RAND_296 = {1{`RANDOM}};
  recv_1_data_12 = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  recv_1_data_13 = _RAND_297[7:0];
  _RAND_298 = {1{`RANDOM}};
  recv_1_data_14 = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  recv_1_data_15 = _RAND_299[7:0];
  _RAND_300 = {1{`RANDOM}};
  recv_1_data_16 = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  recv_1_data_17 = _RAND_301[7:0];
  _RAND_302 = {1{`RANDOM}};
  recv_1_data_18 = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  recv_1_data_19 = _RAND_303[7:0];
  _RAND_304 = {1{`RANDOM}};
  recv_1_data_20 = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  recv_1_data_21 = _RAND_305[7:0];
  _RAND_306 = {1{`RANDOM}};
  recv_1_data_22 = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  recv_1_data_23 = _RAND_307[7:0];
  _RAND_308 = {1{`RANDOM}};
  recv_1_data_24 = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  recv_1_data_25 = _RAND_309[7:0];
  _RAND_310 = {1{`RANDOM}};
  recv_1_data_26 = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  recv_1_data_27 = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  recv_1_data_28 = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  recv_1_data_29 = _RAND_313[7:0];
  _RAND_314 = {1{`RANDOM}};
  recv_1_data_30 = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  recv_1_data_31 = _RAND_315[7:0];
  _RAND_316 = {1{`RANDOM}};
  recv_1_data_32 = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  recv_1_data_33 = _RAND_317[7:0];
  _RAND_318 = {1{`RANDOM}};
  recv_1_data_34 = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  recv_1_data_35 = _RAND_319[7:0];
  _RAND_320 = {1{`RANDOM}};
  recv_1_data_36 = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  recv_1_data_37 = _RAND_321[7:0];
  _RAND_322 = {1{`RANDOM}};
  recv_1_data_38 = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  recv_1_data_39 = _RAND_323[7:0];
  _RAND_324 = {1{`RANDOM}};
  recv_1_data_40 = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  recv_1_data_41 = _RAND_325[7:0];
  _RAND_326 = {1{`RANDOM}};
  recv_1_data_42 = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  recv_1_data_43 = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  recv_1_data_44 = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  recv_1_data_45 = _RAND_329[7:0];
  _RAND_330 = {1{`RANDOM}};
  recv_1_data_46 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  recv_1_data_47 = _RAND_331[7:0];
  _RAND_332 = {1{`RANDOM}};
  recv_1_data_48 = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  recv_1_data_49 = _RAND_333[7:0];
  _RAND_334 = {1{`RANDOM}};
  recv_1_data_50 = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  recv_1_data_51 = _RAND_335[7:0];
  _RAND_336 = {1{`RANDOM}};
  recv_1_data_52 = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  recv_1_data_53 = _RAND_337[7:0];
  _RAND_338 = {1{`RANDOM}};
  recv_1_data_54 = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  recv_1_data_55 = _RAND_339[7:0];
  _RAND_340 = {1{`RANDOM}};
  recv_1_data_56 = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  recv_1_data_57 = _RAND_341[7:0];
  _RAND_342 = {1{`RANDOM}};
  recv_1_data_58 = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  recv_1_data_59 = _RAND_343[7:0];
  _RAND_344 = {1{`RANDOM}};
  recv_1_data_60 = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  recv_1_data_61 = _RAND_345[7:0];
  _RAND_346 = {1{`RANDOM}};
  recv_1_data_62 = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  recv_1_data_63 = _RAND_347[7:0];
  _RAND_348 = {1{`RANDOM}};
  recv_1_data_64 = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  recv_1_data_65 = _RAND_349[7:0];
  _RAND_350 = {1{`RANDOM}};
  recv_1_data_66 = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  recv_1_data_67 = _RAND_351[7:0];
  _RAND_352 = {1{`RANDOM}};
  recv_1_data_68 = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  recv_1_data_69 = _RAND_353[7:0];
  _RAND_354 = {1{`RANDOM}};
  recv_1_data_70 = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  recv_1_data_71 = _RAND_355[7:0];
  _RAND_356 = {1{`RANDOM}};
  recv_1_data_72 = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  recv_1_data_73 = _RAND_357[7:0];
  _RAND_358 = {1{`RANDOM}};
  recv_1_data_74 = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  recv_1_data_75 = _RAND_359[7:0];
  _RAND_360 = {1{`RANDOM}};
  recv_1_data_76 = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  recv_1_data_77 = _RAND_361[7:0];
  _RAND_362 = {1{`RANDOM}};
  recv_1_data_78 = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  recv_1_data_79 = _RAND_363[7:0];
  _RAND_364 = {1{`RANDOM}};
  recv_1_data_80 = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  recv_1_data_81 = _RAND_365[7:0];
  _RAND_366 = {1{`RANDOM}};
  recv_1_data_82 = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  recv_1_data_83 = _RAND_367[7:0];
  _RAND_368 = {1{`RANDOM}};
  recv_1_data_84 = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  recv_1_data_85 = _RAND_369[7:0];
  _RAND_370 = {1{`RANDOM}};
  recv_1_data_86 = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  recv_1_data_87 = _RAND_371[7:0];
  _RAND_372 = {1{`RANDOM}};
  recv_1_data_88 = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  recv_1_data_89 = _RAND_373[7:0];
  _RAND_374 = {1{`RANDOM}};
  recv_1_data_90 = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  recv_1_data_91 = _RAND_375[7:0];
  _RAND_376 = {1{`RANDOM}};
  recv_1_data_92 = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  recv_1_data_93 = _RAND_377[7:0];
  _RAND_378 = {1{`RANDOM}};
  recv_1_data_94 = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  recv_1_data_95 = _RAND_379[7:0];
  _RAND_380 = {1{`RANDOM}};
  recv_1_data_96 = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  recv_1_data_97 = _RAND_381[7:0];
  _RAND_382 = {1{`RANDOM}};
  recv_1_data_98 = _RAND_382[7:0];
  _RAND_383 = {1{`RANDOM}};
  recv_1_data_99 = _RAND_383[7:0];
  _RAND_384 = {1{`RANDOM}};
  recv_1_data_100 = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  recv_1_data_101 = _RAND_385[7:0];
  _RAND_386 = {1{`RANDOM}};
  recv_1_data_102 = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  recv_1_data_103 = _RAND_387[7:0];
  _RAND_388 = {1{`RANDOM}};
  recv_1_data_104 = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  recv_1_data_105 = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  recv_1_data_106 = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  recv_1_data_107 = _RAND_391[7:0];
  _RAND_392 = {1{`RANDOM}};
  recv_1_data_108 = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  recv_1_data_109 = _RAND_393[7:0];
  _RAND_394 = {1{`RANDOM}};
  recv_1_data_110 = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  recv_1_data_111 = _RAND_395[7:0];
  _RAND_396 = {1{`RANDOM}};
  recv_1_data_112 = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  recv_1_data_113 = _RAND_397[7:0];
  _RAND_398 = {1{`RANDOM}};
  recv_1_data_114 = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  recv_1_data_115 = _RAND_399[7:0];
  _RAND_400 = {1{`RANDOM}};
  recv_1_data_116 = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  recv_1_data_117 = _RAND_401[7:0];
  _RAND_402 = {1{`RANDOM}};
  recv_1_data_118 = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  recv_1_data_119 = _RAND_403[7:0];
  _RAND_404 = {1{`RANDOM}};
  recv_1_data_120 = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  recv_1_data_121 = _RAND_405[7:0];
  _RAND_406 = {1{`RANDOM}};
  recv_1_data_122 = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  recv_1_data_123 = _RAND_407[7:0];
  _RAND_408 = {1{`RANDOM}};
  recv_1_data_124 = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  recv_1_data_125 = _RAND_409[7:0];
  _RAND_410 = {1{`RANDOM}};
  recv_1_data_126 = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  recv_1_data_127 = _RAND_411[7:0];
  _RAND_412 = {1{`RANDOM}};
  recv_1_data_128 = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  recv_1_data_129 = _RAND_413[7:0];
  _RAND_414 = {1{`RANDOM}};
  recv_1_data_130 = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  recv_1_data_131 = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  recv_1_data_132 = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  recv_1_data_133 = _RAND_417[7:0];
  _RAND_418 = {1{`RANDOM}};
  recv_1_data_134 = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  recv_1_data_135 = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  recv_1_data_136 = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  recv_1_data_137 = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  recv_1_data_138 = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  recv_1_data_139 = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  recv_1_data_140 = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  recv_1_data_141 = _RAND_425[7:0];
  _RAND_426 = {1{`RANDOM}};
  recv_1_data_142 = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  recv_1_data_143 = _RAND_427[7:0];
  _RAND_428 = {1{`RANDOM}};
  recv_1_data_144 = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  recv_1_data_145 = _RAND_429[7:0];
  _RAND_430 = {1{`RANDOM}};
  recv_1_data_146 = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  recv_1_data_147 = _RAND_431[7:0];
  _RAND_432 = {1{`RANDOM}};
  recv_1_data_148 = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  recv_1_data_149 = _RAND_433[7:0];
  _RAND_434 = {1{`RANDOM}};
  recv_1_data_150 = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  recv_1_data_151 = _RAND_435[7:0];
  _RAND_436 = {1{`RANDOM}};
  recv_1_data_152 = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  recv_1_data_153 = _RAND_437[7:0];
  _RAND_438 = {1{`RANDOM}};
  recv_1_data_154 = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  recv_1_data_155 = _RAND_439[7:0];
  _RAND_440 = {1{`RANDOM}};
  recv_1_data_156 = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  recv_1_data_157 = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  recv_1_data_158 = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  recv_1_data_159 = _RAND_443[7:0];
  _RAND_444 = {1{`RANDOM}};
  recv_1_data_160 = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  recv_1_data_161 = _RAND_445[7:0];
  _RAND_446 = {1{`RANDOM}};
  recv_1_data_162 = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  recv_1_data_163 = _RAND_447[7:0];
  _RAND_448 = {1{`RANDOM}};
  recv_1_data_164 = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  recv_1_data_165 = _RAND_449[7:0];
  _RAND_450 = {1{`RANDOM}};
  recv_1_data_166 = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  recv_1_data_167 = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  recv_1_data_168 = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  recv_1_data_169 = _RAND_453[7:0];
  _RAND_454 = {1{`RANDOM}};
  recv_1_data_170 = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  recv_1_data_171 = _RAND_455[7:0];
  _RAND_456 = {1{`RANDOM}};
  recv_1_data_172 = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  recv_1_data_173 = _RAND_457[7:0];
  _RAND_458 = {1{`RANDOM}};
  recv_1_data_174 = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  recv_1_data_175 = _RAND_459[7:0];
  _RAND_460 = {1{`RANDOM}};
  recv_1_data_176 = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  recv_1_data_177 = _RAND_461[7:0];
  _RAND_462 = {1{`RANDOM}};
  recv_1_data_178 = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  recv_1_data_179 = _RAND_463[7:0];
  _RAND_464 = {1{`RANDOM}};
  recv_1_data_180 = _RAND_464[7:0];
  _RAND_465 = {1{`RANDOM}};
  recv_1_data_181 = _RAND_465[7:0];
  _RAND_466 = {1{`RANDOM}};
  recv_1_data_182 = _RAND_466[7:0];
  _RAND_467 = {1{`RANDOM}};
  recv_1_data_183 = _RAND_467[7:0];
  _RAND_468 = {1{`RANDOM}};
  recv_1_data_184 = _RAND_468[7:0];
  _RAND_469 = {1{`RANDOM}};
  recv_1_data_185 = _RAND_469[7:0];
  _RAND_470 = {1{`RANDOM}};
  recv_1_data_186 = _RAND_470[7:0];
  _RAND_471 = {1{`RANDOM}};
  recv_1_data_187 = _RAND_471[7:0];
  _RAND_472 = {1{`RANDOM}};
  recv_1_data_188 = _RAND_472[7:0];
  _RAND_473 = {1{`RANDOM}};
  recv_1_data_189 = _RAND_473[7:0];
  _RAND_474 = {1{`RANDOM}};
  recv_1_data_190 = _RAND_474[7:0];
  _RAND_475 = {1{`RANDOM}};
  recv_1_data_191 = _RAND_475[7:0];
  _RAND_476 = {1{`RANDOM}};
  recv_1_data_192 = _RAND_476[7:0];
  _RAND_477 = {1{`RANDOM}};
  recv_1_data_193 = _RAND_477[7:0];
  _RAND_478 = {1{`RANDOM}};
  recv_1_data_194 = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  recv_1_data_195 = _RAND_479[7:0];
  _RAND_480 = {1{`RANDOM}};
  recv_1_data_196 = _RAND_480[7:0];
  _RAND_481 = {1{`RANDOM}};
  recv_1_data_197 = _RAND_481[7:0];
  _RAND_482 = {1{`RANDOM}};
  recv_1_data_198 = _RAND_482[7:0];
  _RAND_483 = {1{`RANDOM}};
  recv_1_data_199 = _RAND_483[7:0];
  _RAND_484 = {1{`RANDOM}};
  recv_1_data_200 = _RAND_484[7:0];
  _RAND_485 = {1{`RANDOM}};
  recv_1_data_201 = _RAND_485[7:0];
  _RAND_486 = {1{`RANDOM}};
  recv_1_data_202 = _RAND_486[7:0];
  _RAND_487 = {1{`RANDOM}};
  recv_1_data_203 = _RAND_487[7:0];
  _RAND_488 = {1{`RANDOM}};
  recv_1_data_204 = _RAND_488[7:0];
  _RAND_489 = {1{`RANDOM}};
  recv_1_data_205 = _RAND_489[7:0];
  _RAND_490 = {1{`RANDOM}};
  recv_1_data_206 = _RAND_490[7:0];
  _RAND_491 = {1{`RANDOM}};
  recv_1_data_207 = _RAND_491[7:0];
  _RAND_492 = {1{`RANDOM}};
  recv_1_data_208 = _RAND_492[7:0];
  _RAND_493 = {1{`RANDOM}};
  recv_1_data_209 = _RAND_493[7:0];
  _RAND_494 = {1{`RANDOM}};
  recv_1_data_210 = _RAND_494[7:0];
  _RAND_495 = {1{`RANDOM}};
  recv_1_data_211 = _RAND_495[7:0];
  _RAND_496 = {1{`RANDOM}};
  recv_1_data_212 = _RAND_496[7:0];
  _RAND_497 = {1{`RANDOM}};
  recv_1_data_213 = _RAND_497[7:0];
  _RAND_498 = {1{`RANDOM}};
  recv_1_data_214 = _RAND_498[7:0];
  _RAND_499 = {1{`RANDOM}};
  recv_1_data_215 = _RAND_499[7:0];
  _RAND_500 = {1{`RANDOM}};
  recv_1_data_216 = _RAND_500[7:0];
  _RAND_501 = {1{`RANDOM}};
  recv_1_data_217 = _RAND_501[7:0];
  _RAND_502 = {1{`RANDOM}};
  recv_1_data_218 = _RAND_502[7:0];
  _RAND_503 = {1{`RANDOM}};
  recv_1_data_219 = _RAND_503[7:0];
  _RAND_504 = {1{`RANDOM}};
  recv_1_data_220 = _RAND_504[7:0];
  _RAND_505 = {1{`RANDOM}};
  recv_1_data_221 = _RAND_505[7:0];
  _RAND_506 = {1{`RANDOM}};
  recv_1_data_222 = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  recv_1_data_223 = _RAND_507[7:0];
  _RAND_508 = {1{`RANDOM}};
  recv_1_data_224 = _RAND_508[7:0];
  _RAND_509 = {1{`RANDOM}};
  recv_1_data_225 = _RAND_509[7:0];
  _RAND_510 = {1{`RANDOM}};
  recv_1_data_226 = _RAND_510[7:0];
  _RAND_511 = {1{`RANDOM}};
  recv_1_data_227 = _RAND_511[7:0];
  _RAND_512 = {1{`RANDOM}};
  recv_1_data_228 = _RAND_512[7:0];
  _RAND_513 = {1{`RANDOM}};
  recv_1_data_229 = _RAND_513[7:0];
  _RAND_514 = {1{`RANDOM}};
  recv_1_data_230 = _RAND_514[7:0];
  _RAND_515 = {1{`RANDOM}};
  recv_1_data_231 = _RAND_515[7:0];
  _RAND_516 = {1{`RANDOM}};
  recv_1_data_232 = _RAND_516[7:0];
  _RAND_517 = {1{`RANDOM}};
  recv_1_data_233 = _RAND_517[7:0];
  _RAND_518 = {1{`RANDOM}};
  recv_1_data_234 = _RAND_518[7:0];
  _RAND_519 = {1{`RANDOM}};
  recv_1_data_235 = _RAND_519[7:0];
  _RAND_520 = {1{`RANDOM}};
  recv_1_data_236 = _RAND_520[7:0];
  _RAND_521 = {1{`RANDOM}};
  recv_1_data_237 = _RAND_521[7:0];
  _RAND_522 = {1{`RANDOM}};
  recv_1_data_238 = _RAND_522[7:0];
  _RAND_523 = {1{`RANDOM}};
  recv_1_data_239 = _RAND_523[7:0];
  _RAND_524 = {1{`RANDOM}};
  recv_1_data_240 = _RAND_524[7:0];
  _RAND_525 = {1{`RANDOM}};
  recv_1_data_241 = _RAND_525[7:0];
  _RAND_526 = {1{`RANDOM}};
  recv_1_data_242 = _RAND_526[7:0];
  _RAND_527 = {1{`RANDOM}};
  recv_1_data_243 = _RAND_527[7:0];
  _RAND_528 = {1{`RANDOM}};
  recv_1_data_244 = _RAND_528[7:0];
  _RAND_529 = {1{`RANDOM}};
  recv_1_data_245 = _RAND_529[7:0];
  _RAND_530 = {1{`RANDOM}};
  recv_1_data_246 = _RAND_530[7:0];
  _RAND_531 = {1{`RANDOM}};
  recv_1_data_247 = _RAND_531[7:0];
  _RAND_532 = {1{`RANDOM}};
  recv_1_data_248 = _RAND_532[7:0];
  _RAND_533 = {1{`RANDOM}};
  recv_1_data_249 = _RAND_533[7:0];
  _RAND_534 = {1{`RANDOM}};
  recv_1_data_250 = _RAND_534[7:0];
  _RAND_535 = {1{`RANDOM}};
  recv_1_data_251 = _RAND_535[7:0];
  _RAND_536 = {1{`RANDOM}};
  recv_1_data_252 = _RAND_536[7:0];
  _RAND_537 = {1{`RANDOM}};
  recv_1_data_253 = _RAND_537[7:0];
  _RAND_538 = {1{`RANDOM}};
  recv_1_data_254 = _RAND_538[7:0];
  _RAND_539 = {1{`RANDOM}};
  recv_1_data_255 = _RAND_539[7:0];
  _RAND_540 = {1{`RANDOM}};
  recv_1_header_0 = _RAND_540[15:0];
  _RAND_541 = {1{`RANDOM}};
  recv_1_header_1 = _RAND_541[15:0];
  _RAND_542 = {1{`RANDOM}};
  recv_1_header_2 = _RAND_542[15:0];
  _RAND_543 = {1{`RANDOM}};
  recv_1_header_3 = _RAND_543[15:0];
  _RAND_544 = {1{`RANDOM}};
  recv_1_header_4 = _RAND_544[15:0];
  _RAND_545 = {1{`RANDOM}};
  recv_1_header_5 = _RAND_545[15:0];
  _RAND_546 = {1{`RANDOM}};
  recv_1_header_6 = _RAND_546[15:0];
  _RAND_547 = {1{`RANDOM}};
  recv_1_header_7 = _RAND_547[15:0];
  _RAND_548 = {1{`RANDOM}};
  recv_1_header_8 = _RAND_548[15:0];
  _RAND_549 = {1{`RANDOM}};
  recv_1_header_9 = _RAND_549[15:0];
  _RAND_550 = {1{`RANDOM}};
  recv_1_header_10 = _RAND_550[15:0];
  _RAND_551 = {1{`RANDOM}};
  recv_1_header_11 = _RAND_551[15:0];
  _RAND_552 = {1{`RANDOM}};
  recv_1_header_12 = _RAND_552[15:0];
  _RAND_553 = {1{`RANDOM}};
  recv_1_header_13 = _RAND_553[15:0];
  _RAND_554 = {1{`RANDOM}};
  recv_1_header_14 = _RAND_554[15:0];
  _RAND_555 = {1{`RANDOM}};
  recv_1_header_15 = _RAND_555[15:0];
  _RAND_556 = {1{`RANDOM}};
  recv_1_parse_current_state = _RAND_556[7:0];
  _RAND_557 = {1{`RANDOM}};
  recv_1_parse_current_offset = _RAND_557[7:0];
  _RAND_558 = {1{`RANDOM}};
  recv_1_parse_transition_field = _RAND_558[15:0];
  _RAND_559 = {1{`RANDOM}};
  recv_1_next_processor_id = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  recv_1_next_config_id = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  recv_1_is_valid_processor = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  recv_2_data_0 = _RAND_562[7:0];
  _RAND_563 = {1{`RANDOM}};
  recv_2_data_1 = _RAND_563[7:0];
  _RAND_564 = {1{`RANDOM}};
  recv_2_data_2 = _RAND_564[7:0];
  _RAND_565 = {1{`RANDOM}};
  recv_2_data_3 = _RAND_565[7:0];
  _RAND_566 = {1{`RANDOM}};
  recv_2_data_4 = _RAND_566[7:0];
  _RAND_567 = {1{`RANDOM}};
  recv_2_data_5 = _RAND_567[7:0];
  _RAND_568 = {1{`RANDOM}};
  recv_2_data_6 = _RAND_568[7:0];
  _RAND_569 = {1{`RANDOM}};
  recv_2_data_7 = _RAND_569[7:0];
  _RAND_570 = {1{`RANDOM}};
  recv_2_data_8 = _RAND_570[7:0];
  _RAND_571 = {1{`RANDOM}};
  recv_2_data_9 = _RAND_571[7:0];
  _RAND_572 = {1{`RANDOM}};
  recv_2_data_10 = _RAND_572[7:0];
  _RAND_573 = {1{`RANDOM}};
  recv_2_data_11 = _RAND_573[7:0];
  _RAND_574 = {1{`RANDOM}};
  recv_2_data_12 = _RAND_574[7:0];
  _RAND_575 = {1{`RANDOM}};
  recv_2_data_13 = _RAND_575[7:0];
  _RAND_576 = {1{`RANDOM}};
  recv_2_data_14 = _RAND_576[7:0];
  _RAND_577 = {1{`RANDOM}};
  recv_2_data_15 = _RAND_577[7:0];
  _RAND_578 = {1{`RANDOM}};
  recv_2_data_16 = _RAND_578[7:0];
  _RAND_579 = {1{`RANDOM}};
  recv_2_data_17 = _RAND_579[7:0];
  _RAND_580 = {1{`RANDOM}};
  recv_2_data_18 = _RAND_580[7:0];
  _RAND_581 = {1{`RANDOM}};
  recv_2_data_19 = _RAND_581[7:0];
  _RAND_582 = {1{`RANDOM}};
  recv_2_data_20 = _RAND_582[7:0];
  _RAND_583 = {1{`RANDOM}};
  recv_2_data_21 = _RAND_583[7:0];
  _RAND_584 = {1{`RANDOM}};
  recv_2_data_22 = _RAND_584[7:0];
  _RAND_585 = {1{`RANDOM}};
  recv_2_data_23 = _RAND_585[7:0];
  _RAND_586 = {1{`RANDOM}};
  recv_2_data_24 = _RAND_586[7:0];
  _RAND_587 = {1{`RANDOM}};
  recv_2_data_25 = _RAND_587[7:0];
  _RAND_588 = {1{`RANDOM}};
  recv_2_data_26 = _RAND_588[7:0];
  _RAND_589 = {1{`RANDOM}};
  recv_2_data_27 = _RAND_589[7:0];
  _RAND_590 = {1{`RANDOM}};
  recv_2_data_28 = _RAND_590[7:0];
  _RAND_591 = {1{`RANDOM}};
  recv_2_data_29 = _RAND_591[7:0];
  _RAND_592 = {1{`RANDOM}};
  recv_2_data_30 = _RAND_592[7:0];
  _RAND_593 = {1{`RANDOM}};
  recv_2_data_31 = _RAND_593[7:0];
  _RAND_594 = {1{`RANDOM}};
  recv_2_data_32 = _RAND_594[7:0];
  _RAND_595 = {1{`RANDOM}};
  recv_2_data_33 = _RAND_595[7:0];
  _RAND_596 = {1{`RANDOM}};
  recv_2_data_34 = _RAND_596[7:0];
  _RAND_597 = {1{`RANDOM}};
  recv_2_data_35 = _RAND_597[7:0];
  _RAND_598 = {1{`RANDOM}};
  recv_2_data_36 = _RAND_598[7:0];
  _RAND_599 = {1{`RANDOM}};
  recv_2_data_37 = _RAND_599[7:0];
  _RAND_600 = {1{`RANDOM}};
  recv_2_data_38 = _RAND_600[7:0];
  _RAND_601 = {1{`RANDOM}};
  recv_2_data_39 = _RAND_601[7:0];
  _RAND_602 = {1{`RANDOM}};
  recv_2_data_40 = _RAND_602[7:0];
  _RAND_603 = {1{`RANDOM}};
  recv_2_data_41 = _RAND_603[7:0];
  _RAND_604 = {1{`RANDOM}};
  recv_2_data_42 = _RAND_604[7:0];
  _RAND_605 = {1{`RANDOM}};
  recv_2_data_43 = _RAND_605[7:0];
  _RAND_606 = {1{`RANDOM}};
  recv_2_data_44 = _RAND_606[7:0];
  _RAND_607 = {1{`RANDOM}};
  recv_2_data_45 = _RAND_607[7:0];
  _RAND_608 = {1{`RANDOM}};
  recv_2_data_46 = _RAND_608[7:0];
  _RAND_609 = {1{`RANDOM}};
  recv_2_data_47 = _RAND_609[7:0];
  _RAND_610 = {1{`RANDOM}};
  recv_2_data_48 = _RAND_610[7:0];
  _RAND_611 = {1{`RANDOM}};
  recv_2_data_49 = _RAND_611[7:0];
  _RAND_612 = {1{`RANDOM}};
  recv_2_data_50 = _RAND_612[7:0];
  _RAND_613 = {1{`RANDOM}};
  recv_2_data_51 = _RAND_613[7:0];
  _RAND_614 = {1{`RANDOM}};
  recv_2_data_52 = _RAND_614[7:0];
  _RAND_615 = {1{`RANDOM}};
  recv_2_data_53 = _RAND_615[7:0];
  _RAND_616 = {1{`RANDOM}};
  recv_2_data_54 = _RAND_616[7:0];
  _RAND_617 = {1{`RANDOM}};
  recv_2_data_55 = _RAND_617[7:0];
  _RAND_618 = {1{`RANDOM}};
  recv_2_data_56 = _RAND_618[7:0];
  _RAND_619 = {1{`RANDOM}};
  recv_2_data_57 = _RAND_619[7:0];
  _RAND_620 = {1{`RANDOM}};
  recv_2_data_58 = _RAND_620[7:0];
  _RAND_621 = {1{`RANDOM}};
  recv_2_data_59 = _RAND_621[7:0];
  _RAND_622 = {1{`RANDOM}};
  recv_2_data_60 = _RAND_622[7:0];
  _RAND_623 = {1{`RANDOM}};
  recv_2_data_61 = _RAND_623[7:0];
  _RAND_624 = {1{`RANDOM}};
  recv_2_data_62 = _RAND_624[7:0];
  _RAND_625 = {1{`RANDOM}};
  recv_2_data_63 = _RAND_625[7:0];
  _RAND_626 = {1{`RANDOM}};
  recv_2_data_64 = _RAND_626[7:0];
  _RAND_627 = {1{`RANDOM}};
  recv_2_data_65 = _RAND_627[7:0];
  _RAND_628 = {1{`RANDOM}};
  recv_2_data_66 = _RAND_628[7:0];
  _RAND_629 = {1{`RANDOM}};
  recv_2_data_67 = _RAND_629[7:0];
  _RAND_630 = {1{`RANDOM}};
  recv_2_data_68 = _RAND_630[7:0];
  _RAND_631 = {1{`RANDOM}};
  recv_2_data_69 = _RAND_631[7:0];
  _RAND_632 = {1{`RANDOM}};
  recv_2_data_70 = _RAND_632[7:0];
  _RAND_633 = {1{`RANDOM}};
  recv_2_data_71 = _RAND_633[7:0];
  _RAND_634 = {1{`RANDOM}};
  recv_2_data_72 = _RAND_634[7:0];
  _RAND_635 = {1{`RANDOM}};
  recv_2_data_73 = _RAND_635[7:0];
  _RAND_636 = {1{`RANDOM}};
  recv_2_data_74 = _RAND_636[7:0];
  _RAND_637 = {1{`RANDOM}};
  recv_2_data_75 = _RAND_637[7:0];
  _RAND_638 = {1{`RANDOM}};
  recv_2_data_76 = _RAND_638[7:0];
  _RAND_639 = {1{`RANDOM}};
  recv_2_data_77 = _RAND_639[7:0];
  _RAND_640 = {1{`RANDOM}};
  recv_2_data_78 = _RAND_640[7:0];
  _RAND_641 = {1{`RANDOM}};
  recv_2_data_79 = _RAND_641[7:0];
  _RAND_642 = {1{`RANDOM}};
  recv_2_data_80 = _RAND_642[7:0];
  _RAND_643 = {1{`RANDOM}};
  recv_2_data_81 = _RAND_643[7:0];
  _RAND_644 = {1{`RANDOM}};
  recv_2_data_82 = _RAND_644[7:0];
  _RAND_645 = {1{`RANDOM}};
  recv_2_data_83 = _RAND_645[7:0];
  _RAND_646 = {1{`RANDOM}};
  recv_2_data_84 = _RAND_646[7:0];
  _RAND_647 = {1{`RANDOM}};
  recv_2_data_85 = _RAND_647[7:0];
  _RAND_648 = {1{`RANDOM}};
  recv_2_data_86 = _RAND_648[7:0];
  _RAND_649 = {1{`RANDOM}};
  recv_2_data_87 = _RAND_649[7:0];
  _RAND_650 = {1{`RANDOM}};
  recv_2_data_88 = _RAND_650[7:0];
  _RAND_651 = {1{`RANDOM}};
  recv_2_data_89 = _RAND_651[7:0];
  _RAND_652 = {1{`RANDOM}};
  recv_2_data_90 = _RAND_652[7:0];
  _RAND_653 = {1{`RANDOM}};
  recv_2_data_91 = _RAND_653[7:0];
  _RAND_654 = {1{`RANDOM}};
  recv_2_data_92 = _RAND_654[7:0];
  _RAND_655 = {1{`RANDOM}};
  recv_2_data_93 = _RAND_655[7:0];
  _RAND_656 = {1{`RANDOM}};
  recv_2_data_94 = _RAND_656[7:0];
  _RAND_657 = {1{`RANDOM}};
  recv_2_data_95 = _RAND_657[7:0];
  _RAND_658 = {1{`RANDOM}};
  recv_2_data_96 = _RAND_658[7:0];
  _RAND_659 = {1{`RANDOM}};
  recv_2_data_97 = _RAND_659[7:0];
  _RAND_660 = {1{`RANDOM}};
  recv_2_data_98 = _RAND_660[7:0];
  _RAND_661 = {1{`RANDOM}};
  recv_2_data_99 = _RAND_661[7:0];
  _RAND_662 = {1{`RANDOM}};
  recv_2_data_100 = _RAND_662[7:0];
  _RAND_663 = {1{`RANDOM}};
  recv_2_data_101 = _RAND_663[7:0];
  _RAND_664 = {1{`RANDOM}};
  recv_2_data_102 = _RAND_664[7:0];
  _RAND_665 = {1{`RANDOM}};
  recv_2_data_103 = _RAND_665[7:0];
  _RAND_666 = {1{`RANDOM}};
  recv_2_data_104 = _RAND_666[7:0];
  _RAND_667 = {1{`RANDOM}};
  recv_2_data_105 = _RAND_667[7:0];
  _RAND_668 = {1{`RANDOM}};
  recv_2_data_106 = _RAND_668[7:0];
  _RAND_669 = {1{`RANDOM}};
  recv_2_data_107 = _RAND_669[7:0];
  _RAND_670 = {1{`RANDOM}};
  recv_2_data_108 = _RAND_670[7:0];
  _RAND_671 = {1{`RANDOM}};
  recv_2_data_109 = _RAND_671[7:0];
  _RAND_672 = {1{`RANDOM}};
  recv_2_data_110 = _RAND_672[7:0];
  _RAND_673 = {1{`RANDOM}};
  recv_2_data_111 = _RAND_673[7:0];
  _RAND_674 = {1{`RANDOM}};
  recv_2_data_112 = _RAND_674[7:0];
  _RAND_675 = {1{`RANDOM}};
  recv_2_data_113 = _RAND_675[7:0];
  _RAND_676 = {1{`RANDOM}};
  recv_2_data_114 = _RAND_676[7:0];
  _RAND_677 = {1{`RANDOM}};
  recv_2_data_115 = _RAND_677[7:0];
  _RAND_678 = {1{`RANDOM}};
  recv_2_data_116 = _RAND_678[7:0];
  _RAND_679 = {1{`RANDOM}};
  recv_2_data_117 = _RAND_679[7:0];
  _RAND_680 = {1{`RANDOM}};
  recv_2_data_118 = _RAND_680[7:0];
  _RAND_681 = {1{`RANDOM}};
  recv_2_data_119 = _RAND_681[7:0];
  _RAND_682 = {1{`RANDOM}};
  recv_2_data_120 = _RAND_682[7:0];
  _RAND_683 = {1{`RANDOM}};
  recv_2_data_121 = _RAND_683[7:0];
  _RAND_684 = {1{`RANDOM}};
  recv_2_data_122 = _RAND_684[7:0];
  _RAND_685 = {1{`RANDOM}};
  recv_2_data_123 = _RAND_685[7:0];
  _RAND_686 = {1{`RANDOM}};
  recv_2_data_124 = _RAND_686[7:0];
  _RAND_687 = {1{`RANDOM}};
  recv_2_data_125 = _RAND_687[7:0];
  _RAND_688 = {1{`RANDOM}};
  recv_2_data_126 = _RAND_688[7:0];
  _RAND_689 = {1{`RANDOM}};
  recv_2_data_127 = _RAND_689[7:0];
  _RAND_690 = {1{`RANDOM}};
  recv_2_data_128 = _RAND_690[7:0];
  _RAND_691 = {1{`RANDOM}};
  recv_2_data_129 = _RAND_691[7:0];
  _RAND_692 = {1{`RANDOM}};
  recv_2_data_130 = _RAND_692[7:0];
  _RAND_693 = {1{`RANDOM}};
  recv_2_data_131 = _RAND_693[7:0];
  _RAND_694 = {1{`RANDOM}};
  recv_2_data_132 = _RAND_694[7:0];
  _RAND_695 = {1{`RANDOM}};
  recv_2_data_133 = _RAND_695[7:0];
  _RAND_696 = {1{`RANDOM}};
  recv_2_data_134 = _RAND_696[7:0];
  _RAND_697 = {1{`RANDOM}};
  recv_2_data_135 = _RAND_697[7:0];
  _RAND_698 = {1{`RANDOM}};
  recv_2_data_136 = _RAND_698[7:0];
  _RAND_699 = {1{`RANDOM}};
  recv_2_data_137 = _RAND_699[7:0];
  _RAND_700 = {1{`RANDOM}};
  recv_2_data_138 = _RAND_700[7:0];
  _RAND_701 = {1{`RANDOM}};
  recv_2_data_139 = _RAND_701[7:0];
  _RAND_702 = {1{`RANDOM}};
  recv_2_data_140 = _RAND_702[7:0];
  _RAND_703 = {1{`RANDOM}};
  recv_2_data_141 = _RAND_703[7:0];
  _RAND_704 = {1{`RANDOM}};
  recv_2_data_142 = _RAND_704[7:0];
  _RAND_705 = {1{`RANDOM}};
  recv_2_data_143 = _RAND_705[7:0];
  _RAND_706 = {1{`RANDOM}};
  recv_2_data_144 = _RAND_706[7:0];
  _RAND_707 = {1{`RANDOM}};
  recv_2_data_145 = _RAND_707[7:0];
  _RAND_708 = {1{`RANDOM}};
  recv_2_data_146 = _RAND_708[7:0];
  _RAND_709 = {1{`RANDOM}};
  recv_2_data_147 = _RAND_709[7:0];
  _RAND_710 = {1{`RANDOM}};
  recv_2_data_148 = _RAND_710[7:0];
  _RAND_711 = {1{`RANDOM}};
  recv_2_data_149 = _RAND_711[7:0];
  _RAND_712 = {1{`RANDOM}};
  recv_2_data_150 = _RAND_712[7:0];
  _RAND_713 = {1{`RANDOM}};
  recv_2_data_151 = _RAND_713[7:0];
  _RAND_714 = {1{`RANDOM}};
  recv_2_data_152 = _RAND_714[7:0];
  _RAND_715 = {1{`RANDOM}};
  recv_2_data_153 = _RAND_715[7:0];
  _RAND_716 = {1{`RANDOM}};
  recv_2_data_154 = _RAND_716[7:0];
  _RAND_717 = {1{`RANDOM}};
  recv_2_data_155 = _RAND_717[7:0];
  _RAND_718 = {1{`RANDOM}};
  recv_2_data_156 = _RAND_718[7:0];
  _RAND_719 = {1{`RANDOM}};
  recv_2_data_157 = _RAND_719[7:0];
  _RAND_720 = {1{`RANDOM}};
  recv_2_data_158 = _RAND_720[7:0];
  _RAND_721 = {1{`RANDOM}};
  recv_2_data_159 = _RAND_721[7:0];
  _RAND_722 = {1{`RANDOM}};
  recv_2_data_160 = _RAND_722[7:0];
  _RAND_723 = {1{`RANDOM}};
  recv_2_data_161 = _RAND_723[7:0];
  _RAND_724 = {1{`RANDOM}};
  recv_2_data_162 = _RAND_724[7:0];
  _RAND_725 = {1{`RANDOM}};
  recv_2_data_163 = _RAND_725[7:0];
  _RAND_726 = {1{`RANDOM}};
  recv_2_data_164 = _RAND_726[7:0];
  _RAND_727 = {1{`RANDOM}};
  recv_2_data_165 = _RAND_727[7:0];
  _RAND_728 = {1{`RANDOM}};
  recv_2_data_166 = _RAND_728[7:0];
  _RAND_729 = {1{`RANDOM}};
  recv_2_data_167 = _RAND_729[7:0];
  _RAND_730 = {1{`RANDOM}};
  recv_2_data_168 = _RAND_730[7:0];
  _RAND_731 = {1{`RANDOM}};
  recv_2_data_169 = _RAND_731[7:0];
  _RAND_732 = {1{`RANDOM}};
  recv_2_data_170 = _RAND_732[7:0];
  _RAND_733 = {1{`RANDOM}};
  recv_2_data_171 = _RAND_733[7:0];
  _RAND_734 = {1{`RANDOM}};
  recv_2_data_172 = _RAND_734[7:0];
  _RAND_735 = {1{`RANDOM}};
  recv_2_data_173 = _RAND_735[7:0];
  _RAND_736 = {1{`RANDOM}};
  recv_2_data_174 = _RAND_736[7:0];
  _RAND_737 = {1{`RANDOM}};
  recv_2_data_175 = _RAND_737[7:0];
  _RAND_738 = {1{`RANDOM}};
  recv_2_data_176 = _RAND_738[7:0];
  _RAND_739 = {1{`RANDOM}};
  recv_2_data_177 = _RAND_739[7:0];
  _RAND_740 = {1{`RANDOM}};
  recv_2_data_178 = _RAND_740[7:0];
  _RAND_741 = {1{`RANDOM}};
  recv_2_data_179 = _RAND_741[7:0];
  _RAND_742 = {1{`RANDOM}};
  recv_2_data_180 = _RAND_742[7:0];
  _RAND_743 = {1{`RANDOM}};
  recv_2_data_181 = _RAND_743[7:0];
  _RAND_744 = {1{`RANDOM}};
  recv_2_data_182 = _RAND_744[7:0];
  _RAND_745 = {1{`RANDOM}};
  recv_2_data_183 = _RAND_745[7:0];
  _RAND_746 = {1{`RANDOM}};
  recv_2_data_184 = _RAND_746[7:0];
  _RAND_747 = {1{`RANDOM}};
  recv_2_data_185 = _RAND_747[7:0];
  _RAND_748 = {1{`RANDOM}};
  recv_2_data_186 = _RAND_748[7:0];
  _RAND_749 = {1{`RANDOM}};
  recv_2_data_187 = _RAND_749[7:0];
  _RAND_750 = {1{`RANDOM}};
  recv_2_data_188 = _RAND_750[7:0];
  _RAND_751 = {1{`RANDOM}};
  recv_2_data_189 = _RAND_751[7:0];
  _RAND_752 = {1{`RANDOM}};
  recv_2_data_190 = _RAND_752[7:0];
  _RAND_753 = {1{`RANDOM}};
  recv_2_data_191 = _RAND_753[7:0];
  _RAND_754 = {1{`RANDOM}};
  recv_2_data_192 = _RAND_754[7:0];
  _RAND_755 = {1{`RANDOM}};
  recv_2_data_193 = _RAND_755[7:0];
  _RAND_756 = {1{`RANDOM}};
  recv_2_data_194 = _RAND_756[7:0];
  _RAND_757 = {1{`RANDOM}};
  recv_2_data_195 = _RAND_757[7:0];
  _RAND_758 = {1{`RANDOM}};
  recv_2_data_196 = _RAND_758[7:0];
  _RAND_759 = {1{`RANDOM}};
  recv_2_data_197 = _RAND_759[7:0];
  _RAND_760 = {1{`RANDOM}};
  recv_2_data_198 = _RAND_760[7:0];
  _RAND_761 = {1{`RANDOM}};
  recv_2_data_199 = _RAND_761[7:0];
  _RAND_762 = {1{`RANDOM}};
  recv_2_data_200 = _RAND_762[7:0];
  _RAND_763 = {1{`RANDOM}};
  recv_2_data_201 = _RAND_763[7:0];
  _RAND_764 = {1{`RANDOM}};
  recv_2_data_202 = _RAND_764[7:0];
  _RAND_765 = {1{`RANDOM}};
  recv_2_data_203 = _RAND_765[7:0];
  _RAND_766 = {1{`RANDOM}};
  recv_2_data_204 = _RAND_766[7:0];
  _RAND_767 = {1{`RANDOM}};
  recv_2_data_205 = _RAND_767[7:0];
  _RAND_768 = {1{`RANDOM}};
  recv_2_data_206 = _RAND_768[7:0];
  _RAND_769 = {1{`RANDOM}};
  recv_2_data_207 = _RAND_769[7:0];
  _RAND_770 = {1{`RANDOM}};
  recv_2_data_208 = _RAND_770[7:0];
  _RAND_771 = {1{`RANDOM}};
  recv_2_data_209 = _RAND_771[7:0];
  _RAND_772 = {1{`RANDOM}};
  recv_2_data_210 = _RAND_772[7:0];
  _RAND_773 = {1{`RANDOM}};
  recv_2_data_211 = _RAND_773[7:0];
  _RAND_774 = {1{`RANDOM}};
  recv_2_data_212 = _RAND_774[7:0];
  _RAND_775 = {1{`RANDOM}};
  recv_2_data_213 = _RAND_775[7:0];
  _RAND_776 = {1{`RANDOM}};
  recv_2_data_214 = _RAND_776[7:0];
  _RAND_777 = {1{`RANDOM}};
  recv_2_data_215 = _RAND_777[7:0];
  _RAND_778 = {1{`RANDOM}};
  recv_2_data_216 = _RAND_778[7:0];
  _RAND_779 = {1{`RANDOM}};
  recv_2_data_217 = _RAND_779[7:0];
  _RAND_780 = {1{`RANDOM}};
  recv_2_data_218 = _RAND_780[7:0];
  _RAND_781 = {1{`RANDOM}};
  recv_2_data_219 = _RAND_781[7:0];
  _RAND_782 = {1{`RANDOM}};
  recv_2_data_220 = _RAND_782[7:0];
  _RAND_783 = {1{`RANDOM}};
  recv_2_data_221 = _RAND_783[7:0];
  _RAND_784 = {1{`RANDOM}};
  recv_2_data_222 = _RAND_784[7:0];
  _RAND_785 = {1{`RANDOM}};
  recv_2_data_223 = _RAND_785[7:0];
  _RAND_786 = {1{`RANDOM}};
  recv_2_data_224 = _RAND_786[7:0];
  _RAND_787 = {1{`RANDOM}};
  recv_2_data_225 = _RAND_787[7:0];
  _RAND_788 = {1{`RANDOM}};
  recv_2_data_226 = _RAND_788[7:0];
  _RAND_789 = {1{`RANDOM}};
  recv_2_data_227 = _RAND_789[7:0];
  _RAND_790 = {1{`RANDOM}};
  recv_2_data_228 = _RAND_790[7:0];
  _RAND_791 = {1{`RANDOM}};
  recv_2_data_229 = _RAND_791[7:0];
  _RAND_792 = {1{`RANDOM}};
  recv_2_data_230 = _RAND_792[7:0];
  _RAND_793 = {1{`RANDOM}};
  recv_2_data_231 = _RAND_793[7:0];
  _RAND_794 = {1{`RANDOM}};
  recv_2_data_232 = _RAND_794[7:0];
  _RAND_795 = {1{`RANDOM}};
  recv_2_data_233 = _RAND_795[7:0];
  _RAND_796 = {1{`RANDOM}};
  recv_2_data_234 = _RAND_796[7:0];
  _RAND_797 = {1{`RANDOM}};
  recv_2_data_235 = _RAND_797[7:0];
  _RAND_798 = {1{`RANDOM}};
  recv_2_data_236 = _RAND_798[7:0];
  _RAND_799 = {1{`RANDOM}};
  recv_2_data_237 = _RAND_799[7:0];
  _RAND_800 = {1{`RANDOM}};
  recv_2_data_238 = _RAND_800[7:0];
  _RAND_801 = {1{`RANDOM}};
  recv_2_data_239 = _RAND_801[7:0];
  _RAND_802 = {1{`RANDOM}};
  recv_2_data_240 = _RAND_802[7:0];
  _RAND_803 = {1{`RANDOM}};
  recv_2_data_241 = _RAND_803[7:0];
  _RAND_804 = {1{`RANDOM}};
  recv_2_data_242 = _RAND_804[7:0];
  _RAND_805 = {1{`RANDOM}};
  recv_2_data_243 = _RAND_805[7:0];
  _RAND_806 = {1{`RANDOM}};
  recv_2_data_244 = _RAND_806[7:0];
  _RAND_807 = {1{`RANDOM}};
  recv_2_data_245 = _RAND_807[7:0];
  _RAND_808 = {1{`RANDOM}};
  recv_2_data_246 = _RAND_808[7:0];
  _RAND_809 = {1{`RANDOM}};
  recv_2_data_247 = _RAND_809[7:0];
  _RAND_810 = {1{`RANDOM}};
  recv_2_data_248 = _RAND_810[7:0];
  _RAND_811 = {1{`RANDOM}};
  recv_2_data_249 = _RAND_811[7:0];
  _RAND_812 = {1{`RANDOM}};
  recv_2_data_250 = _RAND_812[7:0];
  _RAND_813 = {1{`RANDOM}};
  recv_2_data_251 = _RAND_813[7:0];
  _RAND_814 = {1{`RANDOM}};
  recv_2_data_252 = _RAND_814[7:0];
  _RAND_815 = {1{`RANDOM}};
  recv_2_data_253 = _RAND_815[7:0];
  _RAND_816 = {1{`RANDOM}};
  recv_2_data_254 = _RAND_816[7:0];
  _RAND_817 = {1{`RANDOM}};
  recv_2_data_255 = _RAND_817[7:0];
  _RAND_818 = {1{`RANDOM}};
  recv_2_header_0 = _RAND_818[15:0];
  _RAND_819 = {1{`RANDOM}};
  recv_2_header_1 = _RAND_819[15:0];
  _RAND_820 = {1{`RANDOM}};
  recv_2_header_2 = _RAND_820[15:0];
  _RAND_821 = {1{`RANDOM}};
  recv_2_header_3 = _RAND_821[15:0];
  _RAND_822 = {1{`RANDOM}};
  recv_2_header_4 = _RAND_822[15:0];
  _RAND_823 = {1{`RANDOM}};
  recv_2_header_5 = _RAND_823[15:0];
  _RAND_824 = {1{`RANDOM}};
  recv_2_header_6 = _RAND_824[15:0];
  _RAND_825 = {1{`RANDOM}};
  recv_2_header_7 = _RAND_825[15:0];
  _RAND_826 = {1{`RANDOM}};
  recv_2_header_8 = _RAND_826[15:0];
  _RAND_827 = {1{`RANDOM}};
  recv_2_header_9 = _RAND_827[15:0];
  _RAND_828 = {1{`RANDOM}};
  recv_2_header_10 = _RAND_828[15:0];
  _RAND_829 = {1{`RANDOM}};
  recv_2_header_11 = _RAND_829[15:0];
  _RAND_830 = {1{`RANDOM}};
  recv_2_header_12 = _RAND_830[15:0];
  _RAND_831 = {1{`RANDOM}};
  recv_2_header_13 = _RAND_831[15:0];
  _RAND_832 = {1{`RANDOM}};
  recv_2_header_14 = _RAND_832[15:0];
  _RAND_833 = {1{`RANDOM}};
  recv_2_header_15 = _RAND_833[15:0];
  _RAND_834 = {1{`RANDOM}};
  recv_2_parse_current_state = _RAND_834[7:0];
  _RAND_835 = {1{`RANDOM}};
  recv_2_parse_current_offset = _RAND_835[7:0];
  _RAND_836 = {1{`RANDOM}};
  recv_2_parse_transition_field = _RAND_836[15:0];
  _RAND_837 = {1{`RANDOM}};
  recv_2_next_processor_id = _RAND_837[1:0];
  _RAND_838 = {1{`RANDOM}};
  recv_2_next_config_id = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  recv_2_is_valid_processor = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  recv_3_data_0 = _RAND_840[7:0];
  _RAND_841 = {1{`RANDOM}};
  recv_3_data_1 = _RAND_841[7:0];
  _RAND_842 = {1{`RANDOM}};
  recv_3_data_2 = _RAND_842[7:0];
  _RAND_843 = {1{`RANDOM}};
  recv_3_data_3 = _RAND_843[7:0];
  _RAND_844 = {1{`RANDOM}};
  recv_3_data_4 = _RAND_844[7:0];
  _RAND_845 = {1{`RANDOM}};
  recv_3_data_5 = _RAND_845[7:0];
  _RAND_846 = {1{`RANDOM}};
  recv_3_data_6 = _RAND_846[7:0];
  _RAND_847 = {1{`RANDOM}};
  recv_3_data_7 = _RAND_847[7:0];
  _RAND_848 = {1{`RANDOM}};
  recv_3_data_8 = _RAND_848[7:0];
  _RAND_849 = {1{`RANDOM}};
  recv_3_data_9 = _RAND_849[7:0];
  _RAND_850 = {1{`RANDOM}};
  recv_3_data_10 = _RAND_850[7:0];
  _RAND_851 = {1{`RANDOM}};
  recv_3_data_11 = _RAND_851[7:0];
  _RAND_852 = {1{`RANDOM}};
  recv_3_data_12 = _RAND_852[7:0];
  _RAND_853 = {1{`RANDOM}};
  recv_3_data_13 = _RAND_853[7:0];
  _RAND_854 = {1{`RANDOM}};
  recv_3_data_14 = _RAND_854[7:0];
  _RAND_855 = {1{`RANDOM}};
  recv_3_data_15 = _RAND_855[7:0];
  _RAND_856 = {1{`RANDOM}};
  recv_3_data_16 = _RAND_856[7:0];
  _RAND_857 = {1{`RANDOM}};
  recv_3_data_17 = _RAND_857[7:0];
  _RAND_858 = {1{`RANDOM}};
  recv_3_data_18 = _RAND_858[7:0];
  _RAND_859 = {1{`RANDOM}};
  recv_3_data_19 = _RAND_859[7:0];
  _RAND_860 = {1{`RANDOM}};
  recv_3_data_20 = _RAND_860[7:0];
  _RAND_861 = {1{`RANDOM}};
  recv_3_data_21 = _RAND_861[7:0];
  _RAND_862 = {1{`RANDOM}};
  recv_3_data_22 = _RAND_862[7:0];
  _RAND_863 = {1{`RANDOM}};
  recv_3_data_23 = _RAND_863[7:0];
  _RAND_864 = {1{`RANDOM}};
  recv_3_data_24 = _RAND_864[7:0];
  _RAND_865 = {1{`RANDOM}};
  recv_3_data_25 = _RAND_865[7:0];
  _RAND_866 = {1{`RANDOM}};
  recv_3_data_26 = _RAND_866[7:0];
  _RAND_867 = {1{`RANDOM}};
  recv_3_data_27 = _RAND_867[7:0];
  _RAND_868 = {1{`RANDOM}};
  recv_3_data_28 = _RAND_868[7:0];
  _RAND_869 = {1{`RANDOM}};
  recv_3_data_29 = _RAND_869[7:0];
  _RAND_870 = {1{`RANDOM}};
  recv_3_data_30 = _RAND_870[7:0];
  _RAND_871 = {1{`RANDOM}};
  recv_3_data_31 = _RAND_871[7:0];
  _RAND_872 = {1{`RANDOM}};
  recv_3_data_32 = _RAND_872[7:0];
  _RAND_873 = {1{`RANDOM}};
  recv_3_data_33 = _RAND_873[7:0];
  _RAND_874 = {1{`RANDOM}};
  recv_3_data_34 = _RAND_874[7:0];
  _RAND_875 = {1{`RANDOM}};
  recv_3_data_35 = _RAND_875[7:0];
  _RAND_876 = {1{`RANDOM}};
  recv_3_data_36 = _RAND_876[7:0];
  _RAND_877 = {1{`RANDOM}};
  recv_3_data_37 = _RAND_877[7:0];
  _RAND_878 = {1{`RANDOM}};
  recv_3_data_38 = _RAND_878[7:0];
  _RAND_879 = {1{`RANDOM}};
  recv_3_data_39 = _RAND_879[7:0];
  _RAND_880 = {1{`RANDOM}};
  recv_3_data_40 = _RAND_880[7:0];
  _RAND_881 = {1{`RANDOM}};
  recv_3_data_41 = _RAND_881[7:0];
  _RAND_882 = {1{`RANDOM}};
  recv_3_data_42 = _RAND_882[7:0];
  _RAND_883 = {1{`RANDOM}};
  recv_3_data_43 = _RAND_883[7:0];
  _RAND_884 = {1{`RANDOM}};
  recv_3_data_44 = _RAND_884[7:0];
  _RAND_885 = {1{`RANDOM}};
  recv_3_data_45 = _RAND_885[7:0];
  _RAND_886 = {1{`RANDOM}};
  recv_3_data_46 = _RAND_886[7:0];
  _RAND_887 = {1{`RANDOM}};
  recv_3_data_47 = _RAND_887[7:0];
  _RAND_888 = {1{`RANDOM}};
  recv_3_data_48 = _RAND_888[7:0];
  _RAND_889 = {1{`RANDOM}};
  recv_3_data_49 = _RAND_889[7:0];
  _RAND_890 = {1{`RANDOM}};
  recv_3_data_50 = _RAND_890[7:0];
  _RAND_891 = {1{`RANDOM}};
  recv_3_data_51 = _RAND_891[7:0];
  _RAND_892 = {1{`RANDOM}};
  recv_3_data_52 = _RAND_892[7:0];
  _RAND_893 = {1{`RANDOM}};
  recv_3_data_53 = _RAND_893[7:0];
  _RAND_894 = {1{`RANDOM}};
  recv_3_data_54 = _RAND_894[7:0];
  _RAND_895 = {1{`RANDOM}};
  recv_3_data_55 = _RAND_895[7:0];
  _RAND_896 = {1{`RANDOM}};
  recv_3_data_56 = _RAND_896[7:0];
  _RAND_897 = {1{`RANDOM}};
  recv_3_data_57 = _RAND_897[7:0];
  _RAND_898 = {1{`RANDOM}};
  recv_3_data_58 = _RAND_898[7:0];
  _RAND_899 = {1{`RANDOM}};
  recv_3_data_59 = _RAND_899[7:0];
  _RAND_900 = {1{`RANDOM}};
  recv_3_data_60 = _RAND_900[7:0];
  _RAND_901 = {1{`RANDOM}};
  recv_3_data_61 = _RAND_901[7:0];
  _RAND_902 = {1{`RANDOM}};
  recv_3_data_62 = _RAND_902[7:0];
  _RAND_903 = {1{`RANDOM}};
  recv_3_data_63 = _RAND_903[7:0];
  _RAND_904 = {1{`RANDOM}};
  recv_3_data_64 = _RAND_904[7:0];
  _RAND_905 = {1{`RANDOM}};
  recv_3_data_65 = _RAND_905[7:0];
  _RAND_906 = {1{`RANDOM}};
  recv_3_data_66 = _RAND_906[7:0];
  _RAND_907 = {1{`RANDOM}};
  recv_3_data_67 = _RAND_907[7:0];
  _RAND_908 = {1{`RANDOM}};
  recv_3_data_68 = _RAND_908[7:0];
  _RAND_909 = {1{`RANDOM}};
  recv_3_data_69 = _RAND_909[7:0];
  _RAND_910 = {1{`RANDOM}};
  recv_3_data_70 = _RAND_910[7:0];
  _RAND_911 = {1{`RANDOM}};
  recv_3_data_71 = _RAND_911[7:0];
  _RAND_912 = {1{`RANDOM}};
  recv_3_data_72 = _RAND_912[7:0];
  _RAND_913 = {1{`RANDOM}};
  recv_3_data_73 = _RAND_913[7:0];
  _RAND_914 = {1{`RANDOM}};
  recv_3_data_74 = _RAND_914[7:0];
  _RAND_915 = {1{`RANDOM}};
  recv_3_data_75 = _RAND_915[7:0];
  _RAND_916 = {1{`RANDOM}};
  recv_3_data_76 = _RAND_916[7:0];
  _RAND_917 = {1{`RANDOM}};
  recv_3_data_77 = _RAND_917[7:0];
  _RAND_918 = {1{`RANDOM}};
  recv_3_data_78 = _RAND_918[7:0];
  _RAND_919 = {1{`RANDOM}};
  recv_3_data_79 = _RAND_919[7:0];
  _RAND_920 = {1{`RANDOM}};
  recv_3_data_80 = _RAND_920[7:0];
  _RAND_921 = {1{`RANDOM}};
  recv_3_data_81 = _RAND_921[7:0];
  _RAND_922 = {1{`RANDOM}};
  recv_3_data_82 = _RAND_922[7:0];
  _RAND_923 = {1{`RANDOM}};
  recv_3_data_83 = _RAND_923[7:0];
  _RAND_924 = {1{`RANDOM}};
  recv_3_data_84 = _RAND_924[7:0];
  _RAND_925 = {1{`RANDOM}};
  recv_3_data_85 = _RAND_925[7:0];
  _RAND_926 = {1{`RANDOM}};
  recv_3_data_86 = _RAND_926[7:0];
  _RAND_927 = {1{`RANDOM}};
  recv_3_data_87 = _RAND_927[7:0];
  _RAND_928 = {1{`RANDOM}};
  recv_3_data_88 = _RAND_928[7:0];
  _RAND_929 = {1{`RANDOM}};
  recv_3_data_89 = _RAND_929[7:0];
  _RAND_930 = {1{`RANDOM}};
  recv_3_data_90 = _RAND_930[7:0];
  _RAND_931 = {1{`RANDOM}};
  recv_3_data_91 = _RAND_931[7:0];
  _RAND_932 = {1{`RANDOM}};
  recv_3_data_92 = _RAND_932[7:0];
  _RAND_933 = {1{`RANDOM}};
  recv_3_data_93 = _RAND_933[7:0];
  _RAND_934 = {1{`RANDOM}};
  recv_3_data_94 = _RAND_934[7:0];
  _RAND_935 = {1{`RANDOM}};
  recv_3_data_95 = _RAND_935[7:0];
  _RAND_936 = {1{`RANDOM}};
  recv_3_data_96 = _RAND_936[7:0];
  _RAND_937 = {1{`RANDOM}};
  recv_3_data_97 = _RAND_937[7:0];
  _RAND_938 = {1{`RANDOM}};
  recv_3_data_98 = _RAND_938[7:0];
  _RAND_939 = {1{`RANDOM}};
  recv_3_data_99 = _RAND_939[7:0];
  _RAND_940 = {1{`RANDOM}};
  recv_3_data_100 = _RAND_940[7:0];
  _RAND_941 = {1{`RANDOM}};
  recv_3_data_101 = _RAND_941[7:0];
  _RAND_942 = {1{`RANDOM}};
  recv_3_data_102 = _RAND_942[7:0];
  _RAND_943 = {1{`RANDOM}};
  recv_3_data_103 = _RAND_943[7:0];
  _RAND_944 = {1{`RANDOM}};
  recv_3_data_104 = _RAND_944[7:0];
  _RAND_945 = {1{`RANDOM}};
  recv_3_data_105 = _RAND_945[7:0];
  _RAND_946 = {1{`RANDOM}};
  recv_3_data_106 = _RAND_946[7:0];
  _RAND_947 = {1{`RANDOM}};
  recv_3_data_107 = _RAND_947[7:0];
  _RAND_948 = {1{`RANDOM}};
  recv_3_data_108 = _RAND_948[7:0];
  _RAND_949 = {1{`RANDOM}};
  recv_3_data_109 = _RAND_949[7:0];
  _RAND_950 = {1{`RANDOM}};
  recv_3_data_110 = _RAND_950[7:0];
  _RAND_951 = {1{`RANDOM}};
  recv_3_data_111 = _RAND_951[7:0];
  _RAND_952 = {1{`RANDOM}};
  recv_3_data_112 = _RAND_952[7:0];
  _RAND_953 = {1{`RANDOM}};
  recv_3_data_113 = _RAND_953[7:0];
  _RAND_954 = {1{`RANDOM}};
  recv_3_data_114 = _RAND_954[7:0];
  _RAND_955 = {1{`RANDOM}};
  recv_3_data_115 = _RAND_955[7:0];
  _RAND_956 = {1{`RANDOM}};
  recv_3_data_116 = _RAND_956[7:0];
  _RAND_957 = {1{`RANDOM}};
  recv_3_data_117 = _RAND_957[7:0];
  _RAND_958 = {1{`RANDOM}};
  recv_3_data_118 = _RAND_958[7:0];
  _RAND_959 = {1{`RANDOM}};
  recv_3_data_119 = _RAND_959[7:0];
  _RAND_960 = {1{`RANDOM}};
  recv_3_data_120 = _RAND_960[7:0];
  _RAND_961 = {1{`RANDOM}};
  recv_3_data_121 = _RAND_961[7:0];
  _RAND_962 = {1{`RANDOM}};
  recv_3_data_122 = _RAND_962[7:0];
  _RAND_963 = {1{`RANDOM}};
  recv_3_data_123 = _RAND_963[7:0];
  _RAND_964 = {1{`RANDOM}};
  recv_3_data_124 = _RAND_964[7:0];
  _RAND_965 = {1{`RANDOM}};
  recv_3_data_125 = _RAND_965[7:0];
  _RAND_966 = {1{`RANDOM}};
  recv_3_data_126 = _RAND_966[7:0];
  _RAND_967 = {1{`RANDOM}};
  recv_3_data_127 = _RAND_967[7:0];
  _RAND_968 = {1{`RANDOM}};
  recv_3_data_128 = _RAND_968[7:0];
  _RAND_969 = {1{`RANDOM}};
  recv_3_data_129 = _RAND_969[7:0];
  _RAND_970 = {1{`RANDOM}};
  recv_3_data_130 = _RAND_970[7:0];
  _RAND_971 = {1{`RANDOM}};
  recv_3_data_131 = _RAND_971[7:0];
  _RAND_972 = {1{`RANDOM}};
  recv_3_data_132 = _RAND_972[7:0];
  _RAND_973 = {1{`RANDOM}};
  recv_3_data_133 = _RAND_973[7:0];
  _RAND_974 = {1{`RANDOM}};
  recv_3_data_134 = _RAND_974[7:0];
  _RAND_975 = {1{`RANDOM}};
  recv_3_data_135 = _RAND_975[7:0];
  _RAND_976 = {1{`RANDOM}};
  recv_3_data_136 = _RAND_976[7:0];
  _RAND_977 = {1{`RANDOM}};
  recv_3_data_137 = _RAND_977[7:0];
  _RAND_978 = {1{`RANDOM}};
  recv_3_data_138 = _RAND_978[7:0];
  _RAND_979 = {1{`RANDOM}};
  recv_3_data_139 = _RAND_979[7:0];
  _RAND_980 = {1{`RANDOM}};
  recv_3_data_140 = _RAND_980[7:0];
  _RAND_981 = {1{`RANDOM}};
  recv_3_data_141 = _RAND_981[7:0];
  _RAND_982 = {1{`RANDOM}};
  recv_3_data_142 = _RAND_982[7:0];
  _RAND_983 = {1{`RANDOM}};
  recv_3_data_143 = _RAND_983[7:0];
  _RAND_984 = {1{`RANDOM}};
  recv_3_data_144 = _RAND_984[7:0];
  _RAND_985 = {1{`RANDOM}};
  recv_3_data_145 = _RAND_985[7:0];
  _RAND_986 = {1{`RANDOM}};
  recv_3_data_146 = _RAND_986[7:0];
  _RAND_987 = {1{`RANDOM}};
  recv_3_data_147 = _RAND_987[7:0];
  _RAND_988 = {1{`RANDOM}};
  recv_3_data_148 = _RAND_988[7:0];
  _RAND_989 = {1{`RANDOM}};
  recv_3_data_149 = _RAND_989[7:0];
  _RAND_990 = {1{`RANDOM}};
  recv_3_data_150 = _RAND_990[7:0];
  _RAND_991 = {1{`RANDOM}};
  recv_3_data_151 = _RAND_991[7:0];
  _RAND_992 = {1{`RANDOM}};
  recv_3_data_152 = _RAND_992[7:0];
  _RAND_993 = {1{`RANDOM}};
  recv_3_data_153 = _RAND_993[7:0];
  _RAND_994 = {1{`RANDOM}};
  recv_3_data_154 = _RAND_994[7:0];
  _RAND_995 = {1{`RANDOM}};
  recv_3_data_155 = _RAND_995[7:0];
  _RAND_996 = {1{`RANDOM}};
  recv_3_data_156 = _RAND_996[7:0];
  _RAND_997 = {1{`RANDOM}};
  recv_3_data_157 = _RAND_997[7:0];
  _RAND_998 = {1{`RANDOM}};
  recv_3_data_158 = _RAND_998[7:0];
  _RAND_999 = {1{`RANDOM}};
  recv_3_data_159 = _RAND_999[7:0];
  _RAND_1000 = {1{`RANDOM}};
  recv_3_data_160 = _RAND_1000[7:0];
  _RAND_1001 = {1{`RANDOM}};
  recv_3_data_161 = _RAND_1001[7:0];
  _RAND_1002 = {1{`RANDOM}};
  recv_3_data_162 = _RAND_1002[7:0];
  _RAND_1003 = {1{`RANDOM}};
  recv_3_data_163 = _RAND_1003[7:0];
  _RAND_1004 = {1{`RANDOM}};
  recv_3_data_164 = _RAND_1004[7:0];
  _RAND_1005 = {1{`RANDOM}};
  recv_3_data_165 = _RAND_1005[7:0];
  _RAND_1006 = {1{`RANDOM}};
  recv_3_data_166 = _RAND_1006[7:0];
  _RAND_1007 = {1{`RANDOM}};
  recv_3_data_167 = _RAND_1007[7:0];
  _RAND_1008 = {1{`RANDOM}};
  recv_3_data_168 = _RAND_1008[7:0];
  _RAND_1009 = {1{`RANDOM}};
  recv_3_data_169 = _RAND_1009[7:0];
  _RAND_1010 = {1{`RANDOM}};
  recv_3_data_170 = _RAND_1010[7:0];
  _RAND_1011 = {1{`RANDOM}};
  recv_3_data_171 = _RAND_1011[7:0];
  _RAND_1012 = {1{`RANDOM}};
  recv_3_data_172 = _RAND_1012[7:0];
  _RAND_1013 = {1{`RANDOM}};
  recv_3_data_173 = _RAND_1013[7:0];
  _RAND_1014 = {1{`RANDOM}};
  recv_3_data_174 = _RAND_1014[7:0];
  _RAND_1015 = {1{`RANDOM}};
  recv_3_data_175 = _RAND_1015[7:0];
  _RAND_1016 = {1{`RANDOM}};
  recv_3_data_176 = _RAND_1016[7:0];
  _RAND_1017 = {1{`RANDOM}};
  recv_3_data_177 = _RAND_1017[7:0];
  _RAND_1018 = {1{`RANDOM}};
  recv_3_data_178 = _RAND_1018[7:0];
  _RAND_1019 = {1{`RANDOM}};
  recv_3_data_179 = _RAND_1019[7:0];
  _RAND_1020 = {1{`RANDOM}};
  recv_3_data_180 = _RAND_1020[7:0];
  _RAND_1021 = {1{`RANDOM}};
  recv_3_data_181 = _RAND_1021[7:0];
  _RAND_1022 = {1{`RANDOM}};
  recv_3_data_182 = _RAND_1022[7:0];
  _RAND_1023 = {1{`RANDOM}};
  recv_3_data_183 = _RAND_1023[7:0];
  _RAND_1024 = {1{`RANDOM}};
  recv_3_data_184 = _RAND_1024[7:0];
  _RAND_1025 = {1{`RANDOM}};
  recv_3_data_185 = _RAND_1025[7:0];
  _RAND_1026 = {1{`RANDOM}};
  recv_3_data_186 = _RAND_1026[7:0];
  _RAND_1027 = {1{`RANDOM}};
  recv_3_data_187 = _RAND_1027[7:0];
  _RAND_1028 = {1{`RANDOM}};
  recv_3_data_188 = _RAND_1028[7:0];
  _RAND_1029 = {1{`RANDOM}};
  recv_3_data_189 = _RAND_1029[7:0];
  _RAND_1030 = {1{`RANDOM}};
  recv_3_data_190 = _RAND_1030[7:0];
  _RAND_1031 = {1{`RANDOM}};
  recv_3_data_191 = _RAND_1031[7:0];
  _RAND_1032 = {1{`RANDOM}};
  recv_3_data_192 = _RAND_1032[7:0];
  _RAND_1033 = {1{`RANDOM}};
  recv_3_data_193 = _RAND_1033[7:0];
  _RAND_1034 = {1{`RANDOM}};
  recv_3_data_194 = _RAND_1034[7:0];
  _RAND_1035 = {1{`RANDOM}};
  recv_3_data_195 = _RAND_1035[7:0];
  _RAND_1036 = {1{`RANDOM}};
  recv_3_data_196 = _RAND_1036[7:0];
  _RAND_1037 = {1{`RANDOM}};
  recv_3_data_197 = _RAND_1037[7:0];
  _RAND_1038 = {1{`RANDOM}};
  recv_3_data_198 = _RAND_1038[7:0];
  _RAND_1039 = {1{`RANDOM}};
  recv_3_data_199 = _RAND_1039[7:0];
  _RAND_1040 = {1{`RANDOM}};
  recv_3_data_200 = _RAND_1040[7:0];
  _RAND_1041 = {1{`RANDOM}};
  recv_3_data_201 = _RAND_1041[7:0];
  _RAND_1042 = {1{`RANDOM}};
  recv_3_data_202 = _RAND_1042[7:0];
  _RAND_1043 = {1{`RANDOM}};
  recv_3_data_203 = _RAND_1043[7:0];
  _RAND_1044 = {1{`RANDOM}};
  recv_3_data_204 = _RAND_1044[7:0];
  _RAND_1045 = {1{`RANDOM}};
  recv_3_data_205 = _RAND_1045[7:0];
  _RAND_1046 = {1{`RANDOM}};
  recv_3_data_206 = _RAND_1046[7:0];
  _RAND_1047 = {1{`RANDOM}};
  recv_3_data_207 = _RAND_1047[7:0];
  _RAND_1048 = {1{`RANDOM}};
  recv_3_data_208 = _RAND_1048[7:0];
  _RAND_1049 = {1{`RANDOM}};
  recv_3_data_209 = _RAND_1049[7:0];
  _RAND_1050 = {1{`RANDOM}};
  recv_3_data_210 = _RAND_1050[7:0];
  _RAND_1051 = {1{`RANDOM}};
  recv_3_data_211 = _RAND_1051[7:0];
  _RAND_1052 = {1{`RANDOM}};
  recv_3_data_212 = _RAND_1052[7:0];
  _RAND_1053 = {1{`RANDOM}};
  recv_3_data_213 = _RAND_1053[7:0];
  _RAND_1054 = {1{`RANDOM}};
  recv_3_data_214 = _RAND_1054[7:0];
  _RAND_1055 = {1{`RANDOM}};
  recv_3_data_215 = _RAND_1055[7:0];
  _RAND_1056 = {1{`RANDOM}};
  recv_3_data_216 = _RAND_1056[7:0];
  _RAND_1057 = {1{`RANDOM}};
  recv_3_data_217 = _RAND_1057[7:0];
  _RAND_1058 = {1{`RANDOM}};
  recv_3_data_218 = _RAND_1058[7:0];
  _RAND_1059 = {1{`RANDOM}};
  recv_3_data_219 = _RAND_1059[7:0];
  _RAND_1060 = {1{`RANDOM}};
  recv_3_data_220 = _RAND_1060[7:0];
  _RAND_1061 = {1{`RANDOM}};
  recv_3_data_221 = _RAND_1061[7:0];
  _RAND_1062 = {1{`RANDOM}};
  recv_3_data_222 = _RAND_1062[7:0];
  _RAND_1063 = {1{`RANDOM}};
  recv_3_data_223 = _RAND_1063[7:0];
  _RAND_1064 = {1{`RANDOM}};
  recv_3_data_224 = _RAND_1064[7:0];
  _RAND_1065 = {1{`RANDOM}};
  recv_3_data_225 = _RAND_1065[7:0];
  _RAND_1066 = {1{`RANDOM}};
  recv_3_data_226 = _RAND_1066[7:0];
  _RAND_1067 = {1{`RANDOM}};
  recv_3_data_227 = _RAND_1067[7:0];
  _RAND_1068 = {1{`RANDOM}};
  recv_3_data_228 = _RAND_1068[7:0];
  _RAND_1069 = {1{`RANDOM}};
  recv_3_data_229 = _RAND_1069[7:0];
  _RAND_1070 = {1{`RANDOM}};
  recv_3_data_230 = _RAND_1070[7:0];
  _RAND_1071 = {1{`RANDOM}};
  recv_3_data_231 = _RAND_1071[7:0];
  _RAND_1072 = {1{`RANDOM}};
  recv_3_data_232 = _RAND_1072[7:0];
  _RAND_1073 = {1{`RANDOM}};
  recv_3_data_233 = _RAND_1073[7:0];
  _RAND_1074 = {1{`RANDOM}};
  recv_3_data_234 = _RAND_1074[7:0];
  _RAND_1075 = {1{`RANDOM}};
  recv_3_data_235 = _RAND_1075[7:0];
  _RAND_1076 = {1{`RANDOM}};
  recv_3_data_236 = _RAND_1076[7:0];
  _RAND_1077 = {1{`RANDOM}};
  recv_3_data_237 = _RAND_1077[7:0];
  _RAND_1078 = {1{`RANDOM}};
  recv_3_data_238 = _RAND_1078[7:0];
  _RAND_1079 = {1{`RANDOM}};
  recv_3_data_239 = _RAND_1079[7:0];
  _RAND_1080 = {1{`RANDOM}};
  recv_3_data_240 = _RAND_1080[7:0];
  _RAND_1081 = {1{`RANDOM}};
  recv_3_data_241 = _RAND_1081[7:0];
  _RAND_1082 = {1{`RANDOM}};
  recv_3_data_242 = _RAND_1082[7:0];
  _RAND_1083 = {1{`RANDOM}};
  recv_3_data_243 = _RAND_1083[7:0];
  _RAND_1084 = {1{`RANDOM}};
  recv_3_data_244 = _RAND_1084[7:0];
  _RAND_1085 = {1{`RANDOM}};
  recv_3_data_245 = _RAND_1085[7:0];
  _RAND_1086 = {1{`RANDOM}};
  recv_3_data_246 = _RAND_1086[7:0];
  _RAND_1087 = {1{`RANDOM}};
  recv_3_data_247 = _RAND_1087[7:0];
  _RAND_1088 = {1{`RANDOM}};
  recv_3_data_248 = _RAND_1088[7:0];
  _RAND_1089 = {1{`RANDOM}};
  recv_3_data_249 = _RAND_1089[7:0];
  _RAND_1090 = {1{`RANDOM}};
  recv_3_data_250 = _RAND_1090[7:0];
  _RAND_1091 = {1{`RANDOM}};
  recv_3_data_251 = _RAND_1091[7:0];
  _RAND_1092 = {1{`RANDOM}};
  recv_3_data_252 = _RAND_1092[7:0];
  _RAND_1093 = {1{`RANDOM}};
  recv_3_data_253 = _RAND_1093[7:0];
  _RAND_1094 = {1{`RANDOM}};
  recv_3_data_254 = _RAND_1094[7:0];
  _RAND_1095 = {1{`RANDOM}};
  recv_3_data_255 = _RAND_1095[7:0];
  _RAND_1096 = {1{`RANDOM}};
  recv_3_header_0 = _RAND_1096[15:0];
  _RAND_1097 = {1{`RANDOM}};
  recv_3_header_1 = _RAND_1097[15:0];
  _RAND_1098 = {1{`RANDOM}};
  recv_3_header_2 = _RAND_1098[15:0];
  _RAND_1099 = {1{`RANDOM}};
  recv_3_header_3 = _RAND_1099[15:0];
  _RAND_1100 = {1{`RANDOM}};
  recv_3_header_4 = _RAND_1100[15:0];
  _RAND_1101 = {1{`RANDOM}};
  recv_3_header_5 = _RAND_1101[15:0];
  _RAND_1102 = {1{`RANDOM}};
  recv_3_header_6 = _RAND_1102[15:0];
  _RAND_1103 = {1{`RANDOM}};
  recv_3_header_7 = _RAND_1103[15:0];
  _RAND_1104 = {1{`RANDOM}};
  recv_3_header_8 = _RAND_1104[15:0];
  _RAND_1105 = {1{`RANDOM}};
  recv_3_header_9 = _RAND_1105[15:0];
  _RAND_1106 = {1{`RANDOM}};
  recv_3_header_10 = _RAND_1106[15:0];
  _RAND_1107 = {1{`RANDOM}};
  recv_3_header_11 = _RAND_1107[15:0];
  _RAND_1108 = {1{`RANDOM}};
  recv_3_header_12 = _RAND_1108[15:0];
  _RAND_1109 = {1{`RANDOM}};
  recv_3_header_13 = _RAND_1109[15:0];
  _RAND_1110 = {1{`RANDOM}};
  recv_3_header_14 = _RAND_1110[15:0];
  _RAND_1111 = {1{`RANDOM}};
  recv_3_header_15 = _RAND_1111[15:0];
  _RAND_1112 = {1{`RANDOM}};
  recv_3_parse_current_state = _RAND_1112[7:0];
  _RAND_1113 = {1{`RANDOM}};
  recv_3_parse_current_offset = _RAND_1113[7:0];
  _RAND_1114 = {1{`RANDOM}};
  recv_3_parse_transition_field = _RAND_1114[15:0];
  _RAND_1115 = {1{`RANDOM}};
  recv_3_next_processor_id = _RAND_1115[1:0];
  _RAND_1116 = {1{`RANDOM}};
  recv_3_next_config_id = _RAND_1116[0:0];
  _RAND_1117 = {1{`RANDOM}};
  recv_3_is_valid_processor = _RAND_1117[0:0];
  _RAND_1118 = {1{`RANDOM}};
  amplifier_0_0_data_0 = _RAND_1118[7:0];
  _RAND_1119 = {1{`RANDOM}};
  amplifier_0_0_data_1 = _RAND_1119[7:0];
  _RAND_1120 = {1{`RANDOM}};
  amplifier_0_0_data_2 = _RAND_1120[7:0];
  _RAND_1121 = {1{`RANDOM}};
  amplifier_0_0_data_3 = _RAND_1121[7:0];
  _RAND_1122 = {1{`RANDOM}};
  amplifier_0_0_data_4 = _RAND_1122[7:0];
  _RAND_1123 = {1{`RANDOM}};
  amplifier_0_0_data_5 = _RAND_1123[7:0];
  _RAND_1124 = {1{`RANDOM}};
  amplifier_0_0_data_6 = _RAND_1124[7:0];
  _RAND_1125 = {1{`RANDOM}};
  amplifier_0_0_data_7 = _RAND_1125[7:0];
  _RAND_1126 = {1{`RANDOM}};
  amplifier_0_0_data_8 = _RAND_1126[7:0];
  _RAND_1127 = {1{`RANDOM}};
  amplifier_0_0_data_9 = _RAND_1127[7:0];
  _RAND_1128 = {1{`RANDOM}};
  amplifier_0_0_data_10 = _RAND_1128[7:0];
  _RAND_1129 = {1{`RANDOM}};
  amplifier_0_0_data_11 = _RAND_1129[7:0];
  _RAND_1130 = {1{`RANDOM}};
  amplifier_0_0_data_12 = _RAND_1130[7:0];
  _RAND_1131 = {1{`RANDOM}};
  amplifier_0_0_data_13 = _RAND_1131[7:0];
  _RAND_1132 = {1{`RANDOM}};
  amplifier_0_0_data_14 = _RAND_1132[7:0];
  _RAND_1133 = {1{`RANDOM}};
  amplifier_0_0_data_15 = _RAND_1133[7:0];
  _RAND_1134 = {1{`RANDOM}};
  amplifier_0_0_data_16 = _RAND_1134[7:0];
  _RAND_1135 = {1{`RANDOM}};
  amplifier_0_0_data_17 = _RAND_1135[7:0];
  _RAND_1136 = {1{`RANDOM}};
  amplifier_0_0_data_18 = _RAND_1136[7:0];
  _RAND_1137 = {1{`RANDOM}};
  amplifier_0_0_data_19 = _RAND_1137[7:0];
  _RAND_1138 = {1{`RANDOM}};
  amplifier_0_0_data_20 = _RAND_1138[7:0];
  _RAND_1139 = {1{`RANDOM}};
  amplifier_0_0_data_21 = _RAND_1139[7:0];
  _RAND_1140 = {1{`RANDOM}};
  amplifier_0_0_data_22 = _RAND_1140[7:0];
  _RAND_1141 = {1{`RANDOM}};
  amplifier_0_0_data_23 = _RAND_1141[7:0];
  _RAND_1142 = {1{`RANDOM}};
  amplifier_0_0_data_24 = _RAND_1142[7:0];
  _RAND_1143 = {1{`RANDOM}};
  amplifier_0_0_data_25 = _RAND_1143[7:0];
  _RAND_1144 = {1{`RANDOM}};
  amplifier_0_0_data_26 = _RAND_1144[7:0];
  _RAND_1145 = {1{`RANDOM}};
  amplifier_0_0_data_27 = _RAND_1145[7:0];
  _RAND_1146 = {1{`RANDOM}};
  amplifier_0_0_data_28 = _RAND_1146[7:0];
  _RAND_1147 = {1{`RANDOM}};
  amplifier_0_0_data_29 = _RAND_1147[7:0];
  _RAND_1148 = {1{`RANDOM}};
  amplifier_0_0_data_30 = _RAND_1148[7:0];
  _RAND_1149 = {1{`RANDOM}};
  amplifier_0_0_data_31 = _RAND_1149[7:0];
  _RAND_1150 = {1{`RANDOM}};
  amplifier_0_0_data_32 = _RAND_1150[7:0];
  _RAND_1151 = {1{`RANDOM}};
  amplifier_0_0_data_33 = _RAND_1151[7:0];
  _RAND_1152 = {1{`RANDOM}};
  amplifier_0_0_data_34 = _RAND_1152[7:0];
  _RAND_1153 = {1{`RANDOM}};
  amplifier_0_0_data_35 = _RAND_1153[7:0];
  _RAND_1154 = {1{`RANDOM}};
  amplifier_0_0_data_36 = _RAND_1154[7:0];
  _RAND_1155 = {1{`RANDOM}};
  amplifier_0_0_data_37 = _RAND_1155[7:0];
  _RAND_1156 = {1{`RANDOM}};
  amplifier_0_0_data_38 = _RAND_1156[7:0];
  _RAND_1157 = {1{`RANDOM}};
  amplifier_0_0_data_39 = _RAND_1157[7:0];
  _RAND_1158 = {1{`RANDOM}};
  amplifier_0_0_data_40 = _RAND_1158[7:0];
  _RAND_1159 = {1{`RANDOM}};
  amplifier_0_0_data_41 = _RAND_1159[7:0];
  _RAND_1160 = {1{`RANDOM}};
  amplifier_0_0_data_42 = _RAND_1160[7:0];
  _RAND_1161 = {1{`RANDOM}};
  amplifier_0_0_data_43 = _RAND_1161[7:0];
  _RAND_1162 = {1{`RANDOM}};
  amplifier_0_0_data_44 = _RAND_1162[7:0];
  _RAND_1163 = {1{`RANDOM}};
  amplifier_0_0_data_45 = _RAND_1163[7:0];
  _RAND_1164 = {1{`RANDOM}};
  amplifier_0_0_data_46 = _RAND_1164[7:0];
  _RAND_1165 = {1{`RANDOM}};
  amplifier_0_0_data_47 = _RAND_1165[7:0];
  _RAND_1166 = {1{`RANDOM}};
  amplifier_0_0_data_48 = _RAND_1166[7:0];
  _RAND_1167 = {1{`RANDOM}};
  amplifier_0_0_data_49 = _RAND_1167[7:0];
  _RAND_1168 = {1{`RANDOM}};
  amplifier_0_0_data_50 = _RAND_1168[7:0];
  _RAND_1169 = {1{`RANDOM}};
  amplifier_0_0_data_51 = _RAND_1169[7:0];
  _RAND_1170 = {1{`RANDOM}};
  amplifier_0_0_data_52 = _RAND_1170[7:0];
  _RAND_1171 = {1{`RANDOM}};
  amplifier_0_0_data_53 = _RAND_1171[7:0];
  _RAND_1172 = {1{`RANDOM}};
  amplifier_0_0_data_54 = _RAND_1172[7:0];
  _RAND_1173 = {1{`RANDOM}};
  amplifier_0_0_data_55 = _RAND_1173[7:0];
  _RAND_1174 = {1{`RANDOM}};
  amplifier_0_0_data_56 = _RAND_1174[7:0];
  _RAND_1175 = {1{`RANDOM}};
  amplifier_0_0_data_57 = _RAND_1175[7:0];
  _RAND_1176 = {1{`RANDOM}};
  amplifier_0_0_data_58 = _RAND_1176[7:0];
  _RAND_1177 = {1{`RANDOM}};
  amplifier_0_0_data_59 = _RAND_1177[7:0];
  _RAND_1178 = {1{`RANDOM}};
  amplifier_0_0_data_60 = _RAND_1178[7:0];
  _RAND_1179 = {1{`RANDOM}};
  amplifier_0_0_data_61 = _RAND_1179[7:0];
  _RAND_1180 = {1{`RANDOM}};
  amplifier_0_0_data_62 = _RAND_1180[7:0];
  _RAND_1181 = {1{`RANDOM}};
  amplifier_0_0_data_63 = _RAND_1181[7:0];
  _RAND_1182 = {1{`RANDOM}};
  amplifier_0_0_data_64 = _RAND_1182[7:0];
  _RAND_1183 = {1{`RANDOM}};
  amplifier_0_0_data_65 = _RAND_1183[7:0];
  _RAND_1184 = {1{`RANDOM}};
  amplifier_0_0_data_66 = _RAND_1184[7:0];
  _RAND_1185 = {1{`RANDOM}};
  amplifier_0_0_data_67 = _RAND_1185[7:0];
  _RAND_1186 = {1{`RANDOM}};
  amplifier_0_0_data_68 = _RAND_1186[7:0];
  _RAND_1187 = {1{`RANDOM}};
  amplifier_0_0_data_69 = _RAND_1187[7:0];
  _RAND_1188 = {1{`RANDOM}};
  amplifier_0_0_data_70 = _RAND_1188[7:0];
  _RAND_1189 = {1{`RANDOM}};
  amplifier_0_0_data_71 = _RAND_1189[7:0];
  _RAND_1190 = {1{`RANDOM}};
  amplifier_0_0_data_72 = _RAND_1190[7:0];
  _RAND_1191 = {1{`RANDOM}};
  amplifier_0_0_data_73 = _RAND_1191[7:0];
  _RAND_1192 = {1{`RANDOM}};
  amplifier_0_0_data_74 = _RAND_1192[7:0];
  _RAND_1193 = {1{`RANDOM}};
  amplifier_0_0_data_75 = _RAND_1193[7:0];
  _RAND_1194 = {1{`RANDOM}};
  amplifier_0_0_data_76 = _RAND_1194[7:0];
  _RAND_1195 = {1{`RANDOM}};
  amplifier_0_0_data_77 = _RAND_1195[7:0];
  _RAND_1196 = {1{`RANDOM}};
  amplifier_0_0_data_78 = _RAND_1196[7:0];
  _RAND_1197 = {1{`RANDOM}};
  amplifier_0_0_data_79 = _RAND_1197[7:0];
  _RAND_1198 = {1{`RANDOM}};
  amplifier_0_0_data_80 = _RAND_1198[7:0];
  _RAND_1199 = {1{`RANDOM}};
  amplifier_0_0_data_81 = _RAND_1199[7:0];
  _RAND_1200 = {1{`RANDOM}};
  amplifier_0_0_data_82 = _RAND_1200[7:0];
  _RAND_1201 = {1{`RANDOM}};
  amplifier_0_0_data_83 = _RAND_1201[7:0];
  _RAND_1202 = {1{`RANDOM}};
  amplifier_0_0_data_84 = _RAND_1202[7:0];
  _RAND_1203 = {1{`RANDOM}};
  amplifier_0_0_data_85 = _RAND_1203[7:0];
  _RAND_1204 = {1{`RANDOM}};
  amplifier_0_0_data_86 = _RAND_1204[7:0];
  _RAND_1205 = {1{`RANDOM}};
  amplifier_0_0_data_87 = _RAND_1205[7:0];
  _RAND_1206 = {1{`RANDOM}};
  amplifier_0_0_data_88 = _RAND_1206[7:0];
  _RAND_1207 = {1{`RANDOM}};
  amplifier_0_0_data_89 = _RAND_1207[7:0];
  _RAND_1208 = {1{`RANDOM}};
  amplifier_0_0_data_90 = _RAND_1208[7:0];
  _RAND_1209 = {1{`RANDOM}};
  amplifier_0_0_data_91 = _RAND_1209[7:0];
  _RAND_1210 = {1{`RANDOM}};
  amplifier_0_0_data_92 = _RAND_1210[7:0];
  _RAND_1211 = {1{`RANDOM}};
  amplifier_0_0_data_93 = _RAND_1211[7:0];
  _RAND_1212 = {1{`RANDOM}};
  amplifier_0_0_data_94 = _RAND_1212[7:0];
  _RAND_1213 = {1{`RANDOM}};
  amplifier_0_0_data_95 = _RAND_1213[7:0];
  _RAND_1214 = {1{`RANDOM}};
  amplifier_0_0_data_96 = _RAND_1214[7:0];
  _RAND_1215 = {1{`RANDOM}};
  amplifier_0_0_data_97 = _RAND_1215[7:0];
  _RAND_1216 = {1{`RANDOM}};
  amplifier_0_0_data_98 = _RAND_1216[7:0];
  _RAND_1217 = {1{`RANDOM}};
  amplifier_0_0_data_99 = _RAND_1217[7:0];
  _RAND_1218 = {1{`RANDOM}};
  amplifier_0_0_data_100 = _RAND_1218[7:0];
  _RAND_1219 = {1{`RANDOM}};
  amplifier_0_0_data_101 = _RAND_1219[7:0];
  _RAND_1220 = {1{`RANDOM}};
  amplifier_0_0_data_102 = _RAND_1220[7:0];
  _RAND_1221 = {1{`RANDOM}};
  amplifier_0_0_data_103 = _RAND_1221[7:0];
  _RAND_1222 = {1{`RANDOM}};
  amplifier_0_0_data_104 = _RAND_1222[7:0];
  _RAND_1223 = {1{`RANDOM}};
  amplifier_0_0_data_105 = _RAND_1223[7:0];
  _RAND_1224 = {1{`RANDOM}};
  amplifier_0_0_data_106 = _RAND_1224[7:0];
  _RAND_1225 = {1{`RANDOM}};
  amplifier_0_0_data_107 = _RAND_1225[7:0];
  _RAND_1226 = {1{`RANDOM}};
  amplifier_0_0_data_108 = _RAND_1226[7:0];
  _RAND_1227 = {1{`RANDOM}};
  amplifier_0_0_data_109 = _RAND_1227[7:0];
  _RAND_1228 = {1{`RANDOM}};
  amplifier_0_0_data_110 = _RAND_1228[7:0];
  _RAND_1229 = {1{`RANDOM}};
  amplifier_0_0_data_111 = _RAND_1229[7:0];
  _RAND_1230 = {1{`RANDOM}};
  amplifier_0_0_data_112 = _RAND_1230[7:0];
  _RAND_1231 = {1{`RANDOM}};
  amplifier_0_0_data_113 = _RAND_1231[7:0];
  _RAND_1232 = {1{`RANDOM}};
  amplifier_0_0_data_114 = _RAND_1232[7:0];
  _RAND_1233 = {1{`RANDOM}};
  amplifier_0_0_data_115 = _RAND_1233[7:0];
  _RAND_1234 = {1{`RANDOM}};
  amplifier_0_0_data_116 = _RAND_1234[7:0];
  _RAND_1235 = {1{`RANDOM}};
  amplifier_0_0_data_117 = _RAND_1235[7:0];
  _RAND_1236 = {1{`RANDOM}};
  amplifier_0_0_data_118 = _RAND_1236[7:0];
  _RAND_1237 = {1{`RANDOM}};
  amplifier_0_0_data_119 = _RAND_1237[7:0];
  _RAND_1238 = {1{`RANDOM}};
  amplifier_0_0_data_120 = _RAND_1238[7:0];
  _RAND_1239 = {1{`RANDOM}};
  amplifier_0_0_data_121 = _RAND_1239[7:0];
  _RAND_1240 = {1{`RANDOM}};
  amplifier_0_0_data_122 = _RAND_1240[7:0];
  _RAND_1241 = {1{`RANDOM}};
  amplifier_0_0_data_123 = _RAND_1241[7:0];
  _RAND_1242 = {1{`RANDOM}};
  amplifier_0_0_data_124 = _RAND_1242[7:0];
  _RAND_1243 = {1{`RANDOM}};
  amplifier_0_0_data_125 = _RAND_1243[7:0];
  _RAND_1244 = {1{`RANDOM}};
  amplifier_0_0_data_126 = _RAND_1244[7:0];
  _RAND_1245 = {1{`RANDOM}};
  amplifier_0_0_data_127 = _RAND_1245[7:0];
  _RAND_1246 = {1{`RANDOM}};
  amplifier_0_0_data_128 = _RAND_1246[7:0];
  _RAND_1247 = {1{`RANDOM}};
  amplifier_0_0_data_129 = _RAND_1247[7:0];
  _RAND_1248 = {1{`RANDOM}};
  amplifier_0_0_data_130 = _RAND_1248[7:0];
  _RAND_1249 = {1{`RANDOM}};
  amplifier_0_0_data_131 = _RAND_1249[7:0];
  _RAND_1250 = {1{`RANDOM}};
  amplifier_0_0_data_132 = _RAND_1250[7:0];
  _RAND_1251 = {1{`RANDOM}};
  amplifier_0_0_data_133 = _RAND_1251[7:0];
  _RAND_1252 = {1{`RANDOM}};
  amplifier_0_0_data_134 = _RAND_1252[7:0];
  _RAND_1253 = {1{`RANDOM}};
  amplifier_0_0_data_135 = _RAND_1253[7:0];
  _RAND_1254 = {1{`RANDOM}};
  amplifier_0_0_data_136 = _RAND_1254[7:0];
  _RAND_1255 = {1{`RANDOM}};
  amplifier_0_0_data_137 = _RAND_1255[7:0];
  _RAND_1256 = {1{`RANDOM}};
  amplifier_0_0_data_138 = _RAND_1256[7:0];
  _RAND_1257 = {1{`RANDOM}};
  amplifier_0_0_data_139 = _RAND_1257[7:0];
  _RAND_1258 = {1{`RANDOM}};
  amplifier_0_0_data_140 = _RAND_1258[7:0];
  _RAND_1259 = {1{`RANDOM}};
  amplifier_0_0_data_141 = _RAND_1259[7:0];
  _RAND_1260 = {1{`RANDOM}};
  amplifier_0_0_data_142 = _RAND_1260[7:0];
  _RAND_1261 = {1{`RANDOM}};
  amplifier_0_0_data_143 = _RAND_1261[7:0];
  _RAND_1262 = {1{`RANDOM}};
  amplifier_0_0_data_144 = _RAND_1262[7:0];
  _RAND_1263 = {1{`RANDOM}};
  amplifier_0_0_data_145 = _RAND_1263[7:0];
  _RAND_1264 = {1{`RANDOM}};
  amplifier_0_0_data_146 = _RAND_1264[7:0];
  _RAND_1265 = {1{`RANDOM}};
  amplifier_0_0_data_147 = _RAND_1265[7:0];
  _RAND_1266 = {1{`RANDOM}};
  amplifier_0_0_data_148 = _RAND_1266[7:0];
  _RAND_1267 = {1{`RANDOM}};
  amplifier_0_0_data_149 = _RAND_1267[7:0];
  _RAND_1268 = {1{`RANDOM}};
  amplifier_0_0_data_150 = _RAND_1268[7:0];
  _RAND_1269 = {1{`RANDOM}};
  amplifier_0_0_data_151 = _RAND_1269[7:0];
  _RAND_1270 = {1{`RANDOM}};
  amplifier_0_0_data_152 = _RAND_1270[7:0];
  _RAND_1271 = {1{`RANDOM}};
  amplifier_0_0_data_153 = _RAND_1271[7:0];
  _RAND_1272 = {1{`RANDOM}};
  amplifier_0_0_data_154 = _RAND_1272[7:0];
  _RAND_1273 = {1{`RANDOM}};
  amplifier_0_0_data_155 = _RAND_1273[7:0];
  _RAND_1274 = {1{`RANDOM}};
  amplifier_0_0_data_156 = _RAND_1274[7:0];
  _RAND_1275 = {1{`RANDOM}};
  amplifier_0_0_data_157 = _RAND_1275[7:0];
  _RAND_1276 = {1{`RANDOM}};
  amplifier_0_0_data_158 = _RAND_1276[7:0];
  _RAND_1277 = {1{`RANDOM}};
  amplifier_0_0_data_159 = _RAND_1277[7:0];
  _RAND_1278 = {1{`RANDOM}};
  amplifier_0_0_data_160 = _RAND_1278[7:0];
  _RAND_1279 = {1{`RANDOM}};
  amplifier_0_0_data_161 = _RAND_1279[7:0];
  _RAND_1280 = {1{`RANDOM}};
  amplifier_0_0_data_162 = _RAND_1280[7:0];
  _RAND_1281 = {1{`RANDOM}};
  amplifier_0_0_data_163 = _RAND_1281[7:0];
  _RAND_1282 = {1{`RANDOM}};
  amplifier_0_0_data_164 = _RAND_1282[7:0];
  _RAND_1283 = {1{`RANDOM}};
  amplifier_0_0_data_165 = _RAND_1283[7:0];
  _RAND_1284 = {1{`RANDOM}};
  amplifier_0_0_data_166 = _RAND_1284[7:0];
  _RAND_1285 = {1{`RANDOM}};
  amplifier_0_0_data_167 = _RAND_1285[7:0];
  _RAND_1286 = {1{`RANDOM}};
  amplifier_0_0_data_168 = _RAND_1286[7:0];
  _RAND_1287 = {1{`RANDOM}};
  amplifier_0_0_data_169 = _RAND_1287[7:0];
  _RAND_1288 = {1{`RANDOM}};
  amplifier_0_0_data_170 = _RAND_1288[7:0];
  _RAND_1289 = {1{`RANDOM}};
  amplifier_0_0_data_171 = _RAND_1289[7:0];
  _RAND_1290 = {1{`RANDOM}};
  amplifier_0_0_data_172 = _RAND_1290[7:0];
  _RAND_1291 = {1{`RANDOM}};
  amplifier_0_0_data_173 = _RAND_1291[7:0];
  _RAND_1292 = {1{`RANDOM}};
  amplifier_0_0_data_174 = _RAND_1292[7:0];
  _RAND_1293 = {1{`RANDOM}};
  amplifier_0_0_data_175 = _RAND_1293[7:0];
  _RAND_1294 = {1{`RANDOM}};
  amplifier_0_0_data_176 = _RAND_1294[7:0];
  _RAND_1295 = {1{`RANDOM}};
  amplifier_0_0_data_177 = _RAND_1295[7:0];
  _RAND_1296 = {1{`RANDOM}};
  amplifier_0_0_data_178 = _RAND_1296[7:0];
  _RAND_1297 = {1{`RANDOM}};
  amplifier_0_0_data_179 = _RAND_1297[7:0];
  _RAND_1298 = {1{`RANDOM}};
  amplifier_0_0_data_180 = _RAND_1298[7:0];
  _RAND_1299 = {1{`RANDOM}};
  amplifier_0_0_data_181 = _RAND_1299[7:0];
  _RAND_1300 = {1{`RANDOM}};
  amplifier_0_0_data_182 = _RAND_1300[7:0];
  _RAND_1301 = {1{`RANDOM}};
  amplifier_0_0_data_183 = _RAND_1301[7:0];
  _RAND_1302 = {1{`RANDOM}};
  amplifier_0_0_data_184 = _RAND_1302[7:0];
  _RAND_1303 = {1{`RANDOM}};
  amplifier_0_0_data_185 = _RAND_1303[7:0];
  _RAND_1304 = {1{`RANDOM}};
  amplifier_0_0_data_186 = _RAND_1304[7:0];
  _RAND_1305 = {1{`RANDOM}};
  amplifier_0_0_data_187 = _RAND_1305[7:0];
  _RAND_1306 = {1{`RANDOM}};
  amplifier_0_0_data_188 = _RAND_1306[7:0];
  _RAND_1307 = {1{`RANDOM}};
  amplifier_0_0_data_189 = _RAND_1307[7:0];
  _RAND_1308 = {1{`RANDOM}};
  amplifier_0_0_data_190 = _RAND_1308[7:0];
  _RAND_1309 = {1{`RANDOM}};
  amplifier_0_0_data_191 = _RAND_1309[7:0];
  _RAND_1310 = {1{`RANDOM}};
  amplifier_0_0_data_192 = _RAND_1310[7:0];
  _RAND_1311 = {1{`RANDOM}};
  amplifier_0_0_data_193 = _RAND_1311[7:0];
  _RAND_1312 = {1{`RANDOM}};
  amplifier_0_0_data_194 = _RAND_1312[7:0];
  _RAND_1313 = {1{`RANDOM}};
  amplifier_0_0_data_195 = _RAND_1313[7:0];
  _RAND_1314 = {1{`RANDOM}};
  amplifier_0_0_data_196 = _RAND_1314[7:0];
  _RAND_1315 = {1{`RANDOM}};
  amplifier_0_0_data_197 = _RAND_1315[7:0];
  _RAND_1316 = {1{`RANDOM}};
  amplifier_0_0_data_198 = _RAND_1316[7:0];
  _RAND_1317 = {1{`RANDOM}};
  amplifier_0_0_data_199 = _RAND_1317[7:0];
  _RAND_1318 = {1{`RANDOM}};
  amplifier_0_0_data_200 = _RAND_1318[7:0];
  _RAND_1319 = {1{`RANDOM}};
  amplifier_0_0_data_201 = _RAND_1319[7:0];
  _RAND_1320 = {1{`RANDOM}};
  amplifier_0_0_data_202 = _RAND_1320[7:0];
  _RAND_1321 = {1{`RANDOM}};
  amplifier_0_0_data_203 = _RAND_1321[7:0];
  _RAND_1322 = {1{`RANDOM}};
  amplifier_0_0_data_204 = _RAND_1322[7:0];
  _RAND_1323 = {1{`RANDOM}};
  amplifier_0_0_data_205 = _RAND_1323[7:0];
  _RAND_1324 = {1{`RANDOM}};
  amplifier_0_0_data_206 = _RAND_1324[7:0];
  _RAND_1325 = {1{`RANDOM}};
  amplifier_0_0_data_207 = _RAND_1325[7:0];
  _RAND_1326 = {1{`RANDOM}};
  amplifier_0_0_data_208 = _RAND_1326[7:0];
  _RAND_1327 = {1{`RANDOM}};
  amplifier_0_0_data_209 = _RAND_1327[7:0];
  _RAND_1328 = {1{`RANDOM}};
  amplifier_0_0_data_210 = _RAND_1328[7:0];
  _RAND_1329 = {1{`RANDOM}};
  amplifier_0_0_data_211 = _RAND_1329[7:0];
  _RAND_1330 = {1{`RANDOM}};
  amplifier_0_0_data_212 = _RAND_1330[7:0];
  _RAND_1331 = {1{`RANDOM}};
  amplifier_0_0_data_213 = _RAND_1331[7:0];
  _RAND_1332 = {1{`RANDOM}};
  amplifier_0_0_data_214 = _RAND_1332[7:0];
  _RAND_1333 = {1{`RANDOM}};
  amplifier_0_0_data_215 = _RAND_1333[7:0];
  _RAND_1334 = {1{`RANDOM}};
  amplifier_0_0_data_216 = _RAND_1334[7:0];
  _RAND_1335 = {1{`RANDOM}};
  amplifier_0_0_data_217 = _RAND_1335[7:0];
  _RAND_1336 = {1{`RANDOM}};
  amplifier_0_0_data_218 = _RAND_1336[7:0];
  _RAND_1337 = {1{`RANDOM}};
  amplifier_0_0_data_219 = _RAND_1337[7:0];
  _RAND_1338 = {1{`RANDOM}};
  amplifier_0_0_data_220 = _RAND_1338[7:0];
  _RAND_1339 = {1{`RANDOM}};
  amplifier_0_0_data_221 = _RAND_1339[7:0];
  _RAND_1340 = {1{`RANDOM}};
  amplifier_0_0_data_222 = _RAND_1340[7:0];
  _RAND_1341 = {1{`RANDOM}};
  amplifier_0_0_data_223 = _RAND_1341[7:0];
  _RAND_1342 = {1{`RANDOM}};
  amplifier_0_0_data_224 = _RAND_1342[7:0];
  _RAND_1343 = {1{`RANDOM}};
  amplifier_0_0_data_225 = _RAND_1343[7:0];
  _RAND_1344 = {1{`RANDOM}};
  amplifier_0_0_data_226 = _RAND_1344[7:0];
  _RAND_1345 = {1{`RANDOM}};
  amplifier_0_0_data_227 = _RAND_1345[7:0];
  _RAND_1346 = {1{`RANDOM}};
  amplifier_0_0_data_228 = _RAND_1346[7:0];
  _RAND_1347 = {1{`RANDOM}};
  amplifier_0_0_data_229 = _RAND_1347[7:0];
  _RAND_1348 = {1{`RANDOM}};
  amplifier_0_0_data_230 = _RAND_1348[7:0];
  _RAND_1349 = {1{`RANDOM}};
  amplifier_0_0_data_231 = _RAND_1349[7:0];
  _RAND_1350 = {1{`RANDOM}};
  amplifier_0_0_data_232 = _RAND_1350[7:0];
  _RAND_1351 = {1{`RANDOM}};
  amplifier_0_0_data_233 = _RAND_1351[7:0];
  _RAND_1352 = {1{`RANDOM}};
  amplifier_0_0_data_234 = _RAND_1352[7:0];
  _RAND_1353 = {1{`RANDOM}};
  amplifier_0_0_data_235 = _RAND_1353[7:0];
  _RAND_1354 = {1{`RANDOM}};
  amplifier_0_0_data_236 = _RAND_1354[7:0];
  _RAND_1355 = {1{`RANDOM}};
  amplifier_0_0_data_237 = _RAND_1355[7:0];
  _RAND_1356 = {1{`RANDOM}};
  amplifier_0_0_data_238 = _RAND_1356[7:0];
  _RAND_1357 = {1{`RANDOM}};
  amplifier_0_0_data_239 = _RAND_1357[7:0];
  _RAND_1358 = {1{`RANDOM}};
  amplifier_0_0_data_240 = _RAND_1358[7:0];
  _RAND_1359 = {1{`RANDOM}};
  amplifier_0_0_data_241 = _RAND_1359[7:0];
  _RAND_1360 = {1{`RANDOM}};
  amplifier_0_0_data_242 = _RAND_1360[7:0];
  _RAND_1361 = {1{`RANDOM}};
  amplifier_0_0_data_243 = _RAND_1361[7:0];
  _RAND_1362 = {1{`RANDOM}};
  amplifier_0_0_data_244 = _RAND_1362[7:0];
  _RAND_1363 = {1{`RANDOM}};
  amplifier_0_0_data_245 = _RAND_1363[7:0];
  _RAND_1364 = {1{`RANDOM}};
  amplifier_0_0_data_246 = _RAND_1364[7:0];
  _RAND_1365 = {1{`RANDOM}};
  amplifier_0_0_data_247 = _RAND_1365[7:0];
  _RAND_1366 = {1{`RANDOM}};
  amplifier_0_0_data_248 = _RAND_1366[7:0];
  _RAND_1367 = {1{`RANDOM}};
  amplifier_0_0_data_249 = _RAND_1367[7:0];
  _RAND_1368 = {1{`RANDOM}};
  amplifier_0_0_data_250 = _RAND_1368[7:0];
  _RAND_1369 = {1{`RANDOM}};
  amplifier_0_0_data_251 = _RAND_1369[7:0];
  _RAND_1370 = {1{`RANDOM}};
  amplifier_0_0_data_252 = _RAND_1370[7:0];
  _RAND_1371 = {1{`RANDOM}};
  amplifier_0_0_data_253 = _RAND_1371[7:0];
  _RAND_1372 = {1{`RANDOM}};
  amplifier_0_0_data_254 = _RAND_1372[7:0];
  _RAND_1373 = {1{`RANDOM}};
  amplifier_0_0_data_255 = _RAND_1373[7:0];
  _RAND_1374 = {1{`RANDOM}};
  amplifier_0_0_header_0 = _RAND_1374[15:0];
  _RAND_1375 = {1{`RANDOM}};
  amplifier_0_0_header_1 = _RAND_1375[15:0];
  _RAND_1376 = {1{`RANDOM}};
  amplifier_0_0_header_2 = _RAND_1376[15:0];
  _RAND_1377 = {1{`RANDOM}};
  amplifier_0_0_header_3 = _RAND_1377[15:0];
  _RAND_1378 = {1{`RANDOM}};
  amplifier_0_0_header_4 = _RAND_1378[15:0];
  _RAND_1379 = {1{`RANDOM}};
  amplifier_0_0_header_5 = _RAND_1379[15:0];
  _RAND_1380 = {1{`RANDOM}};
  amplifier_0_0_header_6 = _RAND_1380[15:0];
  _RAND_1381 = {1{`RANDOM}};
  amplifier_0_0_header_7 = _RAND_1381[15:0];
  _RAND_1382 = {1{`RANDOM}};
  amplifier_0_0_header_8 = _RAND_1382[15:0];
  _RAND_1383 = {1{`RANDOM}};
  amplifier_0_0_header_9 = _RAND_1383[15:0];
  _RAND_1384 = {1{`RANDOM}};
  amplifier_0_0_header_10 = _RAND_1384[15:0];
  _RAND_1385 = {1{`RANDOM}};
  amplifier_0_0_header_11 = _RAND_1385[15:0];
  _RAND_1386 = {1{`RANDOM}};
  amplifier_0_0_header_12 = _RAND_1386[15:0];
  _RAND_1387 = {1{`RANDOM}};
  amplifier_0_0_header_13 = _RAND_1387[15:0];
  _RAND_1388 = {1{`RANDOM}};
  amplifier_0_0_header_14 = _RAND_1388[15:0];
  _RAND_1389 = {1{`RANDOM}};
  amplifier_0_0_header_15 = _RAND_1389[15:0];
  _RAND_1390 = {1{`RANDOM}};
  amplifier_0_0_parse_current_state = _RAND_1390[7:0];
  _RAND_1391 = {1{`RANDOM}};
  amplifier_0_0_parse_current_offset = _RAND_1391[7:0];
  _RAND_1392 = {1{`RANDOM}};
  amplifier_0_0_parse_transition_field = _RAND_1392[15:0];
  _RAND_1393 = {1{`RANDOM}};
  amplifier_0_0_next_processor_id = _RAND_1393[1:0];
  _RAND_1394 = {1{`RANDOM}};
  amplifier_0_0_next_config_id = _RAND_1394[0:0];
  _RAND_1395 = {1{`RANDOM}};
  amplifier_0_0_is_valid_processor = _RAND_1395[0:0];
  _RAND_1396 = {1{`RANDOM}};
  amplifier_0_1_data_0 = _RAND_1396[7:0];
  _RAND_1397 = {1{`RANDOM}};
  amplifier_0_1_data_1 = _RAND_1397[7:0];
  _RAND_1398 = {1{`RANDOM}};
  amplifier_0_1_data_2 = _RAND_1398[7:0];
  _RAND_1399 = {1{`RANDOM}};
  amplifier_0_1_data_3 = _RAND_1399[7:0];
  _RAND_1400 = {1{`RANDOM}};
  amplifier_0_1_data_4 = _RAND_1400[7:0];
  _RAND_1401 = {1{`RANDOM}};
  amplifier_0_1_data_5 = _RAND_1401[7:0];
  _RAND_1402 = {1{`RANDOM}};
  amplifier_0_1_data_6 = _RAND_1402[7:0];
  _RAND_1403 = {1{`RANDOM}};
  amplifier_0_1_data_7 = _RAND_1403[7:0];
  _RAND_1404 = {1{`RANDOM}};
  amplifier_0_1_data_8 = _RAND_1404[7:0];
  _RAND_1405 = {1{`RANDOM}};
  amplifier_0_1_data_9 = _RAND_1405[7:0];
  _RAND_1406 = {1{`RANDOM}};
  amplifier_0_1_data_10 = _RAND_1406[7:0];
  _RAND_1407 = {1{`RANDOM}};
  amplifier_0_1_data_11 = _RAND_1407[7:0];
  _RAND_1408 = {1{`RANDOM}};
  amplifier_0_1_data_12 = _RAND_1408[7:0];
  _RAND_1409 = {1{`RANDOM}};
  amplifier_0_1_data_13 = _RAND_1409[7:0];
  _RAND_1410 = {1{`RANDOM}};
  amplifier_0_1_data_14 = _RAND_1410[7:0];
  _RAND_1411 = {1{`RANDOM}};
  amplifier_0_1_data_15 = _RAND_1411[7:0];
  _RAND_1412 = {1{`RANDOM}};
  amplifier_0_1_data_16 = _RAND_1412[7:0];
  _RAND_1413 = {1{`RANDOM}};
  amplifier_0_1_data_17 = _RAND_1413[7:0];
  _RAND_1414 = {1{`RANDOM}};
  amplifier_0_1_data_18 = _RAND_1414[7:0];
  _RAND_1415 = {1{`RANDOM}};
  amplifier_0_1_data_19 = _RAND_1415[7:0];
  _RAND_1416 = {1{`RANDOM}};
  amplifier_0_1_data_20 = _RAND_1416[7:0];
  _RAND_1417 = {1{`RANDOM}};
  amplifier_0_1_data_21 = _RAND_1417[7:0];
  _RAND_1418 = {1{`RANDOM}};
  amplifier_0_1_data_22 = _RAND_1418[7:0];
  _RAND_1419 = {1{`RANDOM}};
  amplifier_0_1_data_23 = _RAND_1419[7:0];
  _RAND_1420 = {1{`RANDOM}};
  amplifier_0_1_data_24 = _RAND_1420[7:0];
  _RAND_1421 = {1{`RANDOM}};
  amplifier_0_1_data_25 = _RAND_1421[7:0];
  _RAND_1422 = {1{`RANDOM}};
  amplifier_0_1_data_26 = _RAND_1422[7:0];
  _RAND_1423 = {1{`RANDOM}};
  amplifier_0_1_data_27 = _RAND_1423[7:0];
  _RAND_1424 = {1{`RANDOM}};
  amplifier_0_1_data_28 = _RAND_1424[7:0];
  _RAND_1425 = {1{`RANDOM}};
  amplifier_0_1_data_29 = _RAND_1425[7:0];
  _RAND_1426 = {1{`RANDOM}};
  amplifier_0_1_data_30 = _RAND_1426[7:0];
  _RAND_1427 = {1{`RANDOM}};
  amplifier_0_1_data_31 = _RAND_1427[7:0];
  _RAND_1428 = {1{`RANDOM}};
  amplifier_0_1_data_32 = _RAND_1428[7:0];
  _RAND_1429 = {1{`RANDOM}};
  amplifier_0_1_data_33 = _RAND_1429[7:0];
  _RAND_1430 = {1{`RANDOM}};
  amplifier_0_1_data_34 = _RAND_1430[7:0];
  _RAND_1431 = {1{`RANDOM}};
  amplifier_0_1_data_35 = _RAND_1431[7:0];
  _RAND_1432 = {1{`RANDOM}};
  amplifier_0_1_data_36 = _RAND_1432[7:0];
  _RAND_1433 = {1{`RANDOM}};
  amplifier_0_1_data_37 = _RAND_1433[7:0];
  _RAND_1434 = {1{`RANDOM}};
  amplifier_0_1_data_38 = _RAND_1434[7:0];
  _RAND_1435 = {1{`RANDOM}};
  amplifier_0_1_data_39 = _RAND_1435[7:0];
  _RAND_1436 = {1{`RANDOM}};
  amplifier_0_1_data_40 = _RAND_1436[7:0];
  _RAND_1437 = {1{`RANDOM}};
  amplifier_0_1_data_41 = _RAND_1437[7:0];
  _RAND_1438 = {1{`RANDOM}};
  amplifier_0_1_data_42 = _RAND_1438[7:0];
  _RAND_1439 = {1{`RANDOM}};
  amplifier_0_1_data_43 = _RAND_1439[7:0];
  _RAND_1440 = {1{`RANDOM}};
  amplifier_0_1_data_44 = _RAND_1440[7:0];
  _RAND_1441 = {1{`RANDOM}};
  amplifier_0_1_data_45 = _RAND_1441[7:0];
  _RAND_1442 = {1{`RANDOM}};
  amplifier_0_1_data_46 = _RAND_1442[7:0];
  _RAND_1443 = {1{`RANDOM}};
  amplifier_0_1_data_47 = _RAND_1443[7:0];
  _RAND_1444 = {1{`RANDOM}};
  amplifier_0_1_data_48 = _RAND_1444[7:0];
  _RAND_1445 = {1{`RANDOM}};
  amplifier_0_1_data_49 = _RAND_1445[7:0];
  _RAND_1446 = {1{`RANDOM}};
  amplifier_0_1_data_50 = _RAND_1446[7:0];
  _RAND_1447 = {1{`RANDOM}};
  amplifier_0_1_data_51 = _RAND_1447[7:0];
  _RAND_1448 = {1{`RANDOM}};
  amplifier_0_1_data_52 = _RAND_1448[7:0];
  _RAND_1449 = {1{`RANDOM}};
  amplifier_0_1_data_53 = _RAND_1449[7:0];
  _RAND_1450 = {1{`RANDOM}};
  amplifier_0_1_data_54 = _RAND_1450[7:0];
  _RAND_1451 = {1{`RANDOM}};
  amplifier_0_1_data_55 = _RAND_1451[7:0];
  _RAND_1452 = {1{`RANDOM}};
  amplifier_0_1_data_56 = _RAND_1452[7:0];
  _RAND_1453 = {1{`RANDOM}};
  amplifier_0_1_data_57 = _RAND_1453[7:0];
  _RAND_1454 = {1{`RANDOM}};
  amplifier_0_1_data_58 = _RAND_1454[7:0];
  _RAND_1455 = {1{`RANDOM}};
  amplifier_0_1_data_59 = _RAND_1455[7:0];
  _RAND_1456 = {1{`RANDOM}};
  amplifier_0_1_data_60 = _RAND_1456[7:0];
  _RAND_1457 = {1{`RANDOM}};
  amplifier_0_1_data_61 = _RAND_1457[7:0];
  _RAND_1458 = {1{`RANDOM}};
  amplifier_0_1_data_62 = _RAND_1458[7:0];
  _RAND_1459 = {1{`RANDOM}};
  amplifier_0_1_data_63 = _RAND_1459[7:0];
  _RAND_1460 = {1{`RANDOM}};
  amplifier_0_1_data_64 = _RAND_1460[7:0];
  _RAND_1461 = {1{`RANDOM}};
  amplifier_0_1_data_65 = _RAND_1461[7:0];
  _RAND_1462 = {1{`RANDOM}};
  amplifier_0_1_data_66 = _RAND_1462[7:0];
  _RAND_1463 = {1{`RANDOM}};
  amplifier_0_1_data_67 = _RAND_1463[7:0];
  _RAND_1464 = {1{`RANDOM}};
  amplifier_0_1_data_68 = _RAND_1464[7:0];
  _RAND_1465 = {1{`RANDOM}};
  amplifier_0_1_data_69 = _RAND_1465[7:0];
  _RAND_1466 = {1{`RANDOM}};
  amplifier_0_1_data_70 = _RAND_1466[7:0];
  _RAND_1467 = {1{`RANDOM}};
  amplifier_0_1_data_71 = _RAND_1467[7:0];
  _RAND_1468 = {1{`RANDOM}};
  amplifier_0_1_data_72 = _RAND_1468[7:0];
  _RAND_1469 = {1{`RANDOM}};
  amplifier_0_1_data_73 = _RAND_1469[7:0];
  _RAND_1470 = {1{`RANDOM}};
  amplifier_0_1_data_74 = _RAND_1470[7:0];
  _RAND_1471 = {1{`RANDOM}};
  amplifier_0_1_data_75 = _RAND_1471[7:0];
  _RAND_1472 = {1{`RANDOM}};
  amplifier_0_1_data_76 = _RAND_1472[7:0];
  _RAND_1473 = {1{`RANDOM}};
  amplifier_0_1_data_77 = _RAND_1473[7:0];
  _RAND_1474 = {1{`RANDOM}};
  amplifier_0_1_data_78 = _RAND_1474[7:0];
  _RAND_1475 = {1{`RANDOM}};
  amplifier_0_1_data_79 = _RAND_1475[7:0];
  _RAND_1476 = {1{`RANDOM}};
  amplifier_0_1_data_80 = _RAND_1476[7:0];
  _RAND_1477 = {1{`RANDOM}};
  amplifier_0_1_data_81 = _RAND_1477[7:0];
  _RAND_1478 = {1{`RANDOM}};
  amplifier_0_1_data_82 = _RAND_1478[7:0];
  _RAND_1479 = {1{`RANDOM}};
  amplifier_0_1_data_83 = _RAND_1479[7:0];
  _RAND_1480 = {1{`RANDOM}};
  amplifier_0_1_data_84 = _RAND_1480[7:0];
  _RAND_1481 = {1{`RANDOM}};
  amplifier_0_1_data_85 = _RAND_1481[7:0];
  _RAND_1482 = {1{`RANDOM}};
  amplifier_0_1_data_86 = _RAND_1482[7:0];
  _RAND_1483 = {1{`RANDOM}};
  amplifier_0_1_data_87 = _RAND_1483[7:0];
  _RAND_1484 = {1{`RANDOM}};
  amplifier_0_1_data_88 = _RAND_1484[7:0];
  _RAND_1485 = {1{`RANDOM}};
  amplifier_0_1_data_89 = _RAND_1485[7:0];
  _RAND_1486 = {1{`RANDOM}};
  amplifier_0_1_data_90 = _RAND_1486[7:0];
  _RAND_1487 = {1{`RANDOM}};
  amplifier_0_1_data_91 = _RAND_1487[7:0];
  _RAND_1488 = {1{`RANDOM}};
  amplifier_0_1_data_92 = _RAND_1488[7:0];
  _RAND_1489 = {1{`RANDOM}};
  amplifier_0_1_data_93 = _RAND_1489[7:0];
  _RAND_1490 = {1{`RANDOM}};
  amplifier_0_1_data_94 = _RAND_1490[7:0];
  _RAND_1491 = {1{`RANDOM}};
  amplifier_0_1_data_95 = _RAND_1491[7:0];
  _RAND_1492 = {1{`RANDOM}};
  amplifier_0_1_data_96 = _RAND_1492[7:0];
  _RAND_1493 = {1{`RANDOM}};
  amplifier_0_1_data_97 = _RAND_1493[7:0];
  _RAND_1494 = {1{`RANDOM}};
  amplifier_0_1_data_98 = _RAND_1494[7:0];
  _RAND_1495 = {1{`RANDOM}};
  amplifier_0_1_data_99 = _RAND_1495[7:0];
  _RAND_1496 = {1{`RANDOM}};
  amplifier_0_1_data_100 = _RAND_1496[7:0];
  _RAND_1497 = {1{`RANDOM}};
  amplifier_0_1_data_101 = _RAND_1497[7:0];
  _RAND_1498 = {1{`RANDOM}};
  amplifier_0_1_data_102 = _RAND_1498[7:0];
  _RAND_1499 = {1{`RANDOM}};
  amplifier_0_1_data_103 = _RAND_1499[7:0];
  _RAND_1500 = {1{`RANDOM}};
  amplifier_0_1_data_104 = _RAND_1500[7:0];
  _RAND_1501 = {1{`RANDOM}};
  amplifier_0_1_data_105 = _RAND_1501[7:0];
  _RAND_1502 = {1{`RANDOM}};
  amplifier_0_1_data_106 = _RAND_1502[7:0];
  _RAND_1503 = {1{`RANDOM}};
  amplifier_0_1_data_107 = _RAND_1503[7:0];
  _RAND_1504 = {1{`RANDOM}};
  amplifier_0_1_data_108 = _RAND_1504[7:0];
  _RAND_1505 = {1{`RANDOM}};
  amplifier_0_1_data_109 = _RAND_1505[7:0];
  _RAND_1506 = {1{`RANDOM}};
  amplifier_0_1_data_110 = _RAND_1506[7:0];
  _RAND_1507 = {1{`RANDOM}};
  amplifier_0_1_data_111 = _RAND_1507[7:0];
  _RAND_1508 = {1{`RANDOM}};
  amplifier_0_1_data_112 = _RAND_1508[7:0];
  _RAND_1509 = {1{`RANDOM}};
  amplifier_0_1_data_113 = _RAND_1509[7:0];
  _RAND_1510 = {1{`RANDOM}};
  amplifier_0_1_data_114 = _RAND_1510[7:0];
  _RAND_1511 = {1{`RANDOM}};
  amplifier_0_1_data_115 = _RAND_1511[7:0];
  _RAND_1512 = {1{`RANDOM}};
  amplifier_0_1_data_116 = _RAND_1512[7:0];
  _RAND_1513 = {1{`RANDOM}};
  amplifier_0_1_data_117 = _RAND_1513[7:0];
  _RAND_1514 = {1{`RANDOM}};
  amplifier_0_1_data_118 = _RAND_1514[7:0];
  _RAND_1515 = {1{`RANDOM}};
  amplifier_0_1_data_119 = _RAND_1515[7:0];
  _RAND_1516 = {1{`RANDOM}};
  amplifier_0_1_data_120 = _RAND_1516[7:0];
  _RAND_1517 = {1{`RANDOM}};
  amplifier_0_1_data_121 = _RAND_1517[7:0];
  _RAND_1518 = {1{`RANDOM}};
  amplifier_0_1_data_122 = _RAND_1518[7:0];
  _RAND_1519 = {1{`RANDOM}};
  amplifier_0_1_data_123 = _RAND_1519[7:0];
  _RAND_1520 = {1{`RANDOM}};
  amplifier_0_1_data_124 = _RAND_1520[7:0];
  _RAND_1521 = {1{`RANDOM}};
  amplifier_0_1_data_125 = _RAND_1521[7:0];
  _RAND_1522 = {1{`RANDOM}};
  amplifier_0_1_data_126 = _RAND_1522[7:0];
  _RAND_1523 = {1{`RANDOM}};
  amplifier_0_1_data_127 = _RAND_1523[7:0];
  _RAND_1524 = {1{`RANDOM}};
  amplifier_0_1_data_128 = _RAND_1524[7:0];
  _RAND_1525 = {1{`RANDOM}};
  amplifier_0_1_data_129 = _RAND_1525[7:0];
  _RAND_1526 = {1{`RANDOM}};
  amplifier_0_1_data_130 = _RAND_1526[7:0];
  _RAND_1527 = {1{`RANDOM}};
  amplifier_0_1_data_131 = _RAND_1527[7:0];
  _RAND_1528 = {1{`RANDOM}};
  amplifier_0_1_data_132 = _RAND_1528[7:0];
  _RAND_1529 = {1{`RANDOM}};
  amplifier_0_1_data_133 = _RAND_1529[7:0];
  _RAND_1530 = {1{`RANDOM}};
  amplifier_0_1_data_134 = _RAND_1530[7:0];
  _RAND_1531 = {1{`RANDOM}};
  amplifier_0_1_data_135 = _RAND_1531[7:0];
  _RAND_1532 = {1{`RANDOM}};
  amplifier_0_1_data_136 = _RAND_1532[7:0];
  _RAND_1533 = {1{`RANDOM}};
  amplifier_0_1_data_137 = _RAND_1533[7:0];
  _RAND_1534 = {1{`RANDOM}};
  amplifier_0_1_data_138 = _RAND_1534[7:0];
  _RAND_1535 = {1{`RANDOM}};
  amplifier_0_1_data_139 = _RAND_1535[7:0];
  _RAND_1536 = {1{`RANDOM}};
  amplifier_0_1_data_140 = _RAND_1536[7:0];
  _RAND_1537 = {1{`RANDOM}};
  amplifier_0_1_data_141 = _RAND_1537[7:0];
  _RAND_1538 = {1{`RANDOM}};
  amplifier_0_1_data_142 = _RAND_1538[7:0];
  _RAND_1539 = {1{`RANDOM}};
  amplifier_0_1_data_143 = _RAND_1539[7:0];
  _RAND_1540 = {1{`RANDOM}};
  amplifier_0_1_data_144 = _RAND_1540[7:0];
  _RAND_1541 = {1{`RANDOM}};
  amplifier_0_1_data_145 = _RAND_1541[7:0];
  _RAND_1542 = {1{`RANDOM}};
  amplifier_0_1_data_146 = _RAND_1542[7:0];
  _RAND_1543 = {1{`RANDOM}};
  amplifier_0_1_data_147 = _RAND_1543[7:0];
  _RAND_1544 = {1{`RANDOM}};
  amplifier_0_1_data_148 = _RAND_1544[7:0];
  _RAND_1545 = {1{`RANDOM}};
  amplifier_0_1_data_149 = _RAND_1545[7:0];
  _RAND_1546 = {1{`RANDOM}};
  amplifier_0_1_data_150 = _RAND_1546[7:0];
  _RAND_1547 = {1{`RANDOM}};
  amplifier_0_1_data_151 = _RAND_1547[7:0];
  _RAND_1548 = {1{`RANDOM}};
  amplifier_0_1_data_152 = _RAND_1548[7:0];
  _RAND_1549 = {1{`RANDOM}};
  amplifier_0_1_data_153 = _RAND_1549[7:0];
  _RAND_1550 = {1{`RANDOM}};
  amplifier_0_1_data_154 = _RAND_1550[7:0];
  _RAND_1551 = {1{`RANDOM}};
  amplifier_0_1_data_155 = _RAND_1551[7:0];
  _RAND_1552 = {1{`RANDOM}};
  amplifier_0_1_data_156 = _RAND_1552[7:0];
  _RAND_1553 = {1{`RANDOM}};
  amplifier_0_1_data_157 = _RAND_1553[7:0];
  _RAND_1554 = {1{`RANDOM}};
  amplifier_0_1_data_158 = _RAND_1554[7:0];
  _RAND_1555 = {1{`RANDOM}};
  amplifier_0_1_data_159 = _RAND_1555[7:0];
  _RAND_1556 = {1{`RANDOM}};
  amplifier_0_1_data_160 = _RAND_1556[7:0];
  _RAND_1557 = {1{`RANDOM}};
  amplifier_0_1_data_161 = _RAND_1557[7:0];
  _RAND_1558 = {1{`RANDOM}};
  amplifier_0_1_data_162 = _RAND_1558[7:0];
  _RAND_1559 = {1{`RANDOM}};
  amplifier_0_1_data_163 = _RAND_1559[7:0];
  _RAND_1560 = {1{`RANDOM}};
  amplifier_0_1_data_164 = _RAND_1560[7:0];
  _RAND_1561 = {1{`RANDOM}};
  amplifier_0_1_data_165 = _RAND_1561[7:0];
  _RAND_1562 = {1{`RANDOM}};
  amplifier_0_1_data_166 = _RAND_1562[7:0];
  _RAND_1563 = {1{`RANDOM}};
  amplifier_0_1_data_167 = _RAND_1563[7:0];
  _RAND_1564 = {1{`RANDOM}};
  amplifier_0_1_data_168 = _RAND_1564[7:0];
  _RAND_1565 = {1{`RANDOM}};
  amplifier_0_1_data_169 = _RAND_1565[7:0];
  _RAND_1566 = {1{`RANDOM}};
  amplifier_0_1_data_170 = _RAND_1566[7:0];
  _RAND_1567 = {1{`RANDOM}};
  amplifier_0_1_data_171 = _RAND_1567[7:0];
  _RAND_1568 = {1{`RANDOM}};
  amplifier_0_1_data_172 = _RAND_1568[7:0];
  _RAND_1569 = {1{`RANDOM}};
  amplifier_0_1_data_173 = _RAND_1569[7:0];
  _RAND_1570 = {1{`RANDOM}};
  amplifier_0_1_data_174 = _RAND_1570[7:0];
  _RAND_1571 = {1{`RANDOM}};
  amplifier_0_1_data_175 = _RAND_1571[7:0];
  _RAND_1572 = {1{`RANDOM}};
  amplifier_0_1_data_176 = _RAND_1572[7:0];
  _RAND_1573 = {1{`RANDOM}};
  amplifier_0_1_data_177 = _RAND_1573[7:0];
  _RAND_1574 = {1{`RANDOM}};
  amplifier_0_1_data_178 = _RAND_1574[7:0];
  _RAND_1575 = {1{`RANDOM}};
  amplifier_0_1_data_179 = _RAND_1575[7:0];
  _RAND_1576 = {1{`RANDOM}};
  amplifier_0_1_data_180 = _RAND_1576[7:0];
  _RAND_1577 = {1{`RANDOM}};
  amplifier_0_1_data_181 = _RAND_1577[7:0];
  _RAND_1578 = {1{`RANDOM}};
  amplifier_0_1_data_182 = _RAND_1578[7:0];
  _RAND_1579 = {1{`RANDOM}};
  amplifier_0_1_data_183 = _RAND_1579[7:0];
  _RAND_1580 = {1{`RANDOM}};
  amplifier_0_1_data_184 = _RAND_1580[7:0];
  _RAND_1581 = {1{`RANDOM}};
  amplifier_0_1_data_185 = _RAND_1581[7:0];
  _RAND_1582 = {1{`RANDOM}};
  amplifier_0_1_data_186 = _RAND_1582[7:0];
  _RAND_1583 = {1{`RANDOM}};
  amplifier_0_1_data_187 = _RAND_1583[7:0];
  _RAND_1584 = {1{`RANDOM}};
  amplifier_0_1_data_188 = _RAND_1584[7:0];
  _RAND_1585 = {1{`RANDOM}};
  amplifier_0_1_data_189 = _RAND_1585[7:0];
  _RAND_1586 = {1{`RANDOM}};
  amplifier_0_1_data_190 = _RAND_1586[7:0];
  _RAND_1587 = {1{`RANDOM}};
  amplifier_0_1_data_191 = _RAND_1587[7:0];
  _RAND_1588 = {1{`RANDOM}};
  amplifier_0_1_data_192 = _RAND_1588[7:0];
  _RAND_1589 = {1{`RANDOM}};
  amplifier_0_1_data_193 = _RAND_1589[7:0];
  _RAND_1590 = {1{`RANDOM}};
  amplifier_0_1_data_194 = _RAND_1590[7:0];
  _RAND_1591 = {1{`RANDOM}};
  amplifier_0_1_data_195 = _RAND_1591[7:0];
  _RAND_1592 = {1{`RANDOM}};
  amplifier_0_1_data_196 = _RAND_1592[7:0];
  _RAND_1593 = {1{`RANDOM}};
  amplifier_0_1_data_197 = _RAND_1593[7:0];
  _RAND_1594 = {1{`RANDOM}};
  amplifier_0_1_data_198 = _RAND_1594[7:0];
  _RAND_1595 = {1{`RANDOM}};
  amplifier_0_1_data_199 = _RAND_1595[7:0];
  _RAND_1596 = {1{`RANDOM}};
  amplifier_0_1_data_200 = _RAND_1596[7:0];
  _RAND_1597 = {1{`RANDOM}};
  amplifier_0_1_data_201 = _RAND_1597[7:0];
  _RAND_1598 = {1{`RANDOM}};
  amplifier_0_1_data_202 = _RAND_1598[7:0];
  _RAND_1599 = {1{`RANDOM}};
  amplifier_0_1_data_203 = _RAND_1599[7:0];
  _RAND_1600 = {1{`RANDOM}};
  amplifier_0_1_data_204 = _RAND_1600[7:0];
  _RAND_1601 = {1{`RANDOM}};
  amplifier_0_1_data_205 = _RAND_1601[7:0];
  _RAND_1602 = {1{`RANDOM}};
  amplifier_0_1_data_206 = _RAND_1602[7:0];
  _RAND_1603 = {1{`RANDOM}};
  amplifier_0_1_data_207 = _RAND_1603[7:0];
  _RAND_1604 = {1{`RANDOM}};
  amplifier_0_1_data_208 = _RAND_1604[7:0];
  _RAND_1605 = {1{`RANDOM}};
  amplifier_0_1_data_209 = _RAND_1605[7:0];
  _RAND_1606 = {1{`RANDOM}};
  amplifier_0_1_data_210 = _RAND_1606[7:0];
  _RAND_1607 = {1{`RANDOM}};
  amplifier_0_1_data_211 = _RAND_1607[7:0];
  _RAND_1608 = {1{`RANDOM}};
  amplifier_0_1_data_212 = _RAND_1608[7:0];
  _RAND_1609 = {1{`RANDOM}};
  amplifier_0_1_data_213 = _RAND_1609[7:0];
  _RAND_1610 = {1{`RANDOM}};
  amplifier_0_1_data_214 = _RAND_1610[7:0];
  _RAND_1611 = {1{`RANDOM}};
  amplifier_0_1_data_215 = _RAND_1611[7:0];
  _RAND_1612 = {1{`RANDOM}};
  amplifier_0_1_data_216 = _RAND_1612[7:0];
  _RAND_1613 = {1{`RANDOM}};
  amplifier_0_1_data_217 = _RAND_1613[7:0];
  _RAND_1614 = {1{`RANDOM}};
  amplifier_0_1_data_218 = _RAND_1614[7:0];
  _RAND_1615 = {1{`RANDOM}};
  amplifier_0_1_data_219 = _RAND_1615[7:0];
  _RAND_1616 = {1{`RANDOM}};
  amplifier_0_1_data_220 = _RAND_1616[7:0];
  _RAND_1617 = {1{`RANDOM}};
  amplifier_0_1_data_221 = _RAND_1617[7:0];
  _RAND_1618 = {1{`RANDOM}};
  amplifier_0_1_data_222 = _RAND_1618[7:0];
  _RAND_1619 = {1{`RANDOM}};
  amplifier_0_1_data_223 = _RAND_1619[7:0];
  _RAND_1620 = {1{`RANDOM}};
  amplifier_0_1_data_224 = _RAND_1620[7:0];
  _RAND_1621 = {1{`RANDOM}};
  amplifier_0_1_data_225 = _RAND_1621[7:0];
  _RAND_1622 = {1{`RANDOM}};
  amplifier_0_1_data_226 = _RAND_1622[7:0];
  _RAND_1623 = {1{`RANDOM}};
  amplifier_0_1_data_227 = _RAND_1623[7:0];
  _RAND_1624 = {1{`RANDOM}};
  amplifier_0_1_data_228 = _RAND_1624[7:0];
  _RAND_1625 = {1{`RANDOM}};
  amplifier_0_1_data_229 = _RAND_1625[7:0];
  _RAND_1626 = {1{`RANDOM}};
  amplifier_0_1_data_230 = _RAND_1626[7:0];
  _RAND_1627 = {1{`RANDOM}};
  amplifier_0_1_data_231 = _RAND_1627[7:0];
  _RAND_1628 = {1{`RANDOM}};
  amplifier_0_1_data_232 = _RAND_1628[7:0];
  _RAND_1629 = {1{`RANDOM}};
  amplifier_0_1_data_233 = _RAND_1629[7:0];
  _RAND_1630 = {1{`RANDOM}};
  amplifier_0_1_data_234 = _RAND_1630[7:0];
  _RAND_1631 = {1{`RANDOM}};
  amplifier_0_1_data_235 = _RAND_1631[7:0];
  _RAND_1632 = {1{`RANDOM}};
  amplifier_0_1_data_236 = _RAND_1632[7:0];
  _RAND_1633 = {1{`RANDOM}};
  amplifier_0_1_data_237 = _RAND_1633[7:0];
  _RAND_1634 = {1{`RANDOM}};
  amplifier_0_1_data_238 = _RAND_1634[7:0];
  _RAND_1635 = {1{`RANDOM}};
  amplifier_0_1_data_239 = _RAND_1635[7:0];
  _RAND_1636 = {1{`RANDOM}};
  amplifier_0_1_data_240 = _RAND_1636[7:0];
  _RAND_1637 = {1{`RANDOM}};
  amplifier_0_1_data_241 = _RAND_1637[7:0];
  _RAND_1638 = {1{`RANDOM}};
  amplifier_0_1_data_242 = _RAND_1638[7:0];
  _RAND_1639 = {1{`RANDOM}};
  amplifier_0_1_data_243 = _RAND_1639[7:0];
  _RAND_1640 = {1{`RANDOM}};
  amplifier_0_1_data_244 = _RAND_1640[7:0];
  _RAND_1641 = {1{`RANDOM}};
  amplifier_0_1_data_245 = _RAND_1641[7:0];
  _RAND_1642 = {1{`RANDOM}};
  amplifier_0_1_data_246 = _RAND_1642[7:0];
  _RAND_1643 = {1{`RANDOM}};
  amplifier_0_1_data_247 = _RAND_1643[7:0];
  _RAND_1644 = {1{`RANDOM}};
  amplifier_0_1_data_248 = _RAND_1644[7:0];
  _RAND_1645 = {1{`RANDOM}};
  amplifier_0_1_data_249 = _RAND_1645[7:0];
  _RAND_1646 = {1{`RANDOM}};
  amplifier_0_1_data_250 = _RAND_1646[7:0];
  _RAND_1647 = {1{`RANDOM}};
  amplifier_0_1_data_251 = _RAND_1647[7:0];
  _RAND_1648 = {1{`RANDOM}};
  amplifier_0_1_data_252 = _RAND_1648[7:0];
  _RAND_1649 = {1{`RANDOM}};
  amplifier_0_1_data_253 = _RAND_1649[7:0];
  _RAND_1650 = {1{`RANDOM}};
  amplifier_0_1_data_254 = _RAND_1650[7:0];
  _RAND_1651 = {1{`RANDOM}};
  amplifier_0_1_data_255 = _RAND_1651[7:0];
  _RAND_1652 = {1{`RANDOM}};
  amplifier_0_1_header_0 = _RAND_1652[15:0];
  _RAND_1653 = {1{`RANDOM}};
  amplifier_0_1_header_1 = _RAND_1653[15:0];
  _RAND_1654 = {1{`RANDOM}};
  amplifier_0_1_header_2 = _RAND_1654[15:0];
  _RAND_1655 = {1{`RANDOM}};
  amplifier_0_1_header_3 = _RAND_1655[15:0];
  _RAND_1656 = {1{`RANDOM}};
  amplifier_0_1_header_4 = _RAND_1656[15:0];
  _RAND_1657 = {1{`RANDOM}};
  amplifier_0_1_header_5 = _RAND_1657[15:0];
  _RAND_1658 = {1{`RANDOM}};
  amplifier_0_1_header_6 = _RAND_1658[15:0];
  _RAND_1659 = {1{`RANDOM}};
  amplifier_0_1_header_7 = _RAND_1659[15:0];
  _RAND_1660 = {1{`RANDOM}};
  amplifier_0_1_header_8 = _RAND_1660[15:0];
  _RAND_1661 = {1{`RANDOM}};
  amplifier_0_1_header_9 = _RAND_1661[15:0];
  _RAND_1662 = {1{`RANDOM}};
  amplifier_0_1_header_10 = _RAND_1662[15:0];
  _RAND_1663 = {1{`RANDOM}};
  amplifier_0_1_header_11 = _RAND_1663[15:0];
  _RAND_1664 = {1{`RANDOM}};
  amplifier_0_1_header_12 = _RAND_1664[15:0];
  _RAND_1665 = {1{`RANDOM}};
  amplifier_0_1_header_13 = _RAND_1665[15:0];
  _RAND_1666 = {1{`RANDOM}};
  amplifier_0_1_header_14 = _RAND_1666[15:0];
  _RAND_1667 = {1{`RANDOM}};
  amplifier_0_1_header_15 = _RAND_1667[15:0];
  _RAND_1668 = {1{`RANDOM}};
  amplifier_0_1_parse_current_state = _RAND_1668[7:0];
  _RAND_1669 = {1{`RANDOM}};
  amplifier_0_1_parse_current_offset = _RAND_1669[7:0];
  _RAND_1670 = {1{`RANDOM}};
  amplifier_0_1_parse_transition_field = _RAND_1670[15:0];
  _RAND_1671 = {1{`RANDOM}};
  amplifier_0_1_next_processor_id = _RAND_1671[1:0];
  _RAND_1672 = {1{`RANDOM}};
  amplifier_0_1_next_config_id = _RAND_1672[0:0];
  _RAND_1673 = {1{`RANDOM}};
  amplifier_0_1_is_valid_processor = _RAND_1673[0:0];
  _RAND_1674 = {1{`RANDOM}};
  amplifier_0_2_data_0 = _RAND_1674[7:0];
  _RAND_1675 = {1{`RANDOM}};
  amplifier_0_2_data_1 = _RAND_1675[7:0];
  _RAND_1676 = {1{`RANDOM}};
  amplifier_0_2_data_2 = _RAND_1676[7:0];
  _RAND_1677 = {1{`RANDOM}};
  amplifier_0_2_data_3 = _RAND_1677[7:0];
  _RAND_1678 = {1{`RANDOM}};
  amplifier_0_2_data_4 = _RAND_1678[7:0];
  _RAND_1679 = {1{`RANDOM}};
  amplifier_0_2_data_5 = _RAND_1679[7:0];
  _RAND_1680 = {1{`RANDOM}};
  amplifier_0_2_data_6 = _RAND_1680[7:0];
  _RAND_1681 = {1{`RANDOM}};
  amplifier_0_2_data_7 = _RAND_1681[7:0];
  _RAND_1682 = {1{`RANDOM}};
  amplifier_0_2_data_8 = _RAND_1682[7:0];
  _RAND_1683 = {1{`RANDOM}};
  amplifier_0_2_data_9 = _RAND_1683[7:0];
  _RAND_1684 = {1{`RANDOM}};
  amplifier_0_2_data_10 = _RAND_1684[7:0];
  _RAND_1685 = {1{`RANDOM}};
  amplifier_0_2_data_11 = _RAND_1685[7:0];
  _RAND_1686 = {1{`RANDOM}};
  amplifier_0_2_data_12 = _RAND_1686[7:0];
  _RAND_1687 = {1{`RANDOM}};
  amplifier_0_2_data_13 = _RAND_1687[7:0];
  _RAND_1688 = {1{`RANDOM}};
  amplifier_0_2_data_14 = _RAND_1688[7:0];
  _RAND_1689 = {1{`RANDOM}};
  amplifier_0_2_data_15 = _RAND_1689[7:0];
  _RAND_1690 = {1{`RANDOM}};
  amplifier_0_2_data_16 = _RAND_1690[7:0];
  _RAND_1691 = {1{`RANDOM}};
  amplifier_0_2_data_17 = _RAND_1691[7:0];
  _RAND_1692 = {1{`RANDOM}};
  amplifier_0_2_data_18 = _RAND_1692[7:0];
  _RAND_1693 = {1{`RANDOM}};
  amplifier_0_2_data_19 = _RAND_1693[7:0];
  _RAND_1694 = {1{`RANDOM}};
  amplifier_0_2_data_20 = _RAND_1694[7:0];
  _RAND_1695 = {1{`RANDOM}};
  amplifier_0_2_data_21 = _RAND_1695[7:0];
  _RAND_1696 = {1{`RANDOM}};
  amplifier_0_2_data_22 = _RAND_1696[7:0];
  _RAND_1697 = {1{`RANDOM}};
  amplifier_0_2_data_23 = _RAND_1697[7:0];
  _RAND_1698 = {1{`RANDOM}};
  amplifier_0_2_data_24 = _RAND_1698[7:0];
  _RAND_1699 = {1{`RANDOM}};
  amplifier_0_2_data_25 = _RAND_1699[7:0];
  _RAND_1700 = {1{`RANDOM}};
  amplifier_0_2_data_26 = _RAND_1700[7:0];
  _RAND_1701 = {1{`RANDOM}};
  amplifier_0_2_data_27 = _RAND_1701[7:0];
  _RAND_1702 = {1{`RANDOM}};
  amplifier_0_2_data_28 = _RAND_1702[7:0];
  _RAND_1703 = {1{`RANDOM}};
  amplifier_0_2_data_29 = _RAND_1703[7:0];
  _RAND_1704 = {1{`RANDOM}};
  amplifier_0_2_data_30 = _RAND_1704[7:0];
  _RAND_1705 = {1{`RANDOM}};
  amplifier_0_2_data_31 = _RAND_1705[7:0];
  _RAND_1706 = {1{`RANDOM}};
  amplifier_0_2_data_32 = _RAND_1706[7:0];
  _RAND_1707 = {1{`RANDOM}};
  amplifier_0_2_data_33 = _RAND_1707[7:0];
  _RAND_1708 = {1{`RANDOM}};
  amplifier_0_2_data_34 = _RAND_1708[7:0];
  _RAND_1709 = {1{`RANDOM}};
  amplifier_0_2_data_35 = _RAND_1709[7:0];
  _RAND_1710 = {1{`RANDOM}};
  amplifier_0_2_data_36 = _RAND_1710[7:0];
  _RAND_1711 = {1{`RANDOM}};
  amplifier_0_2_data_37 = _RAND_1711[7:0];
  _RAND_1712 = {1{`RANDOM}};
  amplifier_0_2_data_38 = _RAND_1712[7:0];
  _RAND_1713 = {1{`RANDOM}};
  amplifier_0_2_data_39 = _RAND_1713[7:0];
  _RAND_1714 = {1{`RANDOM}};
  amplifier_0_2_data_40 = _RAND_1714[7:0];
  _RAND_1715 = {1{`RANDOM}};
  amplifier_0_2_data_41 = _RAND_1715[7:0];
  _RAND_1716 = {1{`RANDOM}};
  amplifier_0_2_data_42 = _RAND_1716[7:0];
  _RAND_1717 = {1{`RANDOM}};
  amplifier_0_2_data_43 = _RAND_1717[7:0];
  _RAND_1718 = {1{`RANDOM}};
  amplifier_0_2_data_44 = _RAND_1718[7:0];
  _RAND_1719 = {1{`RANDOM}};
  amplifier_0_2_data_45 = _RAND_1719[7:0];
  _RAND_1720 = {1{`RANDOM}};
  amplifier_0_2_data_46 = _RAND_1720[7:0];
  _RAND_1721 = {1{`RANDOM}};
  amplifier_0_2_data_47 = _RAND_1721[7:0];
  _RAND_1722 = {1{`RANDOM}};
  amplifier_0_2_data_48 = _RAND_1722[7:0];
  _RAND_1723 = {1{`RANDOM}};
  amplifier_0_2_data_49 = _RAND_1723[7:0];
  _RAND_1724 = {1{`RANDOM}};
  amplifier_0_2_data_50 = _RAND_1724[7:0];
  _RAND_1725 = {1{`RANDOM}};
  amplifier_0_2_data_51 = _RAND_1725[7:0];
  _RAND_1726 = {1{`RANDOM}};
  amplifier_0_2_data_52 = _RAND_1726[7:0];
  _RAND_1727 = {1{`RANDOM}};
  amplifier_0_2_data_53 = _RAND_1727[7:0];
  _RAND_1728 = {1{`RANDOM}};
  amplifier_0_2_data_54 = _RAND_1728[7:0];
  _RAND_1729 = {1{`RANDOM}};
  amplifier_0_2_data_55 = _RAND_1729[7:0];
  _RAND_1730 = {1{`RANDOM}};
  amplifier_0_2_data_56 = _RAND_1730[7:0];
  _RAND_1731 = {1{`RANDOM}};
  amplifier_0_2_data_57 = _RAND_1731[7:0];
  _RAND_1732 = {1{`RANDOM}};
  amplifier_0_2_data_58 = _RAND_1732[7:0];
  _RAND_1733 = {1{`RANDOM}};
  amplifier_0_2_data_59 = _RAND_1733[7:0];
  _RAND_1734 = {1{`RANDOM}};
  amplifier_0_2_data_60 = _RAND_1734[7:0];
  _RAND_1735 = {1{`RANDOM}};
  amplifier_0_2_data_61 = _RAND_1735[7:0];
  _RAND_1736 = {1{`RANDOM}};
  amplifier_0_2_data_62 = _RAND_1736[7:0];
  _RAND_1737 = {1{`RANDOM}};
  amplifier_0_2_data_63 = _RAND_1737[7:0];
  _RAND_1738 = {1{`RANDOM}};
  amplifier_0_2_data_64 = _RAND_1738[7:0];
  _RAND_1739 = {1{`RANDOM}};
  amplifier_0_2_data_65 = _RAND_1739[7:0];
  _RAND_1740 = {1{`RANDOM}};
  amplifier_0_2_data_66 = _RAND_1740[7:0];
  _RAND_1741 = {1{`RANDOM}};
  amplifier_0_2_data_67 = _RAND_1741[7:0];
  _RAND_1742 = {1{`RANDOM}};
  amplifier_0_2_data_68 = _RAND_1742[7:0];
  _RAND_1743 = {1{`RANDOM}};
  amplifier_0_2_data_69 = _RAND_1743[7:0];
  _RAND_1744 = {1{`RANDOM}};
  amplifier_0_2_data_70 = _RAND_1744[7:0];
  _RAND_1745 = {1{`RANDOM}};
  amplifier_0_2_data_71 = _RAND_1745[7:0];
  _RAND_1746 = {1{`RANDOM}};
  amplifier_0_2_data_72 = _RAND_1746[7:0];
  _RAND_1747 = {1{`RANDOM}};
  amplifier_0_2_data_73 = _RAND_1747[7:0];
  _RAND_1748 = {1{`RANDOM}};
  amplifier_0_2_data_74 = _RAND_1748[7:0];
  _RAND_1749 = {1{`RANDOM}};
  amplifier_0_2_data_75 = _RAND_1749[7:0];
  _RAND_1750 = {1{`RANDOM}};
  amplifier_0_2_data_76 = _RAND_1750[7:0];
  _RAND_1751 = {1{`RANDOM}};
  amplifier_0_2_data_77 = _RAND_1751[7:0];
  _RAND_1752 = {1{`RANDOM}};
  amplifier_0_2_data_78 = _RAND_1752[7:0];
  _RAND_1753 = {1{`RANDOM}};
  amplifier_0_2_data_79 = _RAND_1753[7:0];
  _RAND_1754 = {1{`RANDOM}};
  amplifier_0_2_data_80 = _RAND_1754[7:0];
  _RAND_1755 = {1{`RANDOM}};
  amplifier_0_2_data_81 = _RAND_1755[7:0];
  _RAND_1756 = {1{`RANDOM}};
  amplifier_0_2_data_82 = _RAND_1756[7:0];
  _RAND_1757 = {1{`RANDOM}};
  amplifier_0_2_data_83 = _RAND_1757[7:0];
  _RAND_1758 = {1{`RANDOM}};
  amplifier_0_2_data_84 = _RAND_1758[7:0];
  _RAND_1759 = {1{`RANDOM}};
  amplifier_0_2_data_85 = _RAND_1759[7:0];
  _RAND_1760 = {1{`RANDOM}};
  amplifier_0_2_data_86 = _RAND_1760[7:0];
  _RAND_1761 = {1{`RANDOM}};
  amplifier_0_2_data_87 = _RAND_1761[7:0];
  _RAND_1762 = {1{`RANDOM}};
  amplifier_0_2_data_88 = _RAND_1762[7:0];
  _RAND_1763 = {1{`RANDOM}};
  amplifier_0_2_data_89 = _RAND_1763[7:0];
  _RAND_1764 = {1{`RANDOM}};
  amplifier_0_2_data_90 = _RAND_1764[7:0];
  _RAND_1765 = {1{`RANDOM}};
  amplifier_0_2_data_91 = _RAND_1765[7:0];
  _RAND_1766 = {1{`RANDOM}};
  amplifier_0_2_data_92 = _RAND_1766[7:0];
  _RAND_1767 = {1{`RANDOM}};
  amplifier_0_2_data_93 = _RAND_1767[7:0];
  _RAND_1768 = {1{`RANDOM}};
  amplifier_0_2_data_94 = _RAND_1768[7:0];
  _RAND_1769 = {1{`RANDOM}};
  amplifier_0_2_data_95 = _RAND_1769[7:0];
  _RAND_1770 = {1{`RANDOM}};
  amplifier_0_2_data_96 = _RAND_1770[7:0];
  _RAND_1771 = {1{`RANDOM}};
  amplifier_0_2_data_97 = _RAND_1771[7:0];
  _RAND_1772 = {1{`RANDOM}};
  amplifier_0_2_data_98 = _RAND_1772[7:0];
  _RAND_1773 = {1{`RANDOM}};
  amplifier_0_2_data_99 = _RAND_1773[7:0];
  _RAND_1774 = {1{`RANDOM}};
  amplifier_0_2_data_100 = _RAND_1774[7:0];
  _RAND_1775 = {1{`RANDOM}};
  amplifier_0_2_data_101 = _RAND_1775[7:0];
  _RAND_1776 = {1{`RANDOM}};
  amplifier_0_2_data_102 = _RAND_1776[7:0];
  _RAND_1777 = {1{`RANDOM}};
  amplifier_0_2_data_103 = _RAND_1777[7:0];
  _RAND_1778 = {1{`RANDOM}};
  amplifier_0_2_data_104 = _RAND_1778[7:0];
  _RAND_1779 = {1{`RANDOM}};
  amplifier_0_2_data_105 = _RAND_1779[7:0];
  _RAND_1780 = {1{`RANDOM}};
  amplifier_0_2_data_106 = _RAND_1780[7:0];
  _RAND_1781 = {1{`RANDOM}};
  amplifier_0_2_data_107 = _RAND_1781[7:0];
  _RAND_1782 = {1{`RANDOM}};
  amplifier_0_2_data_108 = _RAND_1782[7:0];
  _RAND_1783 = {1{`RANDOM}};
  amplifier_0_2_data_109 = _RAND_1783[7:0];
  _RAND_1784 = {1{`RANDOM}};
  amplifier_0_2_data_110 = _RAND_1784[7:0];
  _RAND_1785 = {1{`RANDOM}};
  amplifier_0_2_data_111 = _RAND_1785[7:0];
  _RAND_1786 = {1{`RANDOM}};
  amplifier_0_2_data_112 = _RAND_1786[7:0];
  _RAND_1787 = {1{`RANDOM}};
  amplifier_0_2_data_113 = _RAND_1787[7:0];
  _RAND_1788 = {1{`RANDOM}};
  amplifier_0_2_data_114 = _RAND_1788[7:0];
  _RAND_1789 = {1{`RANDOM}};
  amplifier_0_2_data_115 = _RAND_1789[7:0];
  _RAND_1790 = {1{`RANDOM}};
  amplifier_0_2_data_116 = _RAND_1790[7:0];
  _RAND_1791 = {1{`RANDOM}};
  amplifier_0_2_data_117 = _RAND_1791[7:0];
  _RAND_1792 = {1{`RANDOM}};
  amplifier_0_2_data_118 = _RAND_1792[7:0];
  _RAND_1793 = {1{`RANDOM}};
  amplifier_0_2_data_119 = _RAND_1793[7:0];
  _RAND_1794 = {1{`RANDOM}};
  amplifier_0_2_data_120 = _RAND_1794[7:0];
  _RAND_1795 = {1{`RANDOM}};
  amplifier_0_2_data_121 = _RAND_1795[7:0];
  _RAND_1796 = {1{`RANDOM}};
  amplifier_0_2_data_122 = _RAND_1796[7:0];
  _RAND_1797 = {1{`RANDOM}};
  amplifier_0_2_data_123 = _RAND_1797[7:0];
  _RAND_1798 = {1{`RANDOM}};
  amplifier_0_2_data_124 = _RAND_1798[7:0];
  _RAND_1799 = {1{`RANDOM}};
  amplifier_0_2_data_125 = _RAND_1799[7:0];
  _RAND_1800 = {1{`RANDOM}};
  amplifier_0_2_data_126 = _RAND_1800[7:0];
  _RAND_1801 = {1{`RANDOM}};
  amplifier_0_2_data_127 = _RAND_1801[7:0];
  _RAND_1802 = {1{`RANDOM}};
  amplifier_0_2_data_128 = _RAND_1802[7:0];
  _RAND_1803 = {1{`RANDOM}};
  amplifier_0_2_data_129 = _RAND_1803[7:0];
  _RAND_1804 = {1{`RANDOM}};
  amplifier_0_2_data_130 = _RAND_1804[7:0];
  _RAND_1805 = {1{`RANDOM}};
  amplifier_0_2_data_131 = _RAND_1805[7:0];
  _RAND_1806 = {1{`RANDOM}};
  amplifier_0_2_data_132 = _RAND_1806[7:0];
  _RAND_1807 = {1{`RANDOM}};
  amplifier_0_2_data_133 = _RAND_1807[7:0];
  _RAND_1808 = {1{`RANDOM}};
  amplifier_0_2_data_134 = _RAND_1808[7:0];
  _RAND_1809 = {1{`RANDOM}};
  amplifier_0_2_data_135 = _RAND_1809[7:0];
  _RAND_1810 = {1{`RANDOM}};
  amplifier_0_2_data_136 = _RAND_1810[7:0];
  _RAND_1811 = {1{`RANDOM}};
  amplifier_0_2_data_137 = _RAND_1811[7:0];
  _RAND_1812 = {1{`RANDOM}};
  amplifier_0_2_data_138 = _RAND_1812[7:0];
  _RAND_1813 = {1{`RANDOM}};
  amplifier_0_2_data_139 = _RAND_1813[7:0];
  _RAND_1814 = {1{`RANDOM}};
  amplifier_0_2_data_140 = _RAND_1814[7:0];
  _RAND_1815 = {1{`RANDOM}};
  amplifier_0_2_data_141 = _RAND_1815[7:0];
  _RAND_1816 = {1{`RANDOM}};
  amplifier_0_2_data_142 = _RAND_1816[7:0];
  _RAND_1817 = {1{`RANDOM}};
  amplifier_0_2_data_143 = _RAND_1817[7:0];
  _RAND_1818 = {1{`RANDOM}};
  amplifier_0_2_data_144 = _RAND_1818[7:0];
  _RAND_1819 = {1{`RANDOM}};
  amplifier_0_2_data_145 = _RAND_1819[7:0];
  _RAND_1820 = {1{`RANDOM}};
  amplifier_0_2_data_146 = _RAND_1820[7:0];
  _RAND_1821 = {1{`RANDOM}};
  amplifier_0_2_data_147 = _RAND_1821[7:0];
  _RAND_1822 = {1{`RANDOM}};
  amplifier_0_2_data_148 = _RAND_1822[7:0];
  _RAND_1823 = {1{`RANDOM}};
  amplifier_0_2_data_149 = _RAND_1823[7:0];
  _RAND_1824 = {1{`RANDOM}};
  amplifier_0_2_data_150 = _RAND_1824[7:0];
  _RAND_1825 = {1{`RANDOM}};
  amplifier_0_2_data_151 = _RAND_1825[7:0];
  _RAND_1826 = {1{`RANDOM}};
  amplifier_0_2_data_152 = _RAND_1826[7:0];
  _RAND_1827 = {1{`RANDOM}};
  amplifier_0_2_data_153 = _RAND_1827[7:0];
  _RAND_1828 = {1{`RANDOM}};
  amplifier_0_2_data_154 = _RAND_1828[7:0];
  _RAND_1829 = {1{`RANDOM}};
  amplifier_0_2_data_155 = _RAND_1829[7:0];
  _RAND_1830 = {1{`RANDOM}};
  amplifier_0_2_data_156 = _RAND_1830[7:0];
  _RAND_1831 = {1{`RANDOM}};
  amplifier_0_2_data_157 = _RAND_1831[7:0];
  _RAND_1832 = {1{`RANDOM}};
  amplifier_0_2_data_158 = _RAND_1832[7:0];
  _RAND_1833 = {1{`RANDOM}};
  amplifier_0_2_data_159 = _RAND_1833[7:0];
  _RAND_1834 = {1{`RANDOM}};
  amplifier_0_2_data_160 = _RAND_1834[7:0];
  _RAND_1835 = {1{`RANDOM}};
  amplifier_0_2_data_161 = _RAND_1835[7:0];
  _RAND_1836 = {1{`RANDOM}};
  amplifier_0_2_data_162 = _RAND_1836[7:0];
  _RAND_1837 = {1{`RANDOM}};
  amplifier_0_2_data_163 = _RAND_1837[7:0];
  _RAND_1838 = {1{`RANDOM}};
  amplifier_0_2_data_164 = _RAND_1838[7:0];
  _RAND_1839 = {1{`RANDOM}};
  amplifier_0_2_data_165 = _RAND_1839[7:0];
  _RAND_1840 = {1{`RANDOM}};
  amplifier_0_2_data_166 = _RAND_1840[7:0];
  _RAND_1841 = {1{`RANDOM}};
  amplifier_0_2_data_167 = _RAND_1841[7:0];
  _RAND_1842 = {1{`RANDOM}};
  amplifier_0_2_data_168 = _RAND_1842[7:0];
  _RAND_1843 = {1{`RANDOM}};
  amplifier_0_2_data_169 = _RAND_1843[7:0];
  _RAND_1844 = {1{`RANDOM}};
  amplifier_0_2_data_170 = _RAND_1844[7:0];
  _RAND_1845 = {1{`RANDOM}};
  amplifier_0_2_data_171 = _RAND_1845[7:0];
  _RAND_1846 = {1{`RANDOM}};
  amplifier_0_2_data_172 = _RAND_1846[7:0];
  _RAND_1847 = {1{`RANDOM}};
  amplifier_0_2_data_173 = _RAND_1847[7:0];
  _RAND_1848 = {1{`RANDOM}};
  amplifier_0_2_data_174 = _RAND_1848[7:0];
  _RAND_1849 = {1{`RANDOM}};
  amplifier_0_2_data_175 = _RAND_1849[7:0];
  _RAND_1850 = {1{`RANDOM}};
  amplifier_0_2_data_176 = _RAND_1850[7:0];
  _RAND_1851 = {1{`RANDOM}};
  amplifier_0_2_data_177 = _RAND_1851[7:0];
  _RAND_1852 = {1{`RANDOM}};
  amplifier_0_2_data_178 = _RAND_1852[7:0];
  _RAND_1853 = {1{`RANDOM}};
  amplifier_0_2_data_179 = _RAND_1853[7:0];
  _RAND_1854 = {1{`RANDOM}};
  amplifier_0_2_data_180 = _RAND_1854[7:0];
  _RAND_1855 = {1{`RANDOM}};
  amplifier_0_2_data_181 = _RAND_1855[7:0];
  _RAND_1856 = {1{`RANDOM}};
  amplifier_0_2_data_182 = _RAND_1856[7:0];
  _RAND_1857 = {1{`RANDOM}};
  amplifier_0_2_data_183 = _RAND_1857[7:0];
  _RAND_1858 = {1{`RANDOM}};
  amplifier_0_2_data_184 = _RAND_1858[7:0];
  _RAND_1859 = {1{`RANDOM}};
  amplifier_0_2_data_185 = _RAND_1859[7:0];
  _RAND_1860 = {1{`RANDOM}};
  amplifier_0_2_data_186 = _RAND_1860[7:0];
  _RAND_1861 = {1{`RANDOM}};
  amplifier_0_2_data_187 = _RAND_1861[7:0];
  _RAND_1862 = {1{`RANDOM}};
  amplifier_0_2_data_188 = _RAND_1862[7:0];
  _RAND_1863 = {1{`RANDOM}};
  amplifier_0_2_data_189 = _RAND_1863[7:0];
  _RAND_1864 = {1{`RANDOM}};
  amplifier_0_2_data_190 = _RAND_1864[7:0];
  _RAND_1865 = {1{`RANDOM}};
  amplifier_0_2_data_191 = _RAND_1865[7:0];
  _RAND_1866 = {1{`RANDOM}};
  amplifier_0_2_data_192 = _RAND_1866[7:0];
  _RAND_1867 = {1{`RANDOM}};
  amplifier_0_2_data_193 = _RAND_1867[7:0];
  _RAND_1868 = {1{`RANDOM}};
  amplifier_0_2_data_194 = _RAND_1868[7:0];
  _RAND_1869 = {1{`RANDOM}};
  amplifier_0_2_data_195 = _RAND_1869[7:0];
  _RAND_1870 = {1{`RANDOM}};
  amplifier_0_2_data_196 = _RAND_1870[7:0];
  _RAND_1871 = {1{`RANDOM}};
  amplifier_0_2_data_197 = _RAND_1871[7:0];
  _RAND_1872 = {1{`RANDOM}};
  amplifier_0_2_data_198 = _RAND_1872[7:0];
  _RAND_1873 = {1{`RANDOM}};
  amplifier_0_2_data_199 = _RAND_1873[7:0];
  _RAND_1874 = {1{`RANDOM}};
  amplifier_0_2_data_200 = _RAND_1874[7:0];
  _RAND_1875 = {1{`RANDOM}};
  amplifier_0_2_data_201 = _RAND_1875[7:0];
  _RAND_1876 = {1{`RANDOM}};
  amplifier_0_2_data_202 = _RAND_1876[7:0];
  _RAND_1877 = {1{`RANDOM}};
  amplifier_0_2_data_203 = _RAND_1877[7:0];
  _RAND_1878 = {1{`RANDOM}};
  amplifier_0_2_data_204 = _RAND_1878[7:0];
  _RAND_1879 = {1{`RANDOM}};
  amplifier_0_2_data_205 = _RAND_1879[7:0];
  _RAND_1880 = {1{`RANDOM}};
  amplifier_0_2_data_206 = _RAND_1880[7:0];
  _RAND_1881 = {1{`RANDOM}};
  amplifier_0_2_data_207 = _RAND_1881[7:0];
  _RAND_1882 = {1{`RANDOM}};
  amplifier_0_2_data_208 = _RAND_1882[7:0];
  _RAND_1883 = {1{`RANDOM}};
  amplifier_0_2_data_209 = _RAND_1883[7:0];
  _RAND_1884 = {1{`RANDOM}};
  amplifier_0_2_data_210 = _RAND_1884[7:0];
  _RAND_1885 = {1{`RANDOM}};
  amplifier_0_2_data_211 = _RAND_1885[7:0];
  _RAND_1886 = {1{`RANDOM}};
  amplifier_0_2_data_212 = _RAND_1886[7:0];
  _RAND_1887 = {1{`RANDOM}};
  amplifier_0_2_data_213 = _RAND_1887[7:0];
  _RAND_1888 = {1{`RANDOM}};
  amplifier_0_2_data_214 = _RAND_1888[7:0];
  _RAND_1889 = {1{`RANDOM}};
  amplifier_0_2_data_215 = _RAND_1889[7:0];
  _RAND_1890 = {1{`RANDOM}};
  amplifier_0_2_data_216 = _RAND_1890[7:0];
  _RAND_1891 = {1{`RANDOM}};
  amplifier_0_2_data_217 = _RAND_1891[7:0];
  _RAND_1892 = {1{`RANDOM}};
  amplifier_0_2_data_218 = _RAND_1892[7:0];
  _RAND_1893 = {1{`RANDOM}};
  amplifier_0_2_data_219 = _RAND_1893[7:0];
  _RAND_1894 = {1{`RANDOM}};
  amplifier_0_2_data_220 = _RAND_1894[7:0];
  _RAND_1895 = {1{`RANDOM}};
  amplifier_0_2_data_221 = _RAND_1895[7:0];
  _RAND_1896 = {1{`RANDOM}};
  amplifier_0_2_data_222 = _RAND_1896[7:0];
  _RAND_1897 = {1{`RANDOM}};
  amplifier_0_2_data_223 = _RAND_1897[7:0];
  _RAND_1898 = {1{`RANDOM}};
  amplifier_0_2_data_224 = _RAND_1898[7:0];
  _RAND_1899 = {1{`RANDOM}};
  amplifier_0_2_data_225 = _RAND_1899[7:0];
  _RAND_1900 = {1{`RANDOM}};
  amplifier_0_2_data_226 = _RAND_1900[7:0];
  _RAND_1901 = {1{`RANDOM}};
  amplifier_0_2_data_227 = _RAND_1901[7:0];
  _RAND_1902 = {1{`RANDOM}};
  amplifier_0_2_data_228 = _RAND_1902[7:0];
  _RAND_1903 = {1{`RANDOM}};
  amplifier_0_2_data_229 = _RAND_1903[7:0];
  _RAND_1904 = {1{`RANDOM}};
  amplifier_0_2_data_230 = _RAND_1904[7:0];
  _RAND_1905 = {1{`RANDOM}};
  amplifier_0_2_data_231 = _RAND_1905[7:0];
  _RAND_1906 = {1{`RANDOM}};
  amplifier_0_2_data_232 = _RAND_1906[7:0];
  _RAND_1907 = {1{`RANDOM}};
  amplifier_0_2_data_233 = _RAND_1907[7:0];
  _RAND_1908 = {1{`RANDOM}};
  amplifier_0_2_data_234 = _RAND_1908[7:0];
  _RAND_1909 = {1{`RANDOM}};
  amplifier_0_2_data_235 = _RAND_1909[7:0];
  _RAND_1910 = {1{`RANDOM}};
  amplifier_0_2_data_236 = _RAND_1910[7:0];
  _RAND_1911 = {1{`RANDOM}};
  amplifier_0_2_data_237 = _RAND_1911[7:0];
  _RAND_1912 = {1{`RANDOM}};
  amplifier_0_2_data_238 = _RAND_1912[7:0];
  _RAND_1913 = {1{`RANDOM}};
  amplifier_0_2_data_239 = _RAND_1913[7:0];
  _RAND_1914 = {1{`RANDOM}};
  amplifier_0_2_data_240 = _RAND_1914[7:0];
  _RAND_1915 = {1{`RANDOM}};
  amplifier_0_2_data_241 = _RAND_1915[7:0];
  _RAND_1916 = {1{`RANDOM}};
  amplifier_0_2_data_242 = _RAND_1916[7:0];
  _RAND_1917 = {1{`RANDOM}};
  amplifier_0_2_data_243 = _RAND_1917[7:0];
  _RAND_1918 = {1{`RANDOM}};
  amplifier_0_2_data_244 = _RAND_1918[7:0];
  _RAND_1919 = {1{`RANDOM}};
  amplifier_0_2_data_245 = _RAND_1919[7:0];
  _RAND_1920 = {1{`RANDOM}};
  amplifier_0_2_data_246 = _RAND_1920[7:0];
  _RAND_1921 = {1{`RANDOM}};
  amplifier_0_2_data_247 = _RAND_1921[7:0];
  _RAND_1922 = {1{`RANDOM}};
  amplifier_0_2_data_248 = _RAND_1922[7:0];
  _RAND_1923 = {1{`RANDOM}};
  amplifier_0_2_data_249 = _RAND_1923[7:0];
  _RAND_1924 = {1{`RANDOM}};
  amplifier_0_2_data_250 = _RAND_1924[7:0];
  _RAND_1925 = {1{`RANDOM}};
  amplifier_0_2_data_251 = _RAND_1925[7:0];
  _RAND_1926 = {1{`RANDOM}};
  amplifier_0_2_data_252 = _RAND_1926[7:0];
  _RAND_1927 = {1{`RANDOM}};
  amplifier_0_2_data_253 = _RAND_1927[7:0];
  _RAND_1928 = {1{`RANDOM}};
  amplifier_0_2_data_254 = _RAND_1928[7:0];
  _RAND_1929 = {1{`RANDOM}};
  amplifier_0_2_data_255 = _RAND_1929[7:0];
  _RAND_1930 = {1{`RANDOM}};
  amplifier_0_2_header_0 = _RAND_1930[15:0];
  _RAND_1931 = {1{`RANDOM}};
  amplifier_0_2_header_1 = _RAND_1931[15:0];
  _RAND_1932 = {1{`RANDOM}};
  amplifier_0_2_header_2 = _RAND_1932[15:0];
  _RAND_1933 = {1{`RANDOM}};
  amplifier_0_2_header_3 = _RAND_1933[15:0];
  _RAND_1934 = {1{`RANDOM}};
  amplifier_0_2_header_4 = _RAND_1934[15:0];
  _RAND_1935 = {1{`RANDOM}};
  amplifier_0_2_header_5 = _RAND_1935[15:0];
  _RAND_1936 = {1{`RANDOM}};
  amplifier_0_2_header_6 = _RAND_1936[15:0];
  _RAND_1937 = {1{`RANDOM}};
  amplifier_0_2_header_7 = _RAND_1937[15:0];
  _RAND_1938 = {1{`RANDOM}};
  amplifier_0_2_header_8 = _RAND_1938[15:0];
  _RAND_1939 = {1{`RANDOM}};
  amplifier_0_2_header_9 = _RAND_1939[15:0];
  _RAND_1940 = {1{`RANDOM}};
  amplifier_0_2_header_10 = _RAND_1940[15:0];
  _RAND_1941 = {1{`RANDOM}};
  amplifier_0_2_header_11 = _RAND_1941[15:0];
  _RAND_1942 = {1{`RANDOM}};
  amplifier_0_2_header_12 = _RAND_1942[15:0];
  _RAND_1943 = {1{`RANDOM}};
  amplifier_0_2_header_13 = _RAND_1943[15:0];
  _RAND_1944 = {1{`RANDOM}};
  amplifier_0_2_header_14 = _RAND_1944[15:0];
  _RAND_1945 = {1{`RANDOM}};
  amplifier_0_2_header_15 = _RAND_1945[15:0];
  _RAND_1946 = {1{`RANDOM}};
  amplifier_0_2_parse_current_state = _RAND_1946[7:0];
  _RAND_1947 = {1{`RANDOM}};
  amplifier_0_2_parse_current_offset = _RAND_1947[7:0];
  _RAND_1948 = {1{`RANDOM}};
  amplifier_0_2_parse_transition_field = _RAND_1948[15:0];
  _RAND_1949 = {1{`RANDOM}};
  amplifier_0_2_next_processor_id = _RAND_1949[1:0];
  _RAND_1950 = {1{`RANDOM}};
  amplifier_0_2_next_config_id = _RAND_1950[0:0];
  _RAND_1951 = {1{`RANDOM}};
  amplifier_0_2_is_valid_processor = _RAND_1951[0:0];
  _RAND_1952 = {1{`RANDOM}};
  amplifier_0_3_data_0 = _RAND_1952[7:0];
  _RAND_1953 = {1{`RANDOM}};
  amplifier_0_3_data_1 = _RAND_1953[7:0];
  _RAND_1954 = {1{`RANDOM}};
  amplifier_0_3_data_2 = _RAND_1954[7:0];
  _RAND_1955 = {1{`RANDOM}};
  amplifier_0_3_data_3 = _RAND_1955[7:0];
  _RAND_1956 = {1{`RANDOM}};
  amplifier_0_3_data_4 = _RAND_1956[7:0];
  _RAND_1957 = {1{`RANDOM}};
  amplifier_0_3_data_5 = _RAND_1957[7:0];
  _RAND_1958 = {1{`RANDOM}};
  amplifier_0_3_data_6 = _RAND_1958[7:0];
  _RAND_1959 = {1{`RANDOM}};
  amplifier_0_3_data_7 = _RAND_1959[7:0];
  _RAND_1960 = {1{`RANDOM}};
  amplifier_0_3_data_8 = _RAND_1960[7:0];
  _RAND_1961 = {1{`RANDOM}};
  amplifier_0_3_data_9 = _RAND_1961[7:0];
  _RAND_1962 = {1{`RANDOM}};
  amplifier_0_3_data_10 = _RAND_1962[7:0];
  _RAND_1963 = {1{`RANDOM}};
  amplifier_0_3_data_11 = _RAND_1963[7:0];
  _RAND_1964 = {1{`RANDOM}};
  amplifier_0_3_data_12 = _RAND_1964[7:0];
  _RAND_1965 = {1{`RANDOM}};
  amplifier_0_3_data_13 = _RAND_1965[7:0];
  _RAND_1966 = {1{`RANDOM}};
  amplifier_0_3_data_14 = _RAND_1966[7:0];
  _RAND_1967 = {1{`RANDOM}};
  amplifier_0_3_data_15 = _RAND_1967[7:0];
  _RAND_1968 = {1{`RANDOM}};
  amplifier_0_3_data_16 = _RAND_1968[7:0];
  _RAND_1969 = {1{`RANDOM}};
  amplifier_0_3_data_17 = _RAND_1969[7:0];
  _RAND_1970 = {1{`RANDOM}};
  amplifier_0_3_data_18 = _RAND_1970[7:0];
  _RAND_1971 = {1{`RANDOM}};
  amplifier_0_3_data_19 = _RAND_1971[7:0];
  _RAND_1972 = {1{`RANDOM}};
  amplifier_0_3_data_20 = _RAND_1972[7:0];
  _RAND_1973 = {1{`RANDOM}};
  amplifier_0_3_data_21 = _RAND_1973[7:0];
  _RAND_1974 = {1{`RANDOM}};
  amplifier_0_3_data_22 = _RAND_1974[7:0];
  _RAND_1975 = {1{`RANDOM}};
  amplifier_0_3_data_23 = _RAND_1975[7:0];
  _RAND_1976 = {1{`RANDOM}};
  amplifier_0_3_data_24 = _RAND_1976[7:0];
  _RAND_1977 = {1{`RANDOM}};
  amplifier_0_3_data_25 = _RAND_1977[7:0];
  _RAND_1978 = {1{`RANDOM}};
  amplifier_0_3_data_26 = _RAND_1978[7:0];
  _RAND_1979 = {1{`RANDOM}};
  amplifier_0_3_data_27 = _RAND_1979[7:0];
  _RAND_1980 = {1{`RANDOM}};
  amplifier_0_3_data_28 = _RAND_1980[7:0];
  _RAND_1981 = {1{`RANDOM}};
  amplifier_0_3_data_29 = _RAND_1981[7:0];
  _RAND_1982 = {1{`RANDOM}};
  amplifier_0_3_data_30 = _RAND_1982[7:0];
  _RAND_1983 = {1{`RANDOM}};
  amplifier_0_3_data_31 = _RAND_1983[7:0];
  _RAND_1984 = {1{`RANDOM}};
  amplifier_0_3_data_32 = _RAND_1984[7:0];
  _RAND_1985 = {1{`RANDOM}};
  amplifier_0_3_data_33 = _RAND_1985[7:0];
  _RAND_1986 = {1{`RANDOM}};
  amplifier_0_3_data_34 = _RAND_1986[7:0];
  _RAND_1987 = {1{`RANDOM}};
  amplifier_0_3_data_35 = _RAND_1987[7:0];
  _RAND_1988 = {1{`RANDOM}};
  amplifier_0_3_data_36 = _RAND_1988[7:0];
  _RAND_1989 = {1{`RANDOM}};
  amplifier_0_3_data_37 = _RAND_1989[7:0];
  _RAND_1990 = {1{`RANDOM}};
  amplifier_0_3_data_38 = _RAND_1990[7:0];
  _RAND_1991 = {1{`RANDOM}};
  amplifier_0_3_data_39 = _RAND_1991[7:0];
  _RAND_1992 = {1{`RANDOM}};
  amplifier_0_3_data_40 = _RAND_1992[7:0];
  _RAND_1993 = {1{`RANDOM}};
  amplifier_0_3_data_41 = _RAND_1993[7:0];
  _RAND_1994 = {1{`RANDOM}};
  amplifier_0_3_data_42 = _RAND_1994[7:0];
  _RAND_1995 = {1{`RANDOM}};
  amplifier_0_3_data_43 = _RAND_1995[7:0];
  _RAND_1996 = {1{`RANDOM}};
  amplifier_0_3_data_44 = _RAND_1996[7:0];
  _RAND_1997 = {1{`RANDOM}};
  amplifier_0_3_data_45 = _RAND_1997[7:0];
  _RAND_1998 = {1{`RANDOM}};
  amplifier_0_3_data_46 = _RAND_1998[7:0];
  _RAND_1999 = {1{`RANDOM}};
  amplifier_0_3_data_47 = _RAND_1999[7:0];
  _RAND_2000 = {1{`RANDOM}};
  amplifier_0_3_data_48 = _RAND_2000[7:0];
  _RAND_2001 = {1{`RANDOM}};
  amplifier_0_3_data_49 = _RAND_2001[7:0];
  _RAND_2002 = {1{`RANDOM}};
  amplifier_0_3_data_50 = _RAND_2002[7:0];
  _RAND_2003 = {1{`RANDOM}};
  amplifier_0_3_data_51 = _RAND_2003[7:0];
  _RAND_2004 = {1{`RANDOM}};
  amplifier_0_3_data_52 = _RAND_2004[7:0];
  _RAND_2005 = {1{`RANDOM}};
  amplifier_0_3_data_53 = _RAND_2005[7:0];
  _RAND_2006 = {1{`RANDOM}};
  amplifier_0_3_data_54 = _RAND_2006[7:0];
  _RAND_2007 = {1{`RANDOM}};
  amplifier_0_3_data_55 = _RAND_2007[7:0];
  _RAND_2008 = {1{`RANDOM}};
  amplifier_0_3_data_56 = _RAND_2008[7:0];
  _RAND_2009 = {1{`RANDOM}};
  amplifier_0_3_data_57 = _RAND_2009[7:0];
  _RAND_2010 = {1{`RANDOM}};
  amplifier_0_3_data_58 = _RAND_2010[7:0];
  _RAND_2011 = {1{`RANDOM}};
  amplifier_0_3_data_59 = _RAND_2011[7:0];
  _RAND_2012 = {1{`RANDOM}};
  amplifier_0_3_data_60 = _RAND_2012[7:0];
  _RAND_2013 = {1{`RANDOM}};
  amplifier_0_3_data_61 = _RAND_2013[7:0];
  _RAND_2014 = {1{`RANDOM}};
  amplifier_0_3_data_62 = _RAND_2014[7:0];
  _RAND_2015 = {1{`RANDOM}};
  amplifier_0_3_data_63 = _RAND_2015[7:0];
  _RAND_2016 = {1{`RANDOM}};
  amplifier_0_3_data_64 = _RAND_2016[7:0];
  _RAND_2017 = {1{`RANDOM}};
  amplifier_0_3_data_65 = _RAND_2017[7:0];
  _RAND_2018 = {1{`RANDOM}};
  amplifier_0_3_data_66 = _RAND_2018[7:0];
  _RAND_2019 = {1{`RANDOM}};
  amplifier_0_3_data_67 = _RAND_2019[7:0];
  _RAND_2020 = {1{`RANDOM}};
  amplifier_0_3_data_68 = _RAND_2020[7:0];
  _RAND_2021 = {1{`RANDOM}};
  amplifier_0_3_data_69 = _RAND_2021[7:0];
  _RAND_2022 = {1{`RANDOM}};
  amplifier_0_3_data_70 = _RAND_2022[7:0];
  _RAND_2023 = {1{`RANDOM}};
  amplifier_0_3_data_71 = _RAND_2023[7:0];
  _RAND_2024 = {1{`RANDOM}};
  amplifier_0_3_data_72 = _RAND_2024[7:0];
  _RAND_2025 = {1{`RANDOM}};
  amplifier_0_3_data_73 = _RAND_2025[7:0];
  _RAND_2026 = {1{`RANDOM}};
  amplifier_0_3_data_74 = _RAND_2026[7:0];
  _RAND_2027 = {1{`RANDOM}};
  amplifier_0_3_data_75 = _RAND_2027[7:0];
  _RAND_2028 = {1{`RANDOM}};
  amplifier_0_3_data_76 = _RAND_2028[7:0];
  _RAND_2029 = {1{`RANDOM}};
  amplifier_0_3_data_77 = _RAND_2029[7:0];
  _RAND_2030 = {1{`RANDOM}};
  amplifier_0_3_data_78 = _RAND_2030[7:0];
  _RAND_2031 = {1{`RANDOM}};
  amplifier_0_3_data_79 = _RAND_2031[7:0];
  _RAND_2032 = {1{`RANDOM}};
  amplifier_0_3_data_80 = _RAND_2032[7:0];
  _RAND_2033 = {1{`RANDOM}};
  amplifier_0_3_data_81 = _RAND_2033[7:0];
  _RAND_2034 = {1{`RANDOM}};
  amplifier_0_3_data_82 = _RAND_2034[7:0];
  _RAND_2035 = {1{`RANDOM}};
  amplifier_0_3_data_83 = _RAND_2035[7:0];
  _RAND_2036 = {1{`RANDOM}};
  amplifier_0_3_data_84 = _RAND_2036[7:0];
  _RAND_2037 = {1{`RANDOM}};
  amplifier_0_3_data_85 = _RAND_2037[7:0];
  _RAND_2038 = {1{`RANDOM}};
  amplifier_0_3_data_86 = _RAND_2038[7:0];
  _RAND_2039 = {1{`RANDOM}};
  amplifier_0_3_data_87 = _RAND_2039[7:0];
  _RAND_2040 = {1{`RANDOM}};
  amplifier_0_3_data_88 = _RAND_2040[7:0];
  _RAND_2041 = {1{`RANDOM}};
  amplifier_0_3_data_89 = _RAND_2041[7:0];
  _RAND_2042 = {1{`RANDOM}};
  amplifier_0_3_data_90 = _RAND_2042[7:0];
  _RAND_2043 = {1{`RANDOM}};
  amplifier_0_3_data_91 = _RAND_2043[7:0];
  _RAND_2044 = {1{`RANDOM}};
  amplifier_0_3_data_92 = _RAND_2044[7:0];
  _RAND_2045 = {1{`RANDOM}};
  amplifier_0_3_data_93 = _RAND_2045[7:0];
  _RAND_2046 = {1{`RANDOM}};
  amplifier_0_3_data_94 = _RAND_2046[7:0];
  _RAND_2047 = {1{`RANDOM}};
  amplifier_0_3_data_95 = _RAND_2047[7:0];
  _RAND_2048 = {1{`RANDOM}};
  amplifier_0_3_data_96 = _RAND_2048[7:0];
  _RAND_2049 = {1{`RANDOM}};
  amplifier_0_3_data_97 = _RAND_2049[7:0];
  _RAND_2050 = {1{`RANDOM}};
  amplifier_0_3_data_98 = _RAND_2050[7:0];
  _RAND_2051 = {1{`RANDOM}};
  amplifier_0_3_data_99 = _RAND_2051[7:0];
  _RAND_2052 = {1{`RANDOM}};
  amplifier_0_3_data_100 = _RAND_2052[7:0];
  _RAND_2053 = {1{`RANDOM}};
  amplifier_0_3_data_101 = _RAND_2053[7:0];
  _RAND_2054 = {1{`RANDOM}};
  amplifier_0_3_data_102 = _RAND_2054[7:0];
  _RAND_2055 = {1{`RANDOM}};
  amplifier_0_3_data_103 = _RAND_2055[7:0];
  _RAND_2056 = {1{`RANDOM}};
  amplifier_0_3_data_104 = _RAND_2056[7:0];
  _RAND_2057 = {1{`RANDOM}};
  amplifier_0_3_data_105 = _RAND_2057[7:0];
  _RAND_2058 = {1{`RANDOM}};
  amplifier_0_3_data_106 = _RAND_2058[7:0];
  _RAND_2059 = {1{`RANDOM}};
  amplifier_0_3_data_107 = _RAND_2059[7:0];
  _RAND_2060 = {1{`RANDOM}};
  amplifier_0_3_data_108 = _RAND_2060[7:0];
  _RAND_2061 = {1{`RANDOM}};
  amplifier_0_3_data_109 = _RAND_2061[7:0];
  _RAND_2062 = {1{`RANDOM}};
  amplifier_0_3_data_110 = _RAND_2062[7:0];
  _RAND_2063 = {1{`RANDOM}};
  amplifier_0_3_data_111 = _RAND_2063[7:0];
  _RAND_2064 = {1{`RANDOM}};
  amplifier_0_3_data_112 = _RAND_2064[7:0];
  _RAND_2065 = {1{`RANDOM}};
  amplifier_0_3_data_113 = _RAND_2065[7:0];
  _RAND_2066 = {1{`RANDOM}};
  amplifier_0_3_data_114 = _RAND_2066[7:0];
  _RAND_2067 = {1{`RANDOM}};
  amplifier_0_3_data_115 = _RAND_2067[7:0];
  _RAND_2068 = {1{`RANDOM}};
  amplifier_0_3_data_116 = _RAND_2068[7:0];
  _RAND_2069 = {1{`RANDOM}};
  amplifier_0_3_data_117 = _RAND_2069[7:0];
  _RAND_2070 = {1{`RANDOM}};
  amplifier_0_3_data_118 = _RAND_2070[7:0];
  _RAND_2071 = {1{`RANDOM}};
  amplifier_0_3_data_119 = _RAND_2071[7:0];
  _RAND_2072 = {1{`RANDOM}};
  amplifier_0_3_data_120 = _RAND_2072[7:0];
  _RAND_2073 = {1{`RANDOM}};
  amplifier_0_3_data_121 = _RAND_2073[7:0];
  _RAND_2074 = {1{`RANDOM}};
  amplifier_0_3_data_122 = _RAND_2074[7:0];
  _RAND_2075 = {1{`RANDOM}};
  amplifier_0_3_data_123 = _RAND_2075[7:0];
  _RAND_2076 = {1{`RANDOM}};
  amplifier_0_3_data_124 = _RAND_2076[7:0];
  _RAND_2077 = {1{`RANDOM}};
  amplifier_0_3_data_125 = _RAND_2077[7:0];
  _RAND_2078 = {1{`RANDOM}};
  amplifier_0_3_data_126 = _RAND_2078[7:0];
  _RAND_2079 = {1{`RANDOM}};
  amplifier_0_3_data_127 = _RAND_2079[7:0];
  _RAND_2080 = {1{`RANDOM}};
  amplifier_0_3_data_128 = _RAND_2080[7:0];
  _RAND_2081 = {1{`RANDOM}};
  amplifier_0_3_data_129 = _RAND_2081[7:0];
  _RAND_2082 = {1{`RANDOM}};
  amplifier_0_3_data_130 = _RAND_2082[7:0];
  _RAND_2083 = {1{`RANDOM}};
  amplifier_0_3_data_131 = _RAND_2083[7:0];
  _RAND_2084 = {1{`RANDOM}};
  amplifier_0_3_data_132 = _RAND_2084[7:0];
  _RAND_2085 = {1{`RANDOM}};
  amplifier_0_3_data_133 = _RAND_2085[7:0];
  _RAND_2086 = {1{`RANDOM}};
  amplifier_0_3_data_134 = _RAND_2086[7:0];
  _RAND_2087 = {1{`RANDOM}};
  amplifier_0_3_data_135 = _RAND_2087[7:0];
  _RAND_2088 = {1{`RANDOM}};
  amplifier_0_3_data_136 = _RAND_2088[7:0];
  _RAND_2089 = {1{`RANDOM}};
  amplifier_0_3_data_137 = _RAND_2089[7:0];
  _RAND_2090 = {1{`RANDOM}};
  amplifier_0_3_data_138 = _RAND_2090[7:0];
  _RAND_2091 = {1{`RANDOM}};
  amplifier_0_3_data_139 = _RAND_2091[7:0];
  _RAND_2092 = {1{`RANDOM}};
  amplifier_0_3_data_140 = _RAND_2092[7:0];
  _RAND_2093 = {1{`RANDOM}};
  amplifier_0_3_data_141 = _RAND_2093[7:0];
  _RAND_2094 = {1{`RANDOM}};
  amplifier_0_3_data_142 = _RAND_2094[7:0];
  _RAND_2095 = {1{`RANDOM}};
  amplifier_0_3_data_143 = _RAND_2095[7:0];
  _RAND_2096 = {1{`RANDOM}};
  amplifier_0_3_data_144 = _RAND_2096[7:0];
  _RAND_2097 = {1{`RANDOM}};
  amplifier_0_3_data_145 = _RAND_2097[7:0];
  _RAND_2098 = {1{`RANDOM}};
  amplifier_0_3_data_146 = _RAND_2098[7:0];
  _RAND_2099 = {1{`RANDOM}};
  amplifier_0_3_data_147 = _RAND_2099[7:0];
  _RAND_2100 = {1{`RANDOM}};
  amplifier_0_3_data_148 = _RAND_2100[7:0];
  _RAND_2101 = {1{`RANDOM}};
  amplifier_0_3_data_149 = _RAND_2101[7:0];
  _RAND_2102 = {1{`RANDOM}};
  amplifier_0_3_data_150 = _RAND_2102[7:0];
  _RAND_2103 = {1{`RANDOM}};
  amplifier_0_3_data_151 = _RAND_2103[7:0];
  _RAND_2104 = {1{`RANDOM}};
  amplifier_0_3_data_152 = _RAND_2104[7:0];
  _RAND_2105 = {1{`RANDOM}};
  amplifier_0_3_data_153 = _RAND_2105[7:0];
  _RAND_2106 = {1{`RANDOM}};
  amplifier_0_3_data_154 = _RAND_2106[7:0];
  _RAND_2107 = {1{`RANDOM}};
  amplifier_0_3_data_155 = _RAND_2107[7:0];
  _RAND_2108 = {1{`RANDOM}};
  amplifier_0_3_data_156 = _RAND_2108[7:0];
  _RAND_2109 = {1{`RANDOM}};
  amplifier_0_3_data_157 = _RAND_2109[7:0];
  _RAND_2110 = {1{`RANDOM}};
  amplifier_0_3_data_158 = _RAND_2110[7:0];
  _RAND_2111 = {1{`RANDOM}};
  amplifier_0_3_data_159 = _RAND_2111[7:0];
  _RAND_2112 = {1{`RANDOM}};
  amplifier_0_3_data_160 = _RAND_2112[7:0];
  _RAND_2113 = {1{`RANDOM}};
  amplifier_0_3_data_161 = _RAND_2113[7:0];
  _RAND_2114 = {1{`RANDOM}};
  amplifier_0_3_data_162 = _RAND_2114[7:0];
  _RAND_2115 = {1{`RANDOM}};
  amplifier_0_3_data_163 = _RAND_2115[7:0];
  _RAND_2116 = {1{`RANDOM}};
  amplifier_0_3_data_164 = _RAND_2116[7:0];
  _RAND_2117 = {1{`RANDOM}};
  amplifier_0_3_data_165 = _RAND_2117[7:0];
  _RAND_2118 = {1{`RANDOM}};
  amplifier_0_3_data_166 = _RAND_2118[7:0];
  _RAND_2119 = {1{`RANDOM}};
  amplifier_0_3_data_167 = _RAND_2119[7:0];
  _RAND_2120 = {1{`RANDOM}};
  amplifier_0_3_data_168 = _RAND_2120[7:0];
  _RAND_2121 = {1{`RANDOM}};
  amplifier_0_3_data_169 = _RAND_2121[7:0];
  _RAND_2122 = {1{`RANDOM}};
  amplifier_0_3_data_170 = _RAND_2122[7:0];
  _RAND_2123 = {1{`RANDOM}};
  amplifier_0_3_data_171 = _RAND_2123[7:0];
  _RAND_2124 = {1{`RANDOM}};
  amplifier_0_3_data_172 = _RAND_2124[7:0];
  _RAND_2125 = {1{`RANDOM}};
  amplifier_0_3_data_173 = _RAND_2125[7:0];
  _RAND_2126 = {1{`RANDOM}};
  amplifier_0_3_data_174 = _RAND_2126[7:0];
  _RAND_2127 = {1{`RANDOM}};
  amplifier_0_3_data_175 = _RAND_2127[7:0];
  _RAND_2128 = {1{`RANDOM}};
  amplifier_0_3_data_176 = _RAND_2128[7:0];
  _RAND_2129 = {1{`RANDOM}};
  amplifier_0_3_data_177 = _RAND_2129[7:0];
  _RAND_2130 = {1{`RANDOM}};
  amplifier_0_3_data_178 = _RAND_2130[7:0];
  _RAND_2131 = {1{`RANDOM}};
  amplifier_0_3_data_179 = _RAND_2131[7:0];
  _RAND_2132 = {1{`RANDOM}};
  amplifier_0_3_data_180 = _RAND_2132[7:0];
  _RAND_2133 = {1{`RANDOM}};
  amplifier_0_3_data_181 = _RAND_2133[7:0];
  _RAND_2134 = {1{`RANDOM}};
  amplifier_0_3_data_182 = _RAND_2134[7:0];
  _RAND_2135 = {1{`RANDOM}};
  amplifier_0_3_data_183 = _RAND_2135[7:0];
  _RAND_2136 = {1{`RANDOM}};
  amplifier_0_3_data_184 = _RAND_2136[7:0];
  _RAND_2137 = {1{`RANDOM}};
  amplifier_0_3_data_185 = _RAND_2137[7:0];
  _RAND_2138 = {1{`RANDOM}};
  amplifier_0_3_data_186 = _RAND_2138[7:0];
  _RAND_2139 = {1{`RANDOM}};
  amplifier_0_3_data_187 = _RAND_2139[7:0];
  _RAND_2140 = {1{`RANDOM}};
  amplifier_0_3_data_188 = _RAND_2140[7:0];
  _RAND_2141 = {1{`RANDOM}};
  amplifier_0_3_data_189 = _RAND_2141[7:0];
  _RAND_2142 = {1{`RANDOM}};
  amplifier_0_3_data_190 = _RAND_2142[7:0];
  _RAND_2143 = {1{`RANDOM}};
  amplifier_0_3_data_191 = _RAND_2143[7:0];
  _RAND_2144 = {1{`RANDOM}};
  amplifier_0_3_data_192 = _RAND_2144[7:0];
  _RAND_2145 = {1{`RANDOM}};
  amplifier_0_3_data_193 = _RAND_2145[7:0];
  _RAND_2146 = {1{`RANDOM}};
  amplifier_0_3_data_194 = _RAND_2146[7:0];
  _RAND_2147 = {1{`RANDOM}};
  amplifier_0_3_data_195 = _RAND_2147[7:0];
  _RAND_2148 = {1{`RANDOM}};
  amplifier_0_3_data_196 = _RAND_2148[7:0];
  _RAND_2149 = {1{`RANDOM}};
  amplifier_0_3_data_197 = _RAND_2149[7:0];
  _RAND_2150 = {1{`RANDOM}};
  amplifier_0_3_data_198 = _RAND_2150[7:0];
  _RAND_2151 = {1{`RANDOM}};
  amplifier_0_3_data_199 = _RAND_2151[7:0];
  _RAND_2152 = {1{`RANDOM}};
  amplifier_0_3_data_200 = _RAND_2152[7:0];
  _RAND_2153 = {1{`RANDOM}};
  amplifier_0_3_data_201 = _RAND_2153[7:0];
  _RAND_2154 = {1{`RANDOM}};
  amplifier_0_3_data_202 = _RAND_2154[7:0];
  _RAND_2155 = {1{`RANDOM}};
  amplifier_0_3_data_203 = _RAND_2155[7:0];
  _RAND_2156 = {1{`RANDOM}};
  amplifier_0_3_data_204 = _RAND_2156[7:0];
  _RAND_2157 = {1{`RANDOM}};
  amplifier_0_3_data_205 = _RAND_2157[7:0];
  _RAND_2158 = {1{`RANDOM}};
  amplifier_0_3_data_206 = _RAND_2158[7:0];
  _RAND_2159 = {1{`RANDOM}};
  amplifier_0_3_data_207 = _RAND_2159[7:0];
  _RAND_2160 = {1{`RANDOM}};
  amplifier_0_3_data_208 = _RAND_2160[7:0];
  _RAND_2161 = {1{`RANDOM}};
  amplifier_0_3_data_209 = _RAND_2161[7:0];
  _RAND_2162 = {1{`RANDOM}};
  amplifier_0_3_data_210 = _RAND_2162[7:0];
  _RAND_2163 = {1{`RANDOM}};
  amplifier_0_3_data_211 = _RAND_2163[7:0];
  _RAND_2164 = {1{`RANDOM}};
  amplifier_0_3_data_212 = _RAND_2164[7:0];
  _RAND_2165 = {1{`RANDOM}};
  amplifier_0_3_data_213 = _RAND_2165[7:0];
  _RAND_2166 = {1{`RANDOM}};
  amplifier_0_3_data_214 = _RAND_2166[7:0];
  _RAND_2167 = {1{`RANDOM}};
  amplifier_0_3_data_215 = _RAND_2167[7:0];
  _RAND_2168 = {1{`RANDOM}};
  amplifier_0_3_data_216 = _RAND_2168[7:0];
  _RAND_2169 = {1{`RANDOM}};
  amplifier_0_3_data_217 = _RAND_2169[7:0];
  _RAND_2170 = {1{`RANDOM}};
  amplifier_0_3_data_218 = _RAND_2170[7:0];
  _RAND_2171 = {1{`RANDOM}};
  amplifier_0_3_data_219 = _RAND_2171[7:0];
  _RAND_2172 = {1{`RANDOM}};
  amplifier_0_3_data_220 = _RAND_2172[7:0];
  _RAND_2173 = {1{`RANDOM}};
  amplifier_0_3_data_221 = _RAND_2173[7:0];
  _RAND_2174 = {1{`RANDOM}};
  amplifier_0_3_data_222 = _RAND_2174[7:0];
  _RAND_2175 = {1{`RANDOM}};
  amplifier_0_3_data_223 = _RAND_2175[7:0];
  _RAND_2176 = {1{`RANDOM}};
  amplifier_0_3_data_224 = _RAND_2176[7:0];
  _RAND_2177 = {1{`RANDOM}};
  amplifier_0_3_data_225 = _RAND_2177[7:0];
  _RAND_2178 = {1{`RANDOM}};
  amplifier_0_3_data_226 = _RAND_2178[7:0];
  _RAND_2179 = {1{`RANDOM}};
  amplifier_0_3_data_227 = _RAND_2179[7:0];
  _RAND_2180 = {1{`RANDOM}};
  amplifier_0_3_data_228 = _RAND_2180[7:0];
  _RAND_2181 = {1{`RANDOM}};
  amplifier_0_3_data_229 = _RAND_2181[7:0];
  _RAND_2182 = {1{`RANDOM}};
  amplifier_0_3_data_230 = _RAND_2182[7:0];
  _RAND_2183 = {1{`RANDOM}};
  amplifier_0_3_data_231 = _RAND_2183[7:0];
  _RAND_2184 = {1{`RANDOM}};
  amplifier_0_3_data_232 = _RAND_2184[7:0];
  _RAND_2185 = {1{`RANDOM}};
  amplifier_0_3_data_233 = _RAND_2185[7:0];
  _RAND_2186 = {1{`RANDOM}};
  amplifier_0_3_data_234 = _RAND_2186[7:0];
  _RAND_2187 = {1{`RANDOM}};
  amplifier_0_3_data_235 = _RAND_2187[7:0];
  _RAND_2188 = {1{`RANDOM}};
  amplifier_0_3_data_236 = _RAND_2188[7:0];
  _RAND_2189 = {1{`RANDOM}};
  amplifier_0_3_data_237 = _RAND_2189[7:0];
  _RAND_2190 = {1{`RANDOM}};
  amplifier_0_3_data_238 = _RAND_2190[7:0];
  _RAND_2191 = {1{`RANDOM}};
  amplifier_0_3_data_239 = _RAND_2191[7:0];
  _RAND_2192 = {1{`RANDOM}};
  amplifier_0_3_data_240 = _RAND_2192[7:0];
  _RAND_2193 = {1{`RANDOM}};
  amplifier_0_3_data_241 = _RAND_2193[7:0];
  _RAND_2194 = {1{`RANDOM}};
  amplifier_0_3_data_242 = _RAND_2194[7:0];
  _RAND_2195 = {1{`RANDOM}};
  amplifier_0_3_data_243 = _RAND_2195[7:0];
  _RAND_2196 = {1{`RANDOM}};
  amplifier_0_3_data_244 = _RAND_2196[7:0];
  _RAND_2197 = {1{`RANDOM}};
  amplifier_0_3_data_245 = _RAND_2197[7:0];
  _RAND_2198 = {1{`RANDOM}};
  amplifier_0_3_data_246 = _RAND_2198[7:0];
  _RAND_2199 = {1{`RANDOM}};
  amplifier_0_3_data_247 = _RAND_2199[7:0];
  _RAND_2200 = {1{`RANDOM}};
  amplifier_0_3_data_248 = _RAND_2200[7:0];
  _RAND_2201 = {1{`RANDOM}};
  amplifier_0_3_data_249 = _RAND_2201[7:0];
  _RAND_2202 = {1{`RANDOM}};
  amplifier_0_3_data_250 = _RAND_2202[7:0];
  _RAND_2203 = {1{`RANDOM}};
  amplifier_0_3_data_251 = _RAND_2203[7:0];
  _RAND_2204 = {1{`RANDOM}};
  amplifier_0_3_data_252 = _RAND_2204[7:0];
  _RAND_2205 = {1{`RANDOM}};
  amplifier_0_3_data_253 = _RAND_2205[7:0];
  _RAND_2206 = {1{`RANDOM}};
  amplifier_0_3_data_254 = _RAND_2206[7:0];
  _RAND_2207 = {1{`RANDOM}};
  amplifier_0_3_data_255 = _RAND_2207[7:0];
  _RAND_2208 = {1{`RANDOM}};
  amplifier_0_3_header_0 = _RAND_2208[15:0];
  _RAND_2209 = {1{`RANDOM}};
  amplifier_0_3_header_1 = _RAND_2209[15:0];
  _RAND_2210 = {1{`RANDOM}};
  amplifier_0_3_header_2 = _RAND_2210[15:0];
  _RAND_2211 = {1{`RANDOM}};
  amplifier_0_3_header_3 = _RAND_2211[15:0];
  _RAND_2212 = {1{`RANDOM}};
  amplifier_0_3_header_4 = _RAND_2212[15:0];
  _RAND_2213 = {1{`RANDOM}};
  amplifier_0_3_header_5 = _RAND_2213[15:0];
  _RAND_2214 = {1{`RANDOM}};
  amplifier_0_3_header_6 = _RAND_2214[15:0];
  _RAND_2215 = {1{`RANDOM}};
  amplifier_0_3_header_7 = _RAND_2215[15:0];
  _RAND_2216 = {1{`RANDOM}};
  amplifier_0_3_header_8 = _RAND_2216[15:0];
  _RAND_2217 = {1{`RANDOM}};
  amplifier_0_3_header_9 = _RAND_2217[15:0];
  _RAND_2218 = {1{`RANDOM}};
  amplifier_0_3_header_10 = _RAND_2218[15:0];
  _RAND_2219 = {1{`RANDOM}};
  amplifier_0_3_header_11 = _RAND_2219[15:0];
  _RAND_2220 = {1{`RANDOM}};
  amplifier_0_3_header_12 = _RAND_2220[15:0];
  _RAND_2221 = {1{`RANDOM}};
  amplifier_0_3_header_13 = _RAND_2221[15:0];
  _RAND_2222 = {1{`RANDOM}};
  amplifier_0_3_header_14 = _RAND_2222[15:0];
  _RAND_2223 = {1{`RANDOM}};
  amplifier_0_3_header_15 = _RAND_2223[15:0];
  _RAND_2224 = {1{`RANDOM}};
  amplifier_0_3_parse_current_state = _RAND_2224[7:0];
  _RAND_2225 = {1{`RANDOM}};
  amplifier_0_3_parse_current_offset = _RAND_2225[7:0];
  _RAND_2226 = {1{`RANDOM}};
  amplifier_0_3_parse_transition_field = _RAND_2226[15:0];
  _RAND_2227 = {1{`RANDOM}};
  amplifier_0_3_next_processor_id = _RAND_2227[1:0];
  _RAND_2228 = {1{`RANDOM}};
  amplifier_0_3_next_config_id = _RAND_2228[0:0];
  _RAND_2229 = {1{`RANDOM}};
  amplifier_0_3_is_valid_processor = _RAND_2229[0:0];
  _RAND_2230 = {1{`RANDOM}};
  amplifier_1_0_data_0 = _RAND_2230[7:0];
  _RAND_2231 = {1{`RANDOM}};
  amplifier_1_0_data_1 = _RAND_2231[7:0];
  _RAND_2232 = {1{`RANDOM}};
  amplifier_1_0_data_2 = _RAND_2232[7:0];
  _RAND_2233 = {1{`RANDOM}};
  amplifier_1_0_data_3 = _RAND_2233[7:0];
  _RAND_2234 = {1{`RANDOM}};
  amplifier_1_0_data_4 = _RAND_2234[7:0];
  _RAND_2235 = {1{`RANDOM}};
  amplifier_1_0_data_5 = _RAND_2235[7:0];
  _RAND_2236 = {1{`RANDOM}};
  amplifier_1_0_data_6 = _RAND_2236[7:0];
  _RAND_2237 = {1{`RANDOM}};
  amplifier_1_0_data_7 = _RAND_2237[7:0];
  _RAND_2238 = {1{`RANDOM}};
  amplifier_1_0_data_8 = _RAND_2238[7:0];
  _RAND_2239 = {1{`RANDOM}};
  amplifier_1_0_data_9 = _RAND_2239[7:0];
  _RAND_2240 = {1{`RANDOM}};
  amplifier_1_0_data_10 = _RAND_2240[7:0];
  _RAND_2241 = {1{`RANDOM}};
  amplifier_1_0_data_11 = _RAND_2241[7:0];
  _RAND_2242 = {1{`RANDOM}};
  amplifier_1_0_data_12 = _RAND_2242[7:0];
  _RAND_2243 = {1{`RANDOM}};
  amplifier_1_0_data_13 = _RAND_2243[7:0];
  _RAND_2244 = {1{`RANDOM}};
  amplifier_1_0_data_14 = _RAND_2244[7:0];
  _RAND_2245 = {1{`RANDOM}};
  amplifier_1_0_data_15 = _RAND_2245[7:0];
  _RAND_2246 = {1{`RANDOM}};
  amplifier_1_0_data_16 = _RAND_2246[7:0];
  _RAND_2247 = {1{`RANDOM}};
  amplifier_1_0_data_17 = _RAND_2247[7:0];
  _RAND_2248 = {1{`RANDOM}};
  amplifier_1_0_data_18 = _RAND_2248[7:0];
  _RAND_2249 = {1{`RANDOM}};
  amplifier_1_0_data_19 = _RAND_2249[7:0];
  _RAND_2250 = {1{`RANDOM}};
  amplifier_1_0_data_20 = _RAND_2250[7:0];
  _RAND_2251 = {1{`RANDOM}};
  amplifier_1_0_data_21 = _RAND_2251[7:0];
  _RAND_2252 = {1{`RANDOM}};
  amplifier_1_0_data_22 = _RAND_2252[7:0];
  _RAND_2253 = {1{`RANDOM}};
  amplifier_1_0_data_23 = _RAND_2253[7:0];
  _RAND_2254 = {1{`RANDOM}};
  amplifier_1_0_data_24 = _RAND_2254[7:0];
  _RAND_2255 = {1{`RANDOM}};
  amplifier_1_0_data_25 = _RAND_2255[7:0];
  _RAND_2256 = {1{`RANDOM}};
  amplifier_1_0_data_26 = _RAND_2256[7:0];
  _RAND_2257 = {1{`RANDOM}};
  amplifier_1_0_data_27 = _RAND_2257[7:0];
  _RAND_2258 = {1{`RANDOM}};
  amplifier_1_0_data_28 = _RAND_2258[7:0];
  _RAND_2259 = {1{`RANDOM}};
  amplifier_1_0_data_29 = _RAND_2259[7:0];
  _RAND_2260 = {1{`RANDOM}};
  amplifier_1_0_data_30 = _RAND_2260[7:0];
  _RAND_2261 = {1{`RANDOM}};
  amplifier_1_0_data_31 = _RAND_2261[7:0];
  _RAND_2262 = {1{`RANDOM}};
  amplifier_1_0_data_32 = _RAND_2262[7:0];
  _RAND_2263 = {1{`RANDOM}};
  amplifier_1_0_data_33 = _RAND_2263[7:0];
  _RAND_2264 = {1{`RANDOM}};
  amplifier_1_0_data_34 = _RAND_2264[7:0];
  _RAND_2265 = {1{`RANDOM}};
  amplifier_1_0_data_35 = _RAND_2265[7:0];
  _RAND_2266 = {1{`RANDOM}};
  amplifier_1_0_data_36 = _RAND_2266[7:0];
  _RAND_2267 = {1{`RANDOM}};
  amplifier_1_0_data_37 = _RAND_2267[7:0];
  _RAND_2268 = {1{`RANDOM}};
  amplifier_1_0_data_38 = _RAND_2268[7:0];
  _RAND_2269 = {1{`RANDOM}};
  amplifier_1_0_data_39 = _RAND_2269[7:0];
  _RAND_2270 = {1{`RANDOM}};
  amplifier_1_0_data_40 = _RAND_2270[7:0];
  _RAND_2271 = {1{`RANDOM}};
  amplifier_1_0_data_41 = _RAND_2271[7:0];
  _RAND_2272 = {1{`RANDOM}};
  amplifier_1_0_data_42 = _RAND_2272[7:0];
  _RAND_2273 = {1{`RANDOM}};
  amplifier_1_0_data_43 = _RAND_2273[7:0];
  _RAND_2274 = {1{`RANDOM}};
  amplifier_1_0_data_44 = _RAND_2274[7:0];
  _RAND_2275 = {1{`RANDOM}};
  amplifier_1_0_data_45 = _RAND_2275[7:0];
  _RAND_2276 = {1{`RANDOM}};
  amplifier_1_0_data_46 = _RAND_2276[7:0];
  _RAND_2277 = {1{`RANDOM}};
  amplifier_1_0_data_47 = _RAND_2277[7:0];
  _RAND_2278 = {1{`RANDOM}};
  amplifier_1_0_data_48 = _RAND_2278[7:0];
  _RAND_2279 = {1{`RANDOM}};
  amplifier_1_0_data_49 = _RAND_2279[7:0];
  _RAND_2280 = {1{`RANDOM}};
  amplifier_1_0_data_50 = _RAND_2280[7:0];
  _RAND_2281 = {1{`RANDOM}};
  amplifier_1_0_data_51 = _RAND_2281[7:0];
  _RAND_2282 = {1{`RANDOM}};
  amplifier_1_0_data_52 = _RAND_2282[7:0];
  _RAND_2283 = {1{`RANDOM}};
  amplifier_1_0_data_53 = _RAND_2283[7:0];
  _RAND_2284 = {1{`RANDOM}};
  amplifier_1_0_data_54 = _RAND_2284[7:0];
  _RAND_2285 = {1{`RANDOM}};
  amplifier_1_0_data_55 = _RAND_2285[7:0];
  _RAND_2286 = {1{`RANDOM}};
  amplifier_1_0_data_56 = _RAND_2286[7:0];
  _RAND_2287 = {1{`RANDOM}};
  amplifier_1_0_data_57 = _RAND_2287[7:0];
  _RAND_2288 = {1{`RANDOM}};
  amplifier_1_0_data_58 = _RAND_2288[7:0];
  _RAND_2289 = {1{`RANDOM}};
  amplifier_1_0_data_59 = _RAND_2289[7:0];
  _RAND_2290 = {1{`RANDOM}};
  amplifier_1_0_data_60 = _RAND_2290[7:0];
  _RAND_2291 = {1{`RANDOM}};
  amplifier_1_0_data_61 = _RAND_2291[7:0];
  _RAND_2292 = {1{`RANDOM}};
  amplifier_1_0_data_62 = _RAND_2292[7:0];
  _RAND_2293 = {1{`RANDOM}};
  amplifier_1_0_data_63 = _RAND_2293[7:0];
  _RAND_2294 = {1{`RANDOM}};
  amplifier_1_0_data_64 = _RAND_2294[7:0];
  _RAND_2295 = {1{`RANDOM}};
  amplifier_1_0_data_65 = _RAND_2295[7:0];
  _RAND_2296 = {1{`RANDOM}};
  amplifier_1_0_data_66 = _RAND_2296[7:0];
  _RAND_2297 = {1{`RANDOM}};
  amplifier_1_0_data_67 = _RAND_2297[7:0];
  _RAND_2298 = {1{`RANDOM}};
  amplifier_1_0_data_68 = _RAND_2298[7:0];
  _RAND_2299 = {1{`RANDOM}};
  amplifier_1_0_data_69 = _RAND_2299[7:0];
  _RAND_2300 = {1{`RANDOM}};
  amplifier_1_0_data_70 = _RAND_2300[7:0];
  _RAND_2301 = {1{`RANDOM}};
  amplifier_1_0_data_71 = _RAND_2301[7:0];
  _RAND_2302 = {1{`RANDOM}};
  amplifier_1_0_data_72 = _RAND_2302[7:0];
  _RAND_2303 = {1{`RANDOM}};
  amplifier_1_0_data_73 = _RAND_2303[7:0];
  _RAND_2304 = {1{`RANDOM}};
  amplifier_1_0_data_74 = _RAND_2304[7:0];
  _RAND_2305 = {1{`RANDOM}};
  amplifier_1_0_data_75 = _RAND_2305[7:0];
  _RAND_2306 = {1{`RANDOM}};
  amplifier_1_0_data_76 = _RAND_2306[7:0];
  _RAND_2307 = {1{`RANDOM}};
  amplifier_1_0_data_77 = _RAND_2307[7:0];
  _RAND_2308 = {1{`RANDOM}};
  amplifier_1_0_data_78 = _RAND_2308[7:0];
  _RAND_2309 = {1{`RANDOM}};
  amplifier_1_0_data_79 = _RAND_2309[7:0];
  _RAND_2310 = {1{`RANDOM}};
  amplifier_1_0_data_80 = _RAND_2310[7:0];
  _RAND_2311 = {1{`RANDOM}};
  amplifier_1_0_data_81 = _RAND_2311[7:0];
  _RAND_2312 = {1{`RANDOM}};
  amplifier_1_0_data_82 = _RAND_2312[7:0];
  _RAND_2313 = {1{`RANDOM}};
  amplifier_1_0_data_83 = _RAND_2313[7:0];
  _RAND_2314 = {1{`RANDOM}};
  amplifier_1_0_data_84 = _RAND_2314[7:0];
  _RAND_2315 = {1{`RANDOM}};
  amplifier_1_0_data_85 = _RAND_2315[7:0];
  _RAND_2316 = {1{`RANDOM}};
  amplifier_1_0_data_86 = _RAND_2316[7:0];
  _RAND_2317 = {1{`RANDOM}};
  amplifier_1_0_data_87 = _RAND_2317[7:0];
  _RAND_2318 = {1{`RANDOM}};
  amplifier_1_0_data_88 = _RAND_2318[7:0];
  _RAND_2319 = {1{`RANDOM}};
  amplifier_1_0_data_89 = _RAND_2319[7:0];
  _RAND_2320 = {1{`RANDOM}};
  amplifier_1_0_data_90 = _RAND_2320[7:0];
  _RAND_2321 = {1{`RANDOM}};
  amplifier_1_0_data_91 = _RAND_2321[7:0];
  _RAND_2322 = {1{`RANDOM}};
  amplifier_1_0_data_92 = _RAND_2322[7:0];
  _RAND_2323 = {1{`RANDOM}};
  amplifier_1_0_data_93 = _RAND_2323[7:0];
  _RAND_2324 = {1{`RANDOM}};
  amplifier_1_0_data_94 = _RAND_2324[7:0];
  _RAND_2325 = {1{`RANDOM}};
  amplifier_1_0_data_95 = _RAND_2325[7:0];
  _RAND_2326 = {1{`RANDOM}};
  amplifier_1_0_data_96 = _RAND_2326[7:0];
  _RAND_2327 = {1{`RANDOM}};
  amplifier_1_0_data_97 = _RAND_2327[7:0];
  _RAND_2328 = {1{`RANDOM}};
  amplifier_1_0_data_98 = _RAND_2328[7:0];
  _RAND_2329 = {1{`RANDOM}};
  amplifier_1_0_data_99 = _RAND_2329[7:0];
  _RAND_2330 = {1{`RANDOM}};
  amplifier_1_0_data_100 = _RAND_2330[7:0];
  _RAND_2331 = {1{`RANDOM}};
  amplifier_1_0_data_101 = _RAND_2331[7:0];
  _RAND_2332 = {1{`RANDOM}};
  amplifier_1_0_data_102 = _RAND_2332[7:0];
  _RAND_2333 = {1{`RANDOM}};
  amplifier_1_0_data_103 = _RAND_2333[7:0];
  _RAND_2334 = {1{`RANDOM}};
  amplifier_1_0_data_104 = _RAND_2334[7:0];
  _RAND_2335 = {1{`RANDOM}};
  amplifier_1_0_data_105 = _RAND_2335[7:0];
  _RAND_2336 = {1{`RANDOM}};
  amplifier_1_0_data_106 = _RAND_2336[7:0];
  _RAND_2337 = {1{`RANDOM}};
  amplifier_1_0_data_107 = _RAND_2337[7:0];
  _RAND_2338 = {1{`RANDOM}};
  amplifier_1_0_data_108 = _RAND_2338[7:0];
  _RAND_2339 = {1{`RANDOM}};
  amplifier_1_0_data_109 = _RAND_2339[7:0];
  _RAND_2340 = {1{`RANDOM}};
  amplifier_1_0_data_110 = _RAND_2340[7:0];
  _RAND_2341 = {1{`RANDOM}};
  amplifier_1_0_data_111 = _RAND_2341[7:0];
  _RAND_2342 = {1{`RANDOM}};
  amplifier_1_0_data_112 = _RAND_2342[7:0];
  _RAND_2343 = {1{`RANDOM}};
  amplifier_1_0_data_113 = _RAND_2343[7:0];
  _RAND_2344 = {1{`RANDOM}};
  amplifier_1_0_data_114 = _RAND_2344[7:0];
  _RAND_2345 = {1{`RANDOM}};
  amplifier_1_0_data_115 = _RAND_2345[7:0];
  _RAND_2346 = {1{`RANDOM}};
  amplifier_1_0_data_116 = _RAND_2346[7:0];
  _RAND_2347 = {1{`RANDOM}};
  amplifier_1_0_data_117 = _RAND_2347[7:0];
  _RAND_2348 = {1{`RANDOM}};
  amplifier_1_0_data_118 = _RAND_2348[7:0];
  _RAND_2349 = {1{`RANDOM}};
  amplifier_1_0_data_119 = _RAND_2349[7:0];
  _RAND_2350 = {1{`RANDOM}};
  amplifier_1_0_data_120 = _RAND_2350[7:0];
  _RAND_2351 = {1{`RANDOM}};
  amplifier_1_0_data_121 = _RAND_2351[7:0];
  _RAND_2352 = {1{`RANDOM}};
  amplifier_1_0_data_122 = _RAND_2352[7:0];
  _RAND_2353 = {1{`RANDOM}};
  amplifier_1_0_data_123 = _RAND_2353[7:0];
  _RAND_2354 = {1{`RANDOM}};
  amplifier_1_0_data_124 = _RAND_2354[7:0];
  _RAND_2355 = {1{`RANDOM}};
  amplifier_1_0_data_125 = _RAND_2355[7:0];
  _RAND_2356 = {1{`RANDOM}};
  amplifier_1_0_data_126 = _RAND_2356[7:0];
  _RAND_2357 = {1{`RANDOM}};
  amplifier_1_0_data_127 = _RAND_2357[7:0];
  _RAND_2358 = {1{`RANDOM}};
  amplifier_1_0_data_128 = _RAND_2358[7:0];
  _RAND_2359 = {1{`RANDOM}};
  amplifier_1_0_data_129 = _RAND_2359[7:0];
  _RAND_2360 = {1{`RANDOM}};
  amplifier_1_0_data_130 = _RAND_2360[7:0];
  _RAND_2361 = {1{`RANDOM}};
  amplifier_1_0_data_131 = _RAND_2361[7:0];
  _RAND_2362 = {1{`RANDOM}};
  amplifier_1_0_data_132 = _RAND_2362[7:0];
  _RAND_2363 = {1{`RANDOM}};
  amplifier_1_0_data_133 = _RAND_2363[7:0];
  _RAND_2364 = {1{`RANDOM}};
  amplifier_1_0_data_134 = _RAND_2364[7:0];
  _RAND_2365 = {1{`RANDOM}};
  amplifier_1_0_data_135 = _RAND_2365[7:0];
  _RAND_2366 = {1{`RANDOM}};
  amplifier_1_0_data_136 = _RAND_2366[7:0];
  _RAND_2367 = {1{`RANDOM}};
  amplifier_1_0_data_137 = _RAND_2367[7:0];
  _RAND_2368 = {1{`RANDOM}};
  amplifier_1_0_data_138 = _RAND_2368[7:0];
  _RAND_2369 = {1{`RANDOM}};
  amplifier_1_0_data_139 = _RAND_2369[7:0];
  _RAND_2370 = {1{`RANDOM}};
  amplifier_1_0_data_140 = _RAND_2370[7:0];
  _RAND_2371 = {1{`RANDOM}};
  amplifier_1_0_data_141 = _RAND_2371[7:0];
  _RAND_2372 = {1{`RANDOM}};
  amplifier_1_0_data_142 = _RAND_2372[7:0];
  _RAND_2373 = {1{`RANDOM}};
  amplifier_1_0_data_143 = _RAND_2373[7:0];
  _RAND_2374 = {1{`RANDOM}};
  amplifier_1_0_data_144 = _RAND_2374[7:0];
  _RAND_2375 = {1{`RANDOM}};
  amplifier_1_0_data_145 = _RAND_2375[7:0];
  _RAND_2376 = {1{`RANDOM}};
  amplifier_1_0_data_146 = _RAND_2376[7:0];
  _RAND_2377 = {1{`RANDOM}};
  amplifier_1_0_data_147 = _RAND_2377[7:0];
  _RAND_2378 = {1{`RANDOM}};
  amplifier_1_0_data_148 = _RAND_2378[7:0];
  _RAND_2379 = {1{`RANDOM}};
  amplifier_1_0_data_149 = _RAND_2379[7:0];
  _RAND_2380 = {1{`RANDOM}};
  amplifier_1_0_data_150 = _RAND_2380[7:0];
  _RAND_2381 = {1{`RANDOM}};
  amplifier_1_0_data_151 = _RAND_2381[7:0];
  _RAND_2382 = {1{`RANDOM}};
  amplifier_1_0_data_152 = _RAND_2382[7:0];
  _RAND_2383 = {1{`RANDOM}};
  amplifier_1_0_data_153 = _RAND_2383[7:0];
  _RAND_2384 = {1{`RANDOM}};
  amplifier_1_0_data_154 = _RAND_2384[7:0];
  _RAND_2385 = {1{`RANDOM}};
  amplifier_1_0_data_155 = _RAND_2385[7:0];
  _RAND_2386 = {1{`RANDOM}};
  amplifier_1_0_data_156 = _RAND_2386[7:0];
  _RAND_2387 = {1{`RANDOM}};
  amplifier_1_0_data_157 = _RAND_2387[7:0];
  _RAND_2388 = {1{`RANDOM}};
  amplifier_1_0_data_158 = _RAND_2388[7:0];
  _RAND_2389 = {1{`RANDOM}};
  amplifier_1_0_data_159 = _RAND_2389[7:0];
  _RAND_2390 = {1{`RANDOM}};
  amplifier_1_0_data_160 = _RAND_2390[7:0];
  _RAND_2391 = {1{`RANDOM}};
  amplifier_1_0_data_161 = _RAND_2391[7:0];
  _RAND_2392 = {1{`RANDOM}};
  amplifier_1_0_data_162 = _RAND_2392[7:0];
  _RAND_2393 = {1{`RANDOM}};
  amplifier_1_0_data_163 = _RAND_2393[7:0];
  _RAND_2394 = {1{`RANDOM}};
  amplifier_1_0_data_164 = _RAND_2394[7:0];
  _RAND_2395 = {1{`RANDOM}};
  amplifier_1_0_data_165 = _RAND_2395[7:0];
  _RAND_2396 = {1{`RANDOM}};
  amplifier_1_0_data_166 = _RAND_2396[7:0];
  _RAND_2397 = {1{`RANDOM}};
  amplifier_1_0_data_167 = _RAND_2397[7:0];
  _RAND_2398 = {1{`RANDOM}};
  amplifier_1_0_data_168 = _RAND_2398[7:0];
  _RAND_2399 = {1{`RANDOM}};
  amplifier_1_0_data_169 = _RAND_2399[7:0];
  _RAND_2400 = {1{`RANDOM}};
  amplifier_1_0_data_170 = _RAND_2400[7:0];
  _RAND_2401 = {1{`RANDOM}};
  amplifier_1_0_data_171 = _RAND_2401[7:0];
  _RAND_2402 = {1{`RANDOM}};
  amplifier_1_0_data_172 = _RAND_2402[7:0];
  _RAND_2403 = {1{`RANDOM}};
  amplifier_1_0_data_173 = _RAND_2403[7:0];
  _RAND_2404 = {1{`RANDOM}};
  amplifier_1_0_data_174 = _RAND_2404[7:0];
  _RAND_2405 = {1{`RANDOM}};
  amplifier_1_0_data_175 = _RAND_2405[7:0];
  _RAND_2406 = {1{`RANDOM}};
  amplifier_1_0_data_176 = _RAND_2406[7:0];
  _RAND_2407 = {1{`RANDOM}};
  amplifier_1_0_data_177 = _RAND_2407[7:0];
  _RAND_2408 = {1{`RANDOM}};
  amplifier_1_0_data_178 = _RAND_2408[7:0];
  _RAND_2409 = {1{`RANDOM}};
  amplifier_1_0_data_179 = _RAND_2409[7:0];
  _RAND_2410 = {1{`RANDOM}};
  amplifier_1_0_data_180 = _RAND_2410[7:0];
  _RAND_2411 = {1{`RANDOM}};
  amplifier_1_0_data_181 = _RAND_2411[7:0];
  _RAND_2412 = {1{`RANDOM}};
  amplifier_1_0_data_182 = _RAND_2412[7:0];
  _RAND_2413 = {1{`RANDOM}};
  amplifier_1_0_data_183 = _RAND_2413[7:0];
  _RAND_2414 = {1{`RANDOM}};
  amplifier_1_0_data_184 = _RAND_2414[7:0];
  _RAND_2415 = {1{`RANDOM}};
  amplifier_1_0_data_185 = _RAND_2415[7:0];
  _RAND_2416 = {1{`RANDOM}};
  amplifier_1_0_data_186 = _RAND_2416[7:0];
  _RAND_2417 = {1{`RANDOM}};
  amplifier_1_0_data_187 = _RAND_2417[7:0];
  _RAND_2418 = {1{`RANDOM}};
  amplifier_1_0_data_188 = _RAND_2418[7:0];
  _RAND_2419 = {1{`RANDOM}};
  amplifier_1_0_data_189 = _RAND_2419[7:0];
  _RAND_2420 = {1{`RANDOM}};
  amplifier_1_0_data_190 = _RAND_2420[7:0];
  _RAND_2421 = {1{`RANDOM}};
  amplifier_1_0_data_191 = _RAND_2421[7:0];
  _RAND_2422 = {1{`RANDOM}};
  amplifier_1_0_data_192 = _RAND_2422[7:0];
  _RAND_2423 = {1{`RANDOM}};
  amplifier_1_0_data_193 = _RAND_2423[7:0];
  _RAND_2424 = {1{`RANDOM}};
  amplifier_1_0_data_194 = _RAND_2424[7:0];
  _RAND_2425 = {1{`RANDOM}};
  amplifier_1_0_data_195 = _RAND_2425[7:0];
  _RAND_2426 = {1{`RANDOM}};
  amplifier_1_0_data_196 = _RAND_2426[7:0];
  _RAND_2427 = {1{`RANDOM}};
  amplifier_1_0_data_197 = _RAND_2427[7:0];
  _RAND_2428 = {1{`RANDOM}};
  amplifier_1_0_data_198 = _RAND_2428[7:0];
  _RAND_2429 = {1{`RANDOM}};
  amplifier_1_0_data_199 = _RAND_2429[7:0];
  _RAND_2430 = {1{`RANDOM}};
  amplifier_1_0_data_200 = _RAND_2430[7:0];
  _RAND_2431 = {1{`RANDOM}};
  amplifier_1_0_data_201 = _RAND_2431[7:0];
  _RAND_2432 = {1{`RANDOM}};
  amplifier_1_0_data_202 = _RAND_2432[7:0];
  _RAND_2433 = {1{`RANDOM}};
  amplifier_1_0_data_203 = _RAND_2433[7:0];
  _RAND_2434 = {1{`RANDOM}};
  amplifier_1_0_data_204 = _RAND_2434[7:0];
  _RAND_2435 = {1{`RANDOM}};
  amplifier_1_0_data_205 = _RAND_2435[7:0];
  _RAND_2436 = {1{`RANDOM}};
  amplifier_1_0_data_206 = _RAND_2436[7:0];
  _RAND_2437 = {1{`RANDOM}};
  amplifier_1_0_data_207 = _RAND_2437[7:0];
  _RAND_2438 = {1{`RANDOM}};
  amplifier_1_0_data_208 = _RAND_2438[7:0];
  _RAND_2439 = {1{`RANDOM}};
  amplifier_1_0_data_209 = _RAND_2439[7:0];
  _RAND_2440 = {1{`RANDOM}};
  amplifier_1_0_data_210 = _RAND_2440[7:0];
  _RAND_2441 = {1{`RANDOM}};
  amplifier_1_0_data_211 = _RAND_2441[7:0];
  _RAND_2442 = {1{`RANDOM}};
  amplifier_1_0_data_212 = _RAND_2442[7:0];
  _RAND_2443 = {1{`RANDOM}};
  amplifier_1_0_data_213 = _RAND_2443[7:0];
  _RAND_2444 = {1{`RANDOM}};
  amplifier_1_0_data_214 = _RAND_2444[7:0];
  _RAND_2445 = {1{`RANDOM}};
  amplifier_1_0_data_215 = _RAND_2445[7:0];
  _RAND_2446 = {1{`RANDOM}};
  amplifier_1_0_data_216 = _RAND_2446[7:0];
  _RAND_2447 = {1{`RANDOM}};
  amplifier_1_0_data_217 = _RAND_2447[7:0];
  _RAND_2448 = {1{`RANDOM}};
  amplifier_1_0_data_218 = _RAND_2448[7:0];
  _RAND_2449 = {1{`RANDOM}};
  amplifier_1_0_data_219 = _RAND_2449[7:0];
  _RAND_2450 = {1{`RANDOM}};
  amplifier_1_0_data_220 = _RAND_2450[7:0];
  _RAND_2451 = {1{`RANDOM}};
  amplifier_1_0_data_221 = _RAND_2451[7:0];
  _RAND_2452 = {1{`RANDOM}};
  amplifier_1_0_data_222 = _RAND_2452[7:0];
  _RAND_2453 = {1{`RANDOM}};
  amplifier_1_0_data_223 = _RAND_2453[7:0];
  _RAND_2454 = {1{`RANDOM}};
  amplifier_1_0_data_224 = _RAND_2454[7:0];
  _RAND_2455 = {1{`RANDOM}};
  amplifier_1_0_data_225 = _RAND_2455[7:0];
  _RAND_2456 = {1{`RANDOM}};
  amplifier_1_0_data_226 = _RAND_2456[7:0];
  _RAND_2457 = {1{`RANDOM}};
  amplifier_1_0_data_227 = _RAND_2457[7:0];
  _RAND_2458 = {1{`RANDOM}};
  amplifier_1_0_data_228 = _RAND_2458[7:0];
  _RAND_2459 = {1{`RANDOM}};
  amplifier_1_0_data_229 = _RAND_2459[7:0];
  _RAND_2460 = {1{`RANDOM}};
  amplifier_1_0_data_230 = _RAND_2460[7:0];
  _RAND_2461 = {1{`RANDOM}};
  amplifier_1_0_data_231 = _RAND_2461[7:0];
  _RAND_2462 = {1{`RANDOM}};
  amplifier_1_0_data_232 = _RAND_2462[7:0];
  _RAND_2463 = {1{`RANDOM}};
  amplifier_1_0_data_233 = _RAND_2463[7:0];
  _RAND_2464 = {1{`RANDOM}};
  amplifier_1_0_data_234 = _RAND_2464[7:0];
  _RAND_2465 = {1{`RANDOM}};
  amplifier_1_0_data_235 = _RAND_2465[7:0];
  _RAND_2466 = {1{`RANDOM}};
  amplifier_1_0_data_236 = _RAND_2466[7:0];
  _RAND_2467 = {1{`RANDOM}};
  amplifier_1_0_data_237 = _RAND_2467[7:0];
  _RAND_2468 = {1{`RANDOM}};
  amplifier_1_0_data_238 = _RAND_2468[7:0];
  _RAND_2469 = {1{`RANDOM}};
  amplifier_1_0_data_239 = _RAND_2469[7:0];
  _RAND_2470 = {1{`RANDOM}};
  amplifier_1_0_data_240 = _RAND_2470[7:0];
  _RAND_2471 = {1{`RANDOM}};
  amplifier_1_0_data_241 = _RAND_2471[7:0];
  _RAND_2472 = {1{`RANDOM}};
  amplifier_1_0_data_242 = _RAND_2472[7:0];
  _RAND_2473 = {1{`RANDOM}};
  amplifier_1_0_data_243 = _RAND_2473[7:0];
  _RAND_2474 = {1{`RANDOM}};
  amplifier_1_0_data_244 = _RAND_2474[7:0];
  _RAND_2475 = {1{`RANDOM}};
  amplifier_1_0_data_245 = _RAND_2475[7:0];
  _RAND_2476 = {1{`RANDOM}};
  amplifier_1_0_data_246 = _RAND_2476[7:0];
  _RAND_2477 = {1{`RANDOM}};
  amplifier_1_0_data_247 = _RAND_2477[7:0];
  _RAND_2478 = {1{`RANDOM}};
  amplifier_1_0_data_248 = _RAND_2478[7:0];
  _RAND_2479 = {1{`RANDOM}};
  amplifier_1_0_data_249 = _RAND_2479[7:0];
  _RAND_2480 = {1{`RANDOM}};
  amplifier_1_0_data_250 = _RAND_2480[7:0];
  _RAND_2481 = {1{`RANDOM}};
  amplifier_1_0_data_251 = _RAND_2481[7:0];
  _RAND_2482 = {1{`RANDOM}};
  amplifier_1_0_data_252 = _RAND_2482[7:0];
  _RAND_2483 = {1{`RANDOM}};
  amplifier_1_0_data_253 = _RAND_2483[7:0];
  _RAND_2484 = {1{`RANDOM}};
  amplifier_1_0_data_254 = _RAND_2484[7:0];
  _RAND_2485 = {1{`RANDOM}};
  amplifier_1_0_data_255 = _RAND_2485[7:0];
  _RAND_2486 = {1{`RANDOM}};
  amplifier_1_0_header_0 = _RAND_2486[15:0];
  _RAND_2487 = {1{`RANDOM}};
  amplifier_1_0_header_1 = _RAND_2487[15:0];
  _RAND_2488 = {1{`RANDOM}};
  amplifier_1_0_header_2 = _RAND_2488[15:0];
  _RAND_2489 = {1{`RANDOM}};
  amplifier_1_0_header_3 = _RAND_2489[15:0];
  _RAND_2490 = {1{`RANDOM}};
  amplifier_1_0_header_4 = _RAND_2490[15:0];
  _RAND_2491 = {1{`RANDOM}};
  amplifier_1_0_header_5 = _RAND_2491[15:0];
  _RAND_2492 = {1{`RANDOM}};
  amplifier_1_0_header_6 = _RAND_2492[15:0];
  _RAND_2493 = {1{`RANDOM}};
  amplifier_1_0_header_7 = _RAND_2493[15:0];
  _RAND_2494 = {1{`RANDOM}};
  amplifier_1_0_header_8 = _RAND_2494[15:0];
  _RAND_2495 = {1{`RANDOM}};
  amplifier_1_0_header_9 = _RAND_2495[15:0];
  _RAND_2496 = {1{`RANDOM}};
  amplifier_1_0_header_10 = _RAND_2496[15:0];
  _RAND_2497 = {1{`RANDOM}};
  amplifier_1_0_header_11 = _RAND_2497[15:0];
  _RAND_2498 = {1{`RANDOM}};
  amplifier_1_0_header_12 = _RAND_2498[15:0];
  _RAND_2499 = {1{`RANDOM}};
  amplifier_1_0_header_13 = _RAND_2499[15:0];
  _RAND_2500 = {1{`RANDOM}};
  amplifier_1_0_header_14 = _RAND_2500[15:0];
  _RAND_2501 = {1{`RANDOM}};
  amplifier_1_0_header_15 = _RAND_2501[15:0];
  _RAND_2502 = {1{`RANDOM}};
  amplifier_1_0_parse_current_state = _RAND_2502[7:0];
  _RAND_2503 = {1{`RANDOM}};
  amplifier_1_0_parse_current_offset = _RAND_2503[7:0];
  _RAND_2504 = {1{`RANDOM}};
  amplifier_1_0_parse_transition_field = _RAND_2504[15:0];
  _RAND_2505 = {1{`RANDOM}};
  amplifier_1_0_next_processor_id = _RAND_2505[1:0];
  _RAND_2506 = {1{`RANDOM}};
  amplifier_1_0_next_config_id = _RAND_2506[0:0];
  _RAND_2507 = {1{`RANDOM}};
  amplifier_1_0_is_valid_processor = _RAND_2507[0:0];
  _RAND_2508 = {1{`RANDOM}};
  amplifier_1_1_data_0 = _RAND_2508[7:0];
  _RAND_2509 = {1{`RANDOM}};
  amplifier_1_1_data_1 = _RAND_2509[7:0];
  _RAND_2510 = {1{`RANDOM}};
  amplifier_1_1_data_2 = _RAND_2510[7:0];
  _RAND_2511 = {1{`RANDOM}};
  amplifier_1_1_data_3 = _RAND_2511[7:0];
  _RAND_2512 = {1{`RANDOM}};
  amplifier_1_1_data_4 = _RAND_2512[7:0];
  _RAND_2513 = {1{`RANDOM}};
  amplifier_1_1_data_5 = _RAND_2513[7:0];
  _RAND_2514 = {1{`RANDOM}};
  amplifier_1_1_data_6 = _RAND_2514[7:0];
  _RAND_2515 = {1{`RANDOM}};
  amplifier_1_1_data_7 = _RAND_2515[7:0];
  _RAND_2516 = {1{`RANDOM}};
  amplifier_1_1_data_8 = _RAND_2516[7:0];
  _RAND_2517 = {1{`RANDOM}};
  amplifier_1_1_data_9 = _RAND_2517[7:0];
  _RAND_2518 = {1{`RANDOM}};
  amplifier_1_1_data_10 = _RAND_2518[7:0];
  _RAND_2519 = {1{`RANDOM}};
  amplifier_1_1_data_11 = _RAND_2519[7:0];
  _RAND_2520 = {1{`RANDOM}};
  amplifier_1_1_data_12 = _RAND_2520[7:0];
  _RAND_2521 = {1{`RANDOM}};
  amplifier_1_1_data_13 = _RAND_2521[7:0];
  _RAND_2522 = {1{`RANDOM}};
  amplifier_1_1_data_14 = _RAND_2522[7:0];
  _RAND_2523 = {1{`RANDOM}};
  amplifier_1_1_data_15 = _RAND_2523[7:0];
  _RAND_2524 = {1{`RANDOM}};
  amplifier_1_1_data_16 = _RAND_2524[7:0];
  _RAND_2525 = {1{`RANDOM}};
  amplifier_1_1_data_17 = _RAND_2525[7:0];
  _RAND_2526 = {1{`RANDOM}};
  amplifier_1_1_data_18 = _RAND_2526[7:0];
  _RAND_2527 = {1{`RANDOM}};
  amplifier_1_1_data_19 = _RAND_2527[7:0];
  _RAND_2528 = {1{`RANDOM}};
  amplifier_1_1_data_20 = _RAND_2528[7:0];
  _RAND_2529 = {1{`RANDOM}};
  amplifier_1_1_data_21 = _RAND_2529[7:0];
  _RAND_2530 = {1{`RANDOM}};
  amplifier_1_1_data_22 = _RAND_2530[7:0];
  _RAND_2531 = {1{`RANDOM}};
  amplifier_1_1_data_23 = _RAND_2531[7:0];
  _RAND_2532 = {1{`RANDOM}};
  amplifier_1_1_data_24 = _RAND_2532[7:0];
  _RAND_2533 = {1{`RANDOM}};
  amplifier_1_1_data_25 = _RAND_2533[7:0];
  _RAND_2534 = {1{`RANDOM}};
  amplifier_1_1_data_26 = _RAND_2534[7:0];
  _RAND_2535 = {1{`RANDOM}};
  amplifier_1_1_data_27 = _RAND_2535[7:0];
  _RAND_2536 = {1{`RANDOM}};
  amplifier_1_1_data_28 = _RAND_2536[7:0];
  _RAND_2537 = {1{`RANDOM}};
  amplifier_1_1_data_29 = _RAND_2537[7:0];
  _RAND_2538 = {1{`RANDOM}};
  amplifier_1_1_data_30 = _RAND_2538[7:0];
  _RAND_2539 = {1{`RANDOM}};
  amplifier_1_1_data_31 = _RAND_2539[7:0];
  _RAND_2540 = {1{`RANDOM}};
  amplifier_1_1_data_32 = _RAND_2540[7:0];
  _RAND_2541 = {1{`RANDOM}};
  amplifier_1_1_data_33 = _RAND_2541[7:0];
  _RAND_2542 = {1{`RANDOM}};
  amplifier_1_1_data_34 = _RAND_2542[7:0];
  _RAND_2543 = {1{`RANDOM}};
  amplifier_1_1_data_35 = _RAND_2543[7:0];
  _RAND_2544 = {1{`RANDOM}};
  amplifier_1_1_data_36 = _RAND_2544[7:0];
  _RAND_2545 = {1{`RANDOM}};
  amplifier_1_1_data_37 = _RAND_2545[7:0];
  _RAND_2546 = {1{`RANDOM}};
  amplifier_1_1_data_38 = _RAND_2546[7:0];
  _RAND_2547 = {1{`RANDOM}};
  amplifier_1_1_data_39 = _RAND_2547[7:0];
  _RAND_2548 = {1{`RANDOM}};
  amplifier_1_1_data_40 = _RAND_2548[7:0];
  _RAND_2549 = {1{`RANDOM}};
  amplifier_1_1_data_41 = _RAND_2549[7:0];
  _RAND_2550 = {1{`RANDOM}};
  amplifier_1_1_data_42 = _RAND_2550[7:0];
  _RAND_2551 = {1{`RANDOM}};
  amplifier_1_1_data_43 = _RAND_2551[7:0];
  _RAND_2552 = {1{`RANDOM}};
  amplifier_1_1_data_44 = _RAND_2552[7:0];
  _RAND_2553 = {1{`RANDOM}};
  amplifier_1_1_data_45 = _RAND_2553[7:0];
  _RAND_2554 = {1{`RANDOM}};
  amplifier_1_1_data_46 = _RAND_2554[7:0];
  _RAND_2555 = {1{`RANDOM}};
  amplifier_1_1_data_47 = _RAND_2555[7:0];
  _RAND_2556 = {1{`RANDOM}};
  amplifier_1_1_data_48 = _RAND_2556[7:0];
  _RAND_2557 = {1{`RANDOM}};
  amplifier_1_1_data_49 = _RAND_2557[7:0];
  _RAND_2558 = {1{`RANDOM}};
  amplifier_1_1_data_50 = _RAND_2558[7:0];
  _RAND_2559 = {1{`RANDOM}};
  amplifier_1_1_data_51 = _RAND_2559[7:0];
  _RAND_2560 = {1{`RANDOM}};
  amplifier_1_1_data_52 = _RAND_2560[7:0];
  _RAND_2561 = {1{`RANDOM}};
  amplifier_1_1_data_53 = _RAND_2561[7:0];
  _RAND_2562 = {1{`RANDOM}};
  amplifier_1_1_data_54 = _RAND_2562[7:0];
  _RAND_2563 = {1{`RANDOM}};
  amplifier_1_1_data_55 = _RAND_2563[7:0];
  _RAND_2564 = {1{`RANDOM}};
  amplifier_1_1_data_56 = _RAND_2564[7:0];
  _RAND_2565 = {1{`RANDOM}};
  amplifier_1_1_data_57 = _RAND_2565[7:0];
  _RAND_2566 = {1{`RANDOM}};
  amplifier_1_1_data_58 = _RAND_2566[7:0];
  _RAND_2567 = {1{`RANDOM}};
  amplifier_1_1_data_59 = _RAND_2567[7:0];
  _RAND_2568 = {1{`RANDOM}};
  amplifier_1_1_data_60 = _RAND_2568[7:0];
  _RAND_2569 = {1{`RANDOM}};
  amplifier_1_1_data_61 = _RAND_2569[7:0];
  _RAND_2570 = {1{`RANDOM}};
  amplifier_1_1_data_62 = _RAND_2570[7:0];
  _RAND_2571 = {1{`RANDOM}};
  amplifier_1_1_data_63 = _RAND_2571[7:0];
  _RAND_2572 = {1{`RANDOM}};
  amplifier_1_1_data_64 = _RAND_2572[7:0];
  _RAND_2573 = {1{`RANDOM}};
  amplifier_1_1_data_65 = _RAND_2573[7:0];
  _RAND_2574 = {1{`RANDOM}};
  amplifier_1_1_data_66 = _RAND_2574[7:0];
  _RAND_2575 = {1{`RANDOM}};
  amplifier_1_1_data_67 = _RAND_2575[7:0];
  _RAND_2576 = {1{`RANDOM}};
  amplifier_1_1_data_68 = _RAND_2576[7:0];
  _RAND_2577 = {1{`RANDOM}};
  amplifier_1_1_data_69 = _RAND_2577[7:0];
  _RAND_2578 = {1{`RANDOM}};
  amplifier_1_1_data_70 = _RAND_2578[7:0];
  _RAND_2579 = {1{`RANDOM}};
  amplifier_1_1_data_71 = _RAND_2579[7:0];
  _RAND_2580 = {1{`RANDOM}};
  amplifier_1_1_data_72 = _RAND_2580[7:0];
  _RAND_2581 = {1{`RANDOM}};
  amplifier_1_1_data_73 = _RAND_2581[7:0];
  _RAND_2582 = {1{`RANDOM}};
  amplifier_1_1_data_74 = _RAND_2582[7:0];
  _RAND_2583 = {1{`RANDOM}};
  amplifier_1_1_data_75 = _RAND_2583[7:0];
  _RAND_2584 = {1{`RANDOM}};
  amplifier_1_1_data_76 = _RAND_2584[7:0];
  _RAND_2585 = {1{`RANDOM}};
  amplifier_1_1_data_77 = _RAND_2585[7:0];
  _RAND_2586 = {1{`RANDOM}};
  amplifier_1_1_data_78 = _RAND_2586[7:0];
  _RAND_2587 = {1{`RANDOM}};
  amplifier_1_1_data_79 = _RAND_2587[7:0];
  _RAND_2588 = {1{`RANDOM}};
  amplifier_1_1_data_80 = _RAND_2588[7:0];
  _RAND_2589 = {1{`RANDOM}};
  amplifier_1_1_data_81 = _RAND_2589[7:0];
  _RAND_2590 = {1{`RANDOM}};
  amplifier_1_1_data_82 = _RAND_2590[7:0];
  _RAND_2591 = {1{`RANDOM}};
  amplifier_1_1_data_83 = _RAND_2591[7:0];
  _RAND_2592 = {1{`RANDOM}};
  amplifier_1_1_data_84 = _RAND_2592[7:0];
  _RAND_2593 = {1{`RANDOM}};
  amplifier_1_1_data_85 = _RAND_2593[7:0];
  _RAND_2594 = {1{`RANDOM}};
  amplifier_1_1_data_86 = _RAND_2594[7:0];
  _RAND_2595 = {1{`RANDOM}};
  amplifier_1_1_data_87 = _RAND_2595[7:0];
  _RAND_2596 = {1{`RANDOM}};
  amplifier_1_1_data_88 = _RAND_2596[7:0];
  _RAND_2597 = {1{`RANDOM}};
  amplifier_1_1_data_89 = _RAND_2597[7:0];
  _RAND_2598 = {1{`RANDOM}};
  amplifier_1_1_data_90 = _RAND_2598[7:0];
  _RAND_2599 = {1{`RANDOM}};
  amplifier_1_1_data_91 = _RAND_2599[7:0];
  _RAND_2600 = {1{`RANDOM}};
  amplifier_1_1_data_92 = _RAND_2600[7:0];
  _RAND_2601 = {1{`RANDOM}};
  amplifier_1_1_data_93 = _RAND_2601[7:0];
  _RAND_2602 = {1{`RANDOM}};
  amplifier_1_1_data_94 = _RAND_2602[7:0];
  _RAND_2603 = {1{`RANDOM}};
  amplifier_1_1_data_95 = _RAND_2603[7:0];
  _RAND_2604 = {1{`RANDOM}};
  amplifier_1_1_data_96 = _RAND_2604[7:0];
  _RAND_2605 = {1{`RANDOM}};
  amplifier_1_1_data_97 = _RAND_2605[7:0];
  _RAND_2606 = {1{`RANDOM}};
  amplifier_1_1_data_98 = _RAND_2606[7:0];
  _RAND_2607 = {1{`RANDOM}};
  amplifier_1_1_data_99 = _RAND_2607[7:0];
  _RAND_2608 = {1{`RANDOM}};
  amplifier_1_1_data_100 = _RAND_2608[7:0];
  _RAND_2609 = {1{`RANDOM}};
  amplifier_1_1_data_101 = _RAND_2609[7:0];
  _RAND_2610 = {1{`RANDOM}};
  amplifier_1_1_data_102 = _RAND_2610[7:0];
  _RAND_2611 = {1{`RANDOM}};
  amplifier_1_1_data_103 = _RAND_2611[7:0];
  _RAND_2612 = {1{`RANDOM}};
  amplifier_1_1_data_104 = _RAND_2612[7:0];
  _RAND_2613 = {1{`RANDOM}};
  amplifier_1_1_data_105 = _RAND_2613[7:0];
  _RAND_2614 = {1{`RANDOM}};
  amplifier_1_1_data_106 = _RAND_2614[7:0];
  _RAND_2615 = {1{`RANDOM}};
  amplifier_1_1_data_107 = _RAND_2615[7:0];
  _RAND_2616 = {1{`RANDOM}};
  amplifier_1_1_data_108 = _RAND_2616[7:0];
  _RAND_2617 = {1{`RANDOM}};
  amplifier_1_1_data_109 = _RAND_2617[7:0];
  _RAND_2618 = {1{`RANDOM}};
  amplifier_1_1_data_110 = _RAND_2618[7:0];
  _RAND_2619 = {1{`RANDOM}};
  amplifier_1_1_data_111 = _RAND_2619[7:0];
  _RAND_2620 = {1{`RANDOM}};
  amplifier_1_1_data_112 = _RAND_2620[7:0];
  _RAND_2621 = {1{`RANDOM}};
  amplifier_1_1_data_113 = _RAND_2621[7:0];
  _RAND_2622 = {1{`RANDOM}};
  amplifier_1_1_data_114 = _RAND_2622[7:0];
  _RAND_2623 = {1{`RANDOM}};
  amplifier_1_1_data_115 = _RAND_2623[7:0];
  _RAND_2624 = {1{`RANDOM}};
  amplifier_1_1_data_116 = _RAND_2624[7:0];
  _RAND_2625 = {1{`RANDOM}};
  amplifier_1_1_data_117 = _RAND_2625[7:0];
  _RAND_2626 = {1{`RANDOM}};
  amplifier_1_1_data_118 = _RAND_2626[7:0];
  _RAND_2627 = {1{`RANDOM}};
  amplifier_1_1_data_119 = _RAND_2627[7:0];
  _RAND_2628 = {1{`RANDOM}};
  amplifier_1_1_data_120 = _RAND_2628[7:0];
  _RAND_2629 = {1{`RANDOM}};
  amplifier_1_1_data_121 = _RAND_2629[7:0];
  _RAND_2630 = {1{`RANDOM}};
  amplifier_1_1_data_122 = _RAND_2630[7:0];
  _RAND_2631 = {1{`RANDOM}};
  amplifier_1_1_data_123 = _RAND_2631[7:0];
  _RAND_2632 = {1{`RANDOM}};
  amplifier_1_1_data_124 = _RAND_2632[7:0];
  _RAND_2633 = {1{`RANDOM}};
  amplifier_1_1_data_125 = _RAND_2633[7:0];
  _RAND_2634 = {1{`RANDOM}};
  amplifier_1_1_data_126 = _RAND_2634[7:0];
  _RAND_2635 = {1{`RANDOM}};
  amplifier_1_1_data_127 = _RAND_2635[7:0];
  _RAND_2636 = {1{`RANDOM}};
  amplifier_1_1_data_128 = _RAND_2636[7:0];
  _RAND_2637 = {1{`RANDOM}};
  amplifier_1_1_data_129 = _RAND_2637[7:0];
  _RAND_2638 = {1{`RANDOM}};
  amplifier_1_1_data_130 = _RAND_2638[7:0];
  _RAND_2639 = {1{`RANDOM}};
  amplifier_1_1_data_131 = _RAND_2639[7:0];
  _RAND_2640 = {1{`RANDOM}};
  amplifier_1_1_data_132 = _RAND_2640[7:0];
  _RAND_2641 = {1{`RANDOM}};
  amplifier_1_1_data_133 = _RAND_2641[7:0];
  _RAND_2642 = {1{`RANDOM}};
  amplifier_1_1_data_134 = _RAND_2642[7:0];
  _RAND_2643 = {1{`RANDOM}};
  amplifier_1_1_data_135 = _RAND_2643[7:0];
  _RAND_2644 = {1{`RANDOM}};
  amplifier_1_1_data_136 = _RAND_2644[7:0];
  _RAND_2645 = {1{`RANDOM}};
  amplifier_1_1_data_137 = _RAND_2645[7:0];
  _RAND_2646 = {1{`RANDOM}};
  amplifier_1_1_data_138 = _RAND_2646[7:0];
  _RAND_2647 = {1{`RANDOM}};
  amplifier_1_1_data_139 = _RAND_2647[7:0];
  _RAND_2648 = {1{`RANDOM}};
  amplifier_1_1_data_140 = _RAND_2648[7:0];
  _RAND_2649 = {1{`RANDOM}};
  amplifier_1_1_data_141 = _RAND_2649[7:0];
  _RAND_2650 = {1{`RANDOM}};
  amplifier_1_1_data_142 = _RAND_2650[7:0];
  _RAND_2651 = {1{`RANDOM}};
  amplifier_1_1_data_143 = _RAND_2651[7:0];
  _RAND_2652 = {1{`RANDOM}};
  amplifier_1_1_data_144 = _RAND_2652[7:0];
  _RAND_2653 = {1{`RANDOM}};
  amplifier_1_1_data_145 = _RAND_2653[7:0];
  _RAND_2654 = {1{`RANDOM}};
  amplifier_1_1_data_146 = _RAND_2654[7:0];
  _RAND_2655 = {1{`RANDOM}};
  amplifier_1_1_data_147 = _RAND_2655[7:0];
  _RAND_2656 = {1{`RANDOM}};
  amplifier_1_1_data_148 = _RAND_2656[7:0];
  _RAND_2657 = {1{`RANDOM}};
  amplifier_1_1_data_149 = _RAND_2657[7:0];
  _RAND_2658 = {1{`RANDOM}};
  amplifier_1_1_data_150 = _RAND_2658[7:0];
  _RAND_2659 = {1{`RANDOM}};
  amplifier_1_1_data_151 = _RAND_2659[7:0];
  _RAND_2660 = {1{`RANDOM}};
  amplifier_1_1_data_152 = _RAND_2660[7:0];
  _RAND_2661 = {1{`RANDOM}};
  amplifier_1_1_data_153 = _RAND_2661[7:0];
  _RAND_2662 = {1{`RANDOM}};
  amplifier_1_1_data_154 = _RAND_2662[7:0];
  _RAND_2663 = {1{`RANDOM}};
  amplifier_1_1_data_155 = _RAND_2663[7:0];
  _RAND_2664 = {1{`RANDOM}};
  amplifier_1_1_data_156 = _RAND_2664[7:0];
  _RAND_2665 = {1{`RANDOM}};
  amplifier_1_1_data_157 = _RAND_2665[7:0];
  _RAND_2666 = {1{`RANDOM}};
  amplifier_1_1_data_158 = _RAND_2666[7:0];
  _RAND_2667 = {1{`RANDOM}};
  amplifier_1_1_data_159 = _RAND_2667[7:0];
  _RAND_2668 = {1{`RANDOM}};
  amplifier_1_1_data_160 = _RAND_2668[7:0];
  _RAND_2669 = {1{`RANDOM}};
  amplifier_1_1_data_161 = _RAND_2669[7:0];
  _RAND_2670 = {1{`RANDOM}};
  amplifier_1_1_data_162 = _RAND_2670[7:0];
  _RAND_2671 = {1{`RANDOM}};
  amplifier_1_1_data_163 = _RAND_2671[7:0];
  _RAND_2672 = {1{`RANDOM}};
  amplifier_1_1_data_164 = _RAND_2672[7:0];
  _RAND_2673 = {1{`RANDOM}};
  amplifier_1_1_data_165 = _RAND_2673[7:0];
  _RAND_2674 = {1{`RANDOM}};
  amplifier_1_1_data_166 = _RAND_2674[7:0];
  _RAND_2675 = {1{`RANDOM}};
  amplifier_1_1_data_167 = _RAND_2675[7:0];
  _RAND_2676 = {1{`RANDOM}};
  amplifier_1_1_data_168 = _RAND_2676[7:0];
  _RAND_2677 = {1{`RANDOM}};
  amplifier_1_1_data_169 = _RAND_2677[7:0];
  _RAND_2678 = {1{`RANDOM}};
  amplifier_1_1_data_170 = _RAND_2678[7:0];
  _RAND_2679 = {1{`RANDOM}};
  amplifier_1_1_data_171 = _RAND_2679[7:0];
  _RAND_2680 = {1{`RANDOM}};
  amplifier_1_1_data_172 = _RAND_2680[7:0];
  _RAND_2681 = {1{`RANDOM}};
  amplifier_1_1_data_173 = _RAND_2681[7:0];
  _RAND_2682 = {1{`RANDOM}};
  amplifier_1_1_data_174 = _RAND_2682[7:0];
  _RAND_2683 = {1{`RANDOM}};
  amplifier_1_1_data_175 = _RAND_2683[7:0];
  _RAND_2684 = {1{`RANDOM}};
  amplifier_1_1_data_176 = _RAND_2684[7:0];
  _RAND_2685 = {1{`RANDOM}};
  amplifier_1_1_data_177 = _RAND_2685[7:0];
  _RAND_2686 = {1{`RANDOM}};
  amplifier_1_1_data_178 = _RAND_2686[7:0];
  _RAND_2687 = {1{`RANDOM}};
  amplifier_1_1_data_179 = _RAND_2687[7:0];
  _RAND_2688 = {1{`RANDOM}};
  amplifier_1_1_data_180 = _RAND_2688[7:0];
  _RAND_2689 = {1{`RANDOM}};
  amplifier_1_1_data_181 = _RAND_2689[7:0];
  _RAND_2690 = {1{`RANDOM}};
  amplifier_1_1_data_182 = _RAND_2690[7:0];
  _RAND_2691 = {1{`RANDOM}};
  amplifier_1_1_data_183 = _RAND_2691[7:0];
  _RAND_2692 = {1{`RANDOM}};
  amplifier_1_1_data_184 = _RAND_2692[7:0];
  _RAND_2693 = {1{`RANDOM}};
  amplifier_1_1_data_185 = _RAND_2693[7:0];
  _RAND_2694 = {1{`RANDOM}};
  amplifier_1_1_data_186 = _RAND_2694[7:0];
  _RAND_2695 = {1{`RANDOM}};
  amplifier_1_1_data_187 = _RAND_2695[7:0];
  _RAND_2696 = {1{`RANDOM}};
  amplifier_1_1_data_188 = _RAND_2696[7:0];
  _RAND_2697 = {1{`RANDOM}};
  amplifier_1_1_data_189 = _RAND_2697[7:0];
  _RAND_2698 = {1{`RANDOM}};
  amplifier_1_1_data_190 = _RAND_2698[7:0];
  _RAND_2699 = {1{`RANDOM}};
  amplifier_1_1_data_191 = _RAND_2699[7:0];
  _RAND_2700 = {1{`RANDOM}};
  amplifier_1_1_data_192 = _RAND_2700[7:0];
  _RAND_2701 = {1{`RANDOM}};
  amplifier_1_1_data_193 = _RAND_2701[7:0];
  _RAND_2702 = {1{`RANDOM}};
  amplifier_1_1_data_194 = _RAND_2702[7:0];
  _RAND_2703 = {1{`RANDOM}};
  amplifier_1_1_data_195 = _RAND_2703[7:0];
  _RAND_2704 = {1{`RANDOM}};
  amplifier_1_1_data_196 = _RAND_2704[7:0];
  _RAND_2705 = {1{`RANDOM}};
  amplifier_1_1_data_197 = _RAND_2705[7:0];
  _RAND_2706 = {1{`RANDOM}};
  amplifier_1_1_data_198 = _RAND_2706[7:0];
  _RAND_2707 = {1{`RANDOM}};
  amplifier_1_1_data_199 = _RAND_2707[7:0];
  _RAND_2708 = {1{`RANDOM}};
  amplifier_1_1_data_200 = _RAND_2708[7:0];
  _RAND_2709 = {1{`RANDOM}};
  amplifier_1_1_data_201 = _RAND_2709[7:0];
  _RAND_2710 = {1{`RANDOM}};
  amplifier_1_1_data_202 = _RAND_2710[7:0];
  _RAND_2711 = {1{`RANDOM}};
  amplifier_1_1_data_203 = _RAND_2711[7:0];
  _RAND_2712 = {1{`RANDOM}};
  amplifier_1_1_data_204 = _RAND_2712[7:0];
  _RAND_2713 = {1{`RANDOM}};
  amplifier_1_1_data_205 = _RAND_2713[7:0];
  _RAND_2714 = {1{`RANDOM}};
  amplifier_1_1_data_206 = _RAND_2714[7:0];
  _RAND_2715 = {1{`RANDOM}};
  amplifier_1_1_data_207 = _RAND_2715[7:0];
  _RAND_2716 = {1{`RANDOM}};
  amplifier_1_1_data_208 = _RAND_2716[7:0];
  _RAND_2717 = {1{`RANDOM}};
  amplifier_1_1_data_209 = _RAND_2717[7:0];
  _RAND_2718 = {1{`RANDOM}};
  amplifier_1_1_data_210 = _RAND_2718[7:0];
  _RAND_2719 = {1{`RANDOM}};
  amplifier_1_1_data_211 = _RAND_2719[7:0];
  _RAND_2720 = {1{`RANDOM}};
  amplifier_1_1_data_212 = _RAND_2720[7:0];
  _RAND_2721 = {1{`RANDOM}};
  amplifier_1_1_data_213 = _RAND_2721[7:0];
  _RAND_2722 = {1{`RANDOM}};
  amplifier_1_1_data_214 = _RAND_2722[7:0];
  _RAND_2723 = {1{`RANDOM}};
  amplifier_1_1_data_215 = _RAND_2723[7:0];
  _RAND_2724 = {1{`RANDOM}};
  amplifier_1_1_data_216 = _RAND_2724[7:0];
  _RAND_2725 = {1{`RANDOM}};
  amplifier_1_1_data_217 = _RAND_2725[7:0];
  _RAND_2726 = {1{`RANDOM}};
  amplifier_1_1_data_218 = _RAND_2726[7:0];
  _RAND_2727 = {1{`RANDOM}};
  amplifier_1_1_data_219 = _RAND_2727[7:0];
  _RAND_2728 = {1{`RANDOM}};
  amplifier_1_1_data_220 = _RAND_2728[7:0];
  _RAND_2729 = {1{`RANDOM}};
  amplifier_1_1_data_221 = _RAND_2729[7:0];
  _RAND_2730 = {1{`RANDOM}};
  amplifier_1_1_data_222 = _RAND_2730[7:0];
  _RAND_2731 = {1{`RANDOM}};
  amplifier_1_1_data_223 = _RAND_2731[7:0];
  _RAND_2732 = {1{`RANDOM}};
  amplifier_1_1_data_224 = _RAND_2732[7:0];
  _RAND_2733 = {1{`RANDOM}};
  amplifier_1_1_data_225 = _RAND_2733[7:0];
  _RAND_2734 = {1{`RANDOM}};
  amplifier_1_1_data_226 = _RAND_2734[7:0];
  _RAND_2735 = {1{`RANDOM}};
  amplifier_1_1_data_227 = _RAND_2735[7:0];
  _RAND_2736 = {1{`RANDOM}};
  amplifier_1_1_data_228 = _RAND_2736[7:0];
  _RAND_2737 = {1{`RANDOM}};
  amplifier_1_1_data_229 = _RAND_2737[7:0];
  _RAND_2738 = {1{`RANDOM}};
  amplifier_1_1_data_230 = _RAND_2738[7:0];
  _RAND_2739 = {1{`RANDOM}};
  amplifier_1_1_data_231 = _RAND_2739[7:0];
  _RAND_2740 = {1{`RANDOM}};
  amplifier_1_1_data_232 = _RAND_2740[7:0];
  _RAND_2741 = {1{`RANDOM}};
  amplifier_1_1_data_233 = _RAND_2741[7:0];
  _RAND_2742 = {1{`RANDOM}};
  amplifier_1_1_data_234 = _RAND_2742[7:0];
  _RAND_2743 = {1{`RANDOM}};
  amplifier_1_1_data_235 = _RAND_2743[7:0];
  _RAND_2744 = {1{`RANDOM}};
  amplifier_1_1_data_236 = _RAND_2744[7:0];
  _RAND_2745 = {1{`RANDOM}};
  amplifier_1_1_data_237 = _RAND_2745[7:0];
  _RAND_2746 = {1{`RANDOM}};
  amplifier_1_1_data_238 = _RAND_2746[7:0];
  _RAND_2747 = {1{`RANDOM}};
  amplifier_1_1_data_239 = _RAND_2747[7:0];
  _RAND_2748 = {1{`RANDOM}};
  amplifier_1_1_data_240 = _RAND_2748[7:0];
  _RAND_2749 = {1{`RANDOM}};
  amplifier_1_1_data_241 = _RAND_2749[7:0];
  _RAND_2750 = {1{`RANDOM}};
  amplifier_1_1_data_242 = _RAND_2750[7:0];
  _RAND_2751 = {1{`RANDOM}};
  amplifier_1_1_data_243 = _RAND_2751[7:0];
  _RAND_2752 = {1{`RANDOM}};
  amplifier_1_1_data_244 = _RAND_2752[7:0];
  _RAND_2753 = {1{`RANDOM}};
  amplifier_1_1_data_245 = _RAND_2753[7:0];
  _RAND_2754 = {1{`RANDOM}};
  amplifier_1_1_data_246 = _RAND_2754[7:0];
  _RAND_2755 = {1{`RANDOM}};
  amplifier_1_1_data_247 = _RAND_2755[7:0];
  _RAND_2756 = {1{`RANDOM}};
  amplifier_1_1_data_248 = _RAND_2756[7:0];
  _RAND_2757 = {1{`RANDOM}};
  amplifier_1_1_data_249 = _RAND_2757[7:0];
  _RAND_2758 = {1{`RANDOM}};
  amplifier_1_1_data_250 = _RAND_2758[7:0];
  _RAND_2759 = {1{`RANDOM}};
  amplifier_1_1_data_251 = _RAND_2759[7:0];
  _RAND_2760 = {1{`RANDOM}};
  amplifier_1_1_data_252 = _RAND_2760[7:0];
  _RAND_2761 = {1{`RANDOM}};
  amplifier_1_1_data_253 = _RAND_2761[7:0];
  _RAND_2762 = {1{`RANDOM}};
  amplifier_1_1_data_254 = _RAND_2762[7:0];
  _RAND_2763 = {1{`RANDOM}};
  amplifier_1_1_data_255 = _RAND_2763[7:0];
  _RAND_2764 = {1{`RANDOM}};
  amplifier_1_1_header_0 = _RAND_2764[15:0];
  _RAND_2765 = {1{`RANDOM}};
  amplifier_1_1_header_1 = _RAND_2765[15:0];
  _RAND_2766 = {1{`RANDOM}};
  amplifier_1_1_header_2 = _RAND_2766[15:0];
  _RAND_2767 = {1{`RANDOM}};
  amplifier_1_1_header_3 = _RAND_2767[15:0];
  _RAND_2768 = {1{`RANDOM}};
  amplifier_1_1_header_4 = _RAND_2768[15:0];
  _RAND_2769 = {1{`RANDOM}};
  amplifier_1_1_header_5 = _RAND_2769[15:0];
  _RAND_2770 = {1{`RANDOM}};
  amplifier_1_1_header_6 = _RAND_2770[15:0];
  _RAND_2771 = {1{`RANDOM}};
  amplifier_1_1_header_7 = _RAND_2771[15:0];
  _RAND_2772 = {1{`RANDOM}};
  amplifier_1_1_header_8 = _RAND_2772[15:0];
  _RAND_2773 = {1{`RANDOM}};
  amplifier_1_1_header_9 = _RAND_2773[15:0];
  _RAND_2774 = {1{`RANDOM}};
  amplifier_1_1_header_10 = _RAND_2774[15:0];
  _RAND_2775 = {1{`RANDOM}};
  amplifier_1_1_header_11 = _RAND_2775[15:0];
  _RAND_2776 = {1{`RANDOM}};
  amplifier_1_1_header_12 = _RAND_2776[15:0];
  _RAND_2777 = {1{`RANDOM}};
  amplifier_1_1_header_13 = _RAND_2777[15:0];
  _RAND_2778 = {1{`RANDOM}};
  amplifier_1_1_header_14 = _RAND_2778[15:0];
  _RAND_2779 = {1{`RANDOM}};
  amplifier_1_1_header_15 = _RAND_2779[15:0];
  _RAND_2780 = {1{`RANDOM}};
  amplifier_1_1_parse_current_state = _RAND_2780[7:0];
  _RAND_2781 = {1{`RANDOM}};
  amplifier_1_1_parse_current_offset = _RAND_2781[7:0];
  _RAND_2782 = {1{`RANDOM}};
  amplifier_1_1_parse_transition_field = _RAND_2782[15:0];
  _RAND_2783 = {1{`RANDOM}};
  amplifier_1_1_next_processor_id = _RAND_2783[1:0];
  _RAND_2784 = {1{`RANDOM}};
  amplifier_1_1_next_config_id = _RAND_2784[0:0];
  _RAND_2785 = {1{`RANDOM}};
  amplifier_1_1_is_valid_processor = _RAND_2785[0:0];
  _RAND_2786 = {1{`RANDOM}};
  amplifier_1_2_data_0 = _RAND_2786[7:0];
  _RAND_2787 = {1{`RANDOM}};
  amplifier_1_2_data_1 = _RAND_2787[7:0];
  _RAND_2788 = {1{`RANDOM}};
  amplifier_1_2_data_2 = _RAND_2788[7:0];
  _RAND_2789 = {1{`RANDOM}};
  amplifier_1_2_data_3 = _RAND_2789[7:0];
  _RAND_2790 = {1{`RANDOM}};
  amplifier_1_2_data_4 = _RAND_2790[7:0];
  _RAND_2791 = {1{`RANDOM}};
  amplifier_1_2_data_5 = _RAND_2791[7:0];
  _RAND_2792 = {1{`RANDOM}};
  amplifier_1_2_data_6 = _RAND_2792[7:0];
  _RAND_2793 = {1{`RANDOM}};
  amplifier_1_2_data_7 = _RAND_2793[7:0];
  _RAND_2794 = {1{`RANDOM}};
  amplifier_1_2_data_8 = _RAND_2794[7:0];
  _RAND_2795 = {1{`RANDOM}};
  amplifier_1_2_data_9 = _RAND_2795[7:0];
  _RAND_2796 = {1{`RANDOM}};
  amplifier_1_2_data_10 = _RAND_2796[7:0];
  _RAND_2797 = {1{`RANDOM}};
  amplifier_1_2_data_11 = _RAND_2797[7:0];
  _RAND_2798 = {1{`RANDOM}};
  amplifier_1_2_data_12 = _RAND_2798[7:0];
  _RAND_2799 = {1{`RANDOM}};
  amplifier_1_2_data_13 = _RAND_2799[7:0];
  _RAND_2800 = {1{`RANDOM}};
  amplifier_1_2_data_14 = _RAND_2800[7:0];
  _RAND_2801 = {1{`RANDOM}};
  amplifier_1_2_data_15 = _RAND_2801[7:0];
  _RAND_2802 = {1{`RANDOM}};
  amplifier_1_2_data_16 = _RAND_2802[7:0];
  _RAND_2803 = {1{`RANDOM}};
  amplifier_1_2_data_17 = _RAND_2803[7:0];
  _RAND_2804 = {1{`RANDOM}};
  amplifier_1_2_data_18 = _RAND_2804[7:0];
  _RAND_2805 = {1{`RANDOM}};
  amplifier_1_2_data_19 = _RAND_2805[7:0];
  _RAND_2806 = {1{`RANDOM}};
  amplifier_1_2_data_20 = _RAND_2806[7:0];
  _RAND_2807 = {1{`RANDOM}};
  amplifier_1_2_data_21 = _RAND_2807[7:0];
  _RAND_2808 = {1{`RANDOM}};
  amplifier_1_2_data_22 = _RAND_2808[7:0];
  _RAND_2809 = {1{`RANDOM}};
  amplifier_1_2_data_23 = _RAND_2809[7:0];
  _RAND_2810 = {1{`RANDOM}};
  amplifier_1_2_data_24 = _RAND_2810[7:0];
  _RAND_2811 = {1{`RANDOM}};
  amplifier_1_2_data_25 = _RAND_2811[7:0];
  _RAND_2812 = {1{`RANDOM}};
  amplifier_1_2_data_26 = _RAND_2812[7:0];
  _RAND_2813 = {1{`RANDOM}};
  amplifier_1_2_data_27 = _RAND_2813[7:0];
  _RAND_2814 = {1{`RANDOM}};
  amplifier_1_2_data_28 = _RAND_2814[7:0];
  _RAND_2815 = {1{`RANDOM}};
  amplifier_1_2_data_29 = _RAND_2815[7:0];
  _RAND_2816 = {1{`RANDOM}};
  amplifier_1_2_data_30 = _RAND_2816[7:0];
  _RAND_2817 = {1{`RANDOM}};
  amplifier_1_2_data_31 = _RAND_2817[7:0];
  _RAND_2818 = {1{`RANDOM}};
  amplifier_1_2_data_32 = _RAND_2818[7:0];
  _RAND_2819 = {1{`RANDOM}};
  amplifier_1_2_data_33 = _RAND_2819[7:0];
  _RAND_2820 = {1{`RANDOM}};
  amplifier_1_2_data_34 = _RAND_2820[7:0];
  _RAND_2821 = {1{`RANDOM}};
  amplifier_1_2_data_35 = _RAND_2821[7:0];
  _RAND_2822 = {1{`RANDOM}};
  amplifier_1_2_data_36 = _RAND_2822[7:0];
  _RAND_2823 = {1{`RANDOM}};
  amplifier_1_2_data_37 = _RAND_2823[7:0];
  _RAND_2824 = {1{`RANDOM}};
  amplifier_1_2_data_38 = _RAND_2824[7:0];
  _RAND_2825 = {1{`RANDOM}};
  amplifier_1_2_data_39 = _RAND_2825[7:0];
  _RAND_2826 = {1{`RANDOM}};
  amplifier_1_2_data_40 = _RAND_2826[7:0];
  _RAND_2827 = {1{`RANDOM}};
  amplifier_1_2_data_41 = _RAND_2827[7:0];
  _RAND_2828 = {1{`RANDOM}};
  amplifier_1_2_data_42 = _RAND_2828[7:0];
  _RAND_2829 = {1{`RANDOM}};
  amplifier_1_2_data_43 = _RAND_2829[7:0];
  _RAND_2830 = {1{`RANDOM}};
  amplifier_1_2_data_44 = _RAND_2830[7:0];
  _RAND_2831 = {1{`RANDOM}};
  amplifier_1_2_data_45 = _RAND_2831[7:0];
  _RAND_2832 = {1{`RANDOM}};
  amplifier_1_2_data_46 = _RAND_2832[7:0];
  _RAND_2833 = {1{`RANDOM}};
  amplifier_1_2_data_47 = _RAND_2833[7:0];
  _RAND_2834 = {1{`RANDOM}};
  amplifier_1_2_data_48 = _RAND_2834[7:0];
  _RAND_2835 = {1{`RANDOM}};
  amplifier_1_2_data_49 = _RAND_2835[7:0];
  _RAND_2836 = {1{`RANDOM}};
  amplifier_1_2_data_50 = _RAND_2836[7:0];
  _RAND_2837 = {1{`RANDOM}};
  amplifier_1_2_data_51 = _RAND_2837[7:0];
  _RAND_2838 = {1{`RANDOM}};
  amplifier_1_2_data_52 = _RAND_2838[7:0];
  _RAND_2839 = {1{`RANDOM}};
  amplifier_1_2_data_53 = _RAND_2839[7:0];
  _RAND_2840 = {1{`RANDOM}};
  amplifier_1_2_data_54 = _RAND_2840[7:0];
  _RAND_2841 = {1{`RANDOM}};
  amplifier_1_2_data_55 = _RAND_2841[7:0];
  _RAND_2842 = {1{`RANDOM}};
  amplifier_1_2_data_56 = _RAND_2842[7:0];
  _RAND_2843 = {1{`RANDOM}};
  amplifier_1_2_data_57 = _RAND_2843[7:0];
  _RAND_2844 = {1{`RANDOM}};
  amplifier_1_2_data_58 = _RAND_2844[7:0];
  _RAND_2845 = {1{`RANDOM}};
  amplifier_1_2_data_59 = _RAND_2845[7:0];
  _RAND_2846 = {1{`RANDOM}};
  amplifier_1_2_data_60 = _RAND_2846[7:0];
  _RAND_2847 = {1{`RANDOM}};
  amplifier_1_2_data_61 = _RAND_2847[7:0];
  _RAND_2848 = {1{`RANDOM}};
  amplifier_1_2_data_62 = _RAND_2848[7:0];
  _RAND_2849 = {1{`RANDOM}};
  amplifier_1_2_data_63 = _RAND_2849[7:0];
  _RAND_2850 = {1{`RANDOM}};
  amplifier_1_2_data_64 = _RAND_2850[7:0];
  _RAND_2851 = {1{`RANDOM}};
  amplifier_1_2_data_65 = _RAND_2851[7:0];
  _RAND_2852 = {1{`RANDOM}};
  amplifier_1_2_data_66 = _RAND_2852[7:0];
  _RAND_2853 = {1{`RANDOM}};
  amplifier_1_2_data_67 = _RAND_2853[7:0];
  _RAND_2854 = {1{`RANDOM}};
  amplifier_1_2_data_68 = _RAND_2854[7:0];
  _RAND_2855 = {1{`RANDOM}};
  amplifier_1_2_data_69 = _RAND_2855[7:0];
  _RAND_2856 = {1{`RANDOM}};
  amplifier_1_2_data_70 = _RAND_2856[7:0];
  _RAND_2857 = {1{`RANDOM}};
  amplifier_1_2_data_71 = _RAND_2857[7:0];
  _RAND_2858 = {1{`RANDOM}};
  amplifier_1_2_data_72 = _RAND_2858[7:0];
  _RAND_2859 = {1{`RANDOM}};
  amplifier_1_2_data_73 = _RAND_2859[7:0];
  _RAND_2860 = {1{`RANDOM}};
  amplifier_1_2_data_74 = _RAND_2860[7:0];
  _RAND_2861 = {1{`RANDOM}};
  amplifier_1_2_data_75 = _RAND_2861[7:0];
  _RAND_2862 = {1{`RANDOM}};
  amplifier_1_2_data_76 = _RAND_2862[7:0];
  _RAND_2863 = {1{`RANDOM}};
  amplifier_1_2_data_77 = _RAND_2863[7:0];
  _RAND_2864 = {1{`RANDOM}};
  amplifier_1_2_data_78 = _RAND_2864[7:0];
  _RAND_2865 = {1{`RANDOM}};
  amplifier_1_2_data_79 = _RAND_2865[7:0];
  _RAND_2866 = {1{`RANDOM}};
  amplifier_1_2_data_80 = _RAND_2866[7:0];
  _RAND_2867 = {1{`RANDOM}};
  amplifier_1_2_data_81 = _RAND_2867[7:0];
  _RAND_2868 = {1{`RANDOM}};
  amplifier_1_2_data_82 = _RAND_2868[7:0];
  _RAND_2869 = {1{`RANDOM}};
  amplifier_1_2_data_83 = _RAND_2869[7:0];
  _RAND_2870 = {1{`RANDOM}};
  amplifier_1_2_data_84 = _RAND_2870[7:0];
  _RAND_2871 = {1{`RANDOM}};
  amplifier_1_2_data_85 = _RAND_2871[7:0];
  _RAND_2872 = {1{`RANDOM}};
  amplifier_1_2_data_86 = _RAND_2872[7:0];
  _RAND_2873 = {1{`RANDOM}};
  amplifier_1_2_data_87 = _RAND_2873[7:0];
  _RAND_2874 = {1{`RANDOM}};
  amplifier_1_2_data_88 = _RAND_2874[7:0];
  _RAND_2875 = {1{`RANDOM}};
  amplifier_1_2_data_89 = _RAND_2875[7:0];
  _RAND_2876 = {1{`RANDOM}};
  amplifier_1_2_data_90 = _RAND_2876[7:0];
  _RAND_2877 = {1{`RANDOM}};
  amplifier_1_2_data_91 = _RAND_2877[7:0];
  _RAND_2878 = {1{`RANDOM}};
  amplifier_1_2_data_92 = _RAND_2878[7:0];
  _RAND_2879 = {1{`RANDOM}};
  amplifier_1_2_data_93 = _RAND_2879[7:0];
  _RAND_2880 = {1{`RANDOM}};
  amplifier_1_2_data_94 = _RAND_2880[7:0];
  _RAND_2881 = {1{`RANDOM}};
  amplifier_1_2_data_95 = _RAND_2881[7:0];
  _RAND_2882 = {1{`RANDOM}};
  amplifier_1_2_data_96 = _RAND_2882[7:0];
  _RAND_2883 = {1{`RANDOM}};
  amplifier_1_2_data_97 = _RAND_2883[7:0];
  _RAND_2884 = {1{`RANDOM}};
  amplifier_1_2_data_98 = _RAND_2884[7:0];
  _RAND_2885 = {1{`RANDOM}};
  amplifier_1_2_data_99 = _RAND_2885[7:0];
  _RAND_2886 = {1{`RANDOM}};
  amplifier_1_2_data_100 = _RAND_2886[7:0];
  _RAND_2887 = {1{`RANDOM}};
  amplifier_1_2_data_101 = _RAND_2887[7:0];
  _RAND_2888 = {1{`RANDOM}};
  amplifier_1_2_data_102 = _RAND_2888[7:0];
  _RAND_2889 = {1{`RANDOM}};
  amplifier_1_2_data_103 = _RAND_2889[7:0];
  _RAND_2890 = {1{`RANDOM}};
  amplifier_1_2_data_104 = _RAND_2890[7:0];
  _RAND_2891 = {1{`RANDOM}};
  amplifier_1_2_data_105 = _RAND_2891[7:0];
  _RAND_2892 = {1{`RANDOM}};
  amplifier_1_2_data_106 = _RAND_2892[7:0];
  _RAND_2893 = {1{`RANDOM}};
  amplifier_1_2_data_107 = _RAND_2893[7:0];
  _RAND_2894 = {1{`RANDOM}};
  amplifier_1_2_data_108 = _RAND_2894[7:0];
  _RAND_2895 = {1{`RANDOM}};
  amplifier_1_2_data_109 = _RAND_2895[7:0];
  _RAND_2896 = {1{`RANDOM}};
  amplifier_1_2_data_110 = _RAND_2896[7:0];
  _RAND_2897 = {1{`RANDOM}};
  amplifier_1_2_data_111 = _RAND_2897[7:0];
  _RAND_2898 = {1{`RANDOM}};
  amplifier_1_2_data_112 = _RAND_2898[7:0];
  _RAND_2899 = {1{`RANDOM}};
  amplifier_1_2_data_113 = _RAND_2899[7:0];
  _RAND_2900 = {1{`RANDOM}};
  amplifier_1_2_data_114 = _RAND_2900[7:0];
  _RAND_2901 = {1{`RANDOM}};
  amplifier_1_2_data_115 = _RAND_2901[7:0];
  _RAND_2902 = {1{`RANDOM}};
  amplifier_1_2_data_116 = _RAND_2902[7:0];
  _RAND_2903 = {1{`RANDOM}};
  amplifier_1_2_data_117 = _RAND_2903[7:0];
  _RAND_2904 = {1{`RANDOM}};
  amplifier_1_2_data_118 = _RAND_2904[7:0];
  _RAND_2905 = {1{`RANDOM}};
  amplifier_1_2_data_119 = _RAND_2905[7:0];
  _RAND_2906 = {1{`RANDOM}};
  amplifier_1_2_data_120 = _RAND_2906[7:0];
  _RAND_2907 = {1{`RANDOM}};
  amplifier_1_2_data_121 = _RAND_2907[7:0];
  _RAND_2908 = {1{`RANDOM}};
  amplifier_1_2_data_122 = _RAND_2908[7:0];
  _RAND_2909 = {1{`RANDOM}};
  amplifier_1_2_data_123 = _RAND_2909[7:0];
  _RAND_2910 = {1{`RANDOM}};
  amplifier_1_2_data_124 = _RAND_2910[7:0];
  _RAND_2911 = {1{`RANDOM}};
  amplifier_1_2_data_125 = _RAND_2911[7:0];
  _RAND_2912 = {1{`RANDOM}};
  amplifier_1_2_data_126 = _RAND_2912[7:0];
  _RAND_2913 = {1{`RANDOM}};
  amplifier_1_2_data_127 = _RAND_2913[7:0];
  _RAND_2914 = {1{`RANDOM}};
  amplifier_1_2_data_128 = _RAND_2914[7:0];
  _RAND_2915 = {1{`RANDOM}};
  amplifier_1_2_data_129 = _RAND_2915[7:0];
  _RAND_2916 = {1{`RANDOM}};
  amplifier_1_2_data_130 = _RAND_2916[7:0];
  _RAND_2917 = {1{`RANDOM}};
  amplifier_1_2_data_131 = _RAND_2917[7:0];
  _RAND_2918 = {1{`RANDOM}};
  amplifier_1_2_data_132 = _RAND_2918[7:0];
  _RAND_2919 = {1{`RANDOM}};
  amplifier_1_2_data_133 = _RAND_2919[7:0];
  _RAND_2920 = {1{`RANDOM}};
  amplifier_1_2_data_134 = _RAND_2920[7:0];
  _RAND_2921 = {1{`RANDOM}};
  amplifier_1_2_data_135 = _RAND_2921[7:0];
  _RAND_2922 = {1{`RANDOM}};
  amplifier_1_2_data_136 = _RAND_2922[7:0];
  _RAND_2923 = {1{`RANDOM}};
  amplifier_1_2_data_137 = _RAND_2923[7:0];
  _RAND_2924 = {1{`RANDOM}};
  amplifier_1_2_data_138 = _RAND_2924[7:0];
  _RAND_2925 = {1{`RANDOM}};
  amplifier_1_2_data_139 = _RAND_2925[7:0];
  _RAND_2926 = {1{`RANDOM}};
  amplifier_1_2_data_140 = _RAND_2926[7:0];
  _RAND_2927 = {1{`RANDOM}};
  amplifier_1_2_data_141 = _RAND_2927[7:0];
  _RAND_2928 = {1{`RANDOM}};
  amplifier_1_2_data_142 = _RAND_2928[7:0];
  _RAND_2929 = {1{`RANDOM}};
  amplifier_1_2_data_143 = _RAND_2929[7:0];
  _RAND_2930 = {1{`RANDOM}};
  amplifier_1_2_data_144 = _RAND_2930[7:0];
  _RAND_2931 = {1{`RANDOM}};
  amplifier_1_2_data_145 = _RAND_2931[7:0];
  _RAND_2932 = {1{`RANDOM}};
  amplifier_1_2_data_146 = _RAND_2932[7:0];
  _RAND_2933 = {1{`RANDOM}};
  amplifier_1_2_data_147 = _RAND_2933[7:0];
  _RAND_2934 = {1{`RANDOM}};
  amplifier_1_2_data_148 = _RAND_2934[7:0];
  _RAND_2935 = {1{`RANDOM}};
  amplifier_1_2_data_149 = _RAND_2935[7:0];
  _RAND_2936 = {1{`RANDOM}};
  amplifier_1_2_data_150 = _RAND_2936[7:0];
  _RAND_2937 = {1{`RANDOM}};
  amplifier_1_2_data_151 = _RAND_2937[7:0];
  _RAND_2938 = {1{`RANDOM}};
  amplifier_1_2_data_152 = _RAND_2938[7:0];
  _RAND_2939 = {1{`RANDOM}};
  amplifier_1_2_data_153 = _RAND_2939[7:0];
  _RAND_2940 = {1{`RANDOM}};
  amplifier_1_2_data_154 = _RAND_2940[7:0];
  _RAND_2941 = {1{`RANDOM}};
  amplifier_1_2_data_155 = _RAND_2941[7:0];
  _RAND_2942 = {1{`RANDOM}};
  amplifier_1_2_data_156 = _RAND_2942[7:0];
  _RAND_2943 = {1{`RANDOM}};
  amplifier_1_2_data_157 = _RAND_2943[7:0];
  _RAND_2944 = {1{`RANDOM}};
  amplifier_1_2_data_158 = _RAND_2944[7:0];
  _RAND_2945 = {1{`RANDOM}};
  amplifier_1_2_data_159 = _RAND_2945[7:0];
  _RAND_2946 = {1{`RANDOM}};
  amplifier_1_2_data_160 = _RAND_2946[7:0];
  _RAND_2947 = {1{`RANDOM}};
  amplifier_1_2_data_161 = _RAND_2947[7:0];
  _RAND_2948 = {1{`RANDOM}};
  amplifier_1_2_data_162 = _RAND_2948[7:0];
  _RAND_2949 = {1{`RANDOM}};
  amplifier_1_2_data_163 = _RAND_2949[7:0];
  _RAND_2950 = {1{`RANDOM}};
  amplifier_1_2_data_164 = _RAND_2950[7:0];
  _RAND_2951 = {1{`RANDOM}};
  amplifier_1_2_data_165 = _RAND_2951[7:0];
  _RAND_2952 = {1{`RANDOM}};
  amplifier_1_2_data_166 = _RAND_2952[7:0];
  _RAND_2953 = {1{`RANDOM}};
  amplifier_1_2_data_167 = _RAND_2953[7:0];
  _RAND_2954 = {1{`RANDOM}};
  amplifier_1_2_data_168 = _RAND_2954[7:0];
  _RAND_2955 = {1{`RANDOM}};
  amplifier_1_2_data_169 = _RAND_2955[7:0];
  _RAND_2956 = {1{`RANDOM}};
  amplifier_1_2_data_170 = _RAND_2956[7:0];
  _RAND_2957 = {1{`RANDOM}};
  amplifier_1_2_data_171 = _RAND_2957[7:0];
  _RAND_2958 = {1{`RANDOM}};
  amplifier_1_2_data_172 = _RAND_2958[7:0];
  _RAND_2959 = {1{`RANDOM}};
  amplifier_1_2_data_173 = _RAND_2959[7:0];
  _RAND_2960 = {1{`RANDOM}};
  amplifier_1_2_data_174 = _RAND_2960[7:0];
  _RAND_2961 = {1{`RANDOM}};
  amplifier_1_2_data_175 = _RAND_2961[7:0];
  _RAND_2962 = {1{`RANDOM}};
  amplifier_1_2_data_176 = _RAND_2962[7:0];
  _RAND_2963 = {1{`RANDOM}};
  amplifier_1_2_data_177 = _RAND_2963[7:0];
  _RAND_2964 = {1{`RANDOM}};
  amplifier_1_2_data_178 = _RAND_2964[7:0];
  _RAND_2965 = {1{`RANDOM}};
  amplifier_1_2_data_179 = _RAND_2965[7:0];
  _RAND_2966 = {1{`RANDOM}};
  amplifier_1_2_data_180 = _RAND_2966[7:0];
  _RAND_2967 = {1{`RANDOM}};
  amplifier_1_2_data_181 = _RAND_2967[7:0];
  _RAND_2968 = {1{`RANDOM}};
  amplifier_1_2_data_182 = _RAND_2968[7:0];
  _RAND_2969 = {1{`RANDOM}};
  amplifier_1_2_data_183 = _RAND_2969[7:0];
  _RAND_2970 = {1{`RANDOM}};
  amplifier_1_2_data_184 = _RAND_2970[7:0];
  _RAND_2971 = {1{`RANDOM}};
  amplifier_1_2_data_185 = _RAND_2971[7:0];
  _RAND_2972 = {1{`RANDOM}};
  amplifier_1_2_data_186 = _RAND_2972[7:0];
  _RAND_2973 = {1{`RANDOM}};
  amplifier_1_2_data_187 = _RAND_2973[7:0];
  _RAND_2974 = {1{`RANDOM}};
  amplifier_1_2_data_188 = _RAND_2974[7:0];
  _RAND_2975 = {1{`RANDOM}};
  amplifier_1_2_data_189 = _RAND_2975[7:0];
  _RAND_2976 = {1{`RANDOM}};
  amplifier_1_2_data_190 = _RAND_2976[7:0];
  _RAND_2977 = {1{`RANDOM}};
  amplifier_1_2_data_191 = _RAND_2977[7:0];
  _RAND_2978 = {1{`RANDOM}};
  amplifier_1_2_data_192 = _RAND_2978[7:0];
  _RAND_2979 = {1{`RANDOM}};
  amplifier_1_2_data_193 = _RAND_2979[7:0];
  _RAND_2980 = {1{`RANDOM}};
  amplifier_1_2_data_194 = _RAND_2980[7:0];
  _RAND_2981 = {1{`RANDOM}};
  amplifier_1_2_data_195 = _RAND_2981[7:0];
  _RAND_2982 = {1{`RANDOM}};
  amplifier_1_2_data_196 = _RAND_2982[7:0];
  _RAND_2983 = {1{`RANDOM}};
  amplifier_1_2_data_197 = _RAND_2983[7:0];
  _RAND_2984 = {1{`RANDOM}};
  amplifier_1_2_data_198 = _RAND_2984[7:0];
  _RAND_2985 = {1{`RANDOM}};
  amplifier_1_2_data_199 = _RAND_2985[7:0];
  _RAND_2986 = {1{`RANDOM}};
  amplifier_1_2_data_200 = _RAND_2986[7:0];
  _RAND_2987 = {1{`RANDOM}};
  amplifier_1_2_data_201 = _RAND_2987[7:0];
  _RAND_2988 = {1{`RANDOM}};
  amplifier_1_2_data_202 = _RAND_2988[7:0];
  _RAND_2989 = {1{`RANDOM}};
  amplifier_1_2_data_203 = _RAND_2989[7:0];
  _RAND_2990 = {1{`RANDOM}};
  amplifier_1_2_data_204 = _RAND_2990[7:0];
  _RAND_2991 = {1{`RANDOM}};
  amplifier_1_2_data_205 = _RAND_2991[7:0];
  _RAND_2992 = {1{`RANDOM}};
  amplifier_1_2_data_206 = _RAND_2992[7:0];
  _RAND_2993 = {1{`RANDOM}};
  amplifier_1_2_data_207 = _RAND_2993[7:0];
  _RAND_2994 = {1{`RANDOM}};
  amplifier_1_2_data_208 = _RAND_2994[7:0];
  _RAND_2995 = {1{`RANDOM}};
  amplifier_1_2_data_209 = _RAND_2995[7:0];
  _RAND_2996 = {1{`RANDOM}};
  amplifier_1_2_data_210 = _RAND_2996[7:0];
  _RAND_2997 = {1{`RANDOM}};
  amplifier_1_2_data_211 = _RAND_2997[7:0];
  _RAND_2998 = {1{`RANDOM}};
  amplifier_1_2_data_212 = _RAND_2998[7:0];
  _RAND_2999 = {1{`RANDOM}};
  amplifier_1_2_data_213 = _RAND_2999[7:0];
  _RAND_3000 = {1{`RANDOM}};
  amplifier_1_2_data_214 = _RAND_3000[7:0];
  _RAND_3001 = {1{`RANDOM}};
  amplifier_1_2_data_215 = _RAND_3001[7:0];
  _RAND_3002 = {1{`RANDOM}};
  amplifier_1_2_data_216 = _RAND_3002[7:0];
  _RAND_3003 = {1{`RANDOM}};
  amplifier_1_2_data_217 = _RAND_3003[7:0];
  _RAND_3004 = {1{`RANDOM}};
  amplifier_1_2_data_218 = _RAND_3004[7:0];
  _RAND_3005 = {1{`RANDOM}};
  amplifier_1_2_data_219 = _RAND_3005[7:0];
  _RAND_3006 = {1{`RANDOM}};
  amplifier_1_2_data_220 = _RAND_3006[7:0];
  _RAND_3007 = {1{`RANDOM}};
  amplifier_1_2_data_221 = _RAND_3007[7:0];
  _RAND_3008 = {1{`RANDOM}};
  amplifier_1_2_data_222 = _RAND_3008[7:0];
  _RAND_3009 = {1{`RANDOM}};
  amplifier_1_2_data_223 = _RAND_3009[7:0];
  _RAND_3010 = {1{`RANDOM}};
  amplifier_1_2_data_224 = _RAND_3010[7:0];
  _RAND_3011 = {1{`RANDOM}};
  amplifier_1_2_data_225 = _RAND_3011[7:0];
  _RAND_3012 = {1{`RANDOM}};
  amplifier_1_2_data_226 = _RAND_3012[7:0];
  _RAND_3013 = {1{`RANDOM}};
  amplifier_1_2_data_227 = _RAND_3013[7:0];
  _RAND_3014 = {1{`RANDOM}};
  amplifier_1_2_data_228 = _RAND_3014[7:0];
  _RAND_3015 = {1{`RANDOM}};
  amplifier_1_2_data_229 = _RAND_3015[7:0];
  _RAND_3016 = {1{`RANDOM}};
  amplifier_1_2_data_230 = _RAND_3016[7:0];
  _RAND_3017 = {1{`RANDOM}};
  amplifier_1_2_data_231 = _RAND_3017[7:0];
  _RAND_3018 = {1{`RANDOM}};
  amplifier_1_2_data_232 = _RAND_3018[7:0];
  _RAND_3019 = {1{`RANDOM}};
  amplifier_1_2_data_233 = _RAND_3019[7:0];
  _RAND_3020 = {1{`RANDOM}};
  amplifier_1_2_data_234 = _RAND_3020[7:0];
  _RAND_3021 = {1{`RANDOM}};
  amplifier_1_2_data_235 = _RAND_3021[7:0];
  _RAND_3022 = {1{`RANDOM}};
  amplifier_1_2_data_236 = _RAND_3022[7:0];
  _RAND_3023 = {1{`RANDOM}};
  amplifier_1_2_data_237 = _RAND_3023[7:0];
  _RAND_3024 = {1{`RANDOM}};
  amplifier_1_2_data_238 = _RAND_3024[7:0];
  _RAND_3025 = {1{`RANDOM}};
  amplifier_1_2_data_239 = _RAND_3025[7:0];
  _RAND_3026 = {1{`RANDOM}};
  amplifier_1_2_data_240 = _RAND_3026[7:0];
  _RAND_3027 = {1{`RANDOM}};
  amplifier_1_2_data_241 = _RAND_3027[7:0];
  _RAND_3028 = {1{`RANDOM}};
  amplifier_1_2_data_242 = _RAND_3028[7:0];
  _RAND_3029 = {1{`RANDOM}};
  amplifier_1_2_data_243 = _RAND_3029[7:0];
  _RAND_3030 = {1{`RANDOM}};
  amplifier_1_2_data_244 = _RAND_3030[7:0];
  _RAND_3031 = {1{`RANDOM}};
  amplifier_1_2_data_245 = _RAND_3031[7:0];
  _RAND_3032 = {1{`RANDOM}};
  amplifier_1_2_data_246 = _RAND_3032[7:0];
  _RAND_3033 = {1{`RANDOM}};
  amplifier_1_2_data_247 = _RAND_3033[7:0];
  _RAND_3034 = {1{`RANDOM}};
  amplifier_1_2_data_248 = _RAND_3034[7:0];
  _RAND_3035 = {1{`RANDOM}};
  amplifier_1_2_data_249 = _RAND_3035[7:0];
  _RAND_3036 = {1{`RANDOM}};
  amplifier_1_2_data_250 = _RAND_3036[7:0];
  _RAND_3037 = {1{`RANDOM}};
  amplifier_1_2_data_251 = _RAND_3037[7:0];
  _RAND_3038 = {1{`RANDOM}};
  amplifier_1_2_data_252 = _RAND_3038[7:0];
  _RAND_3039 = {1{`RANDOM}};
  amplifier_1_2_data_253 = _RAND_3039[7:0];
  _RAND_3040 = {1{`RANDOM}};
  amplifier_1_2_data_254 = _RAND_3040[7:0];
  _RAND_3041 = {1{`RANDOM}};
  amplifier_1_2_data_255 = _RAND_3041[7:0];
  _RAND_3042 = {1{`RANDOM}};
  amplifier_1_2_header_0 = _RAND_3042[15:0];
  _RAND_3043 = {1{`RANDOM}};
  amplifier_1_2_header_1 = _RAND_3043[15:0];
  _RAND_3044 = {1{`RANDOM}};
  amplifier_1_2_header_2 = _RAND_3044[15:0];
  _RAND_3045 = {1{`RANDOM}};
  amplifier_1_2_header_3 = _RAND_3045[15:0];
  _RAND_3046 = {1{`RANDOM}};
  amplifier_1_2_header_4 = _RAND_3046[15:0];
  _RAND_3047 = {1{`RANDOM}};
  amplifier_1_2_header_5 = _RAND_3047[15:0];
  _RAND_3048 = {1{`RANDOM}};
  amplifier_1_2_header_6 = _RAND_3048[15:0];
  _RAND_3049 = {1{`RANDOM}};
  amplifier_1_2_header_7 = _RAND_3049[15:0];
  _RAND_3050 = {1{`RANDOM}};
  amplifier_1_2_header_8 = _RAND_3050[15:0];
  _RAND_3051 = {1{`RANDOM}};
  amplifier_1_2_header_9 = _RAND_3051[15:0];
  _RAND_3052 = {1{`RANDOM}};
  amplifier_1_2_header_10 = _RAND_3052[15:0];
  _RAND_3053 = {1{`RANDOM}};
  amplifier_1_2_header_11 = _RAND_3053[15:0];
  _RAND_3054 = {1{`RANDOM}};
  amplifier_1_2_header_12 = _RAND_3054[15:0];
  _RAND_3055 = {1{`RANDOM}};
  amplifier_1_2_header_13 = _RAND_3055[15:0];
  _RAND_3056 = {1{`RANDOM}};
  amplifier_1_2_header_14 = _RAND_3056[15:0];
  _RAND_3057 = {1{`RANDOM}};
  amplifier_1_2_header_15 = _RAND_3057[15:0];
  _RAND_3058 = {1{`RANDOM}};
  amplifier_1_2_parse_current_state = _RAND_3058[7:0];
  _RAND_3059 = {1{`RANDOM}};
  amplifier_1_2_parse_current_offset = _RAND_3059[7:0];
  _RAND_3060 = {1{`RANDOM}};
  amplifier_1_2_parse_transition_field = _RAND_3060[15:0];
  _RAND_3061 = {1{`RANDOM}};
  amplifier_1_2_next_processor_id = _RAND_3061[1:0];
  _RAND_3062 = {1{`RANDOM}};
  amplifier_1_2_next_config_id = _RAND_3062[0:0];
  _RAND_3063 = {1{`RANDOM}};
  amplifier_1_2_is_valid_processor = _RAND_3063[0:0];
  _RAND_3064 = {1{`RANDOM}};
  amplifier_1_3_data_0 = _RAND_3064[7:0];
  _RAND_3065 = {1{`RANDOM}};
  amplifier_1_3_data_1 = _RAND_3065[7:0];
  _RAND_3066 = {1{`RANDOM}};
  amplifier_1_3_data_2 = _RAND_3066[7:0];
  _RAND_3067 = {1{`RANDOM}};
  amplifier_1_3_data_3 = _RAND_3067[7:0];
  _RAND_3068 = {1{`RANDOM}};
  amplifier_1_3_data_4 = _RAND_3068[7:0];
  _RAND_3069 = {1{`RANDOM}};
  amplifier_1_3_data_5 = _RAND_3069[7:0];
  _RAND_3070 = {1{`RANDOM}};
  amplifier_1_3_data_6 = _RAND_3070[7:0];
  _RAND_3071 = {1{`RANDOM}};
  amplifier_1_3_data_7 = _RAND_3071[7:0];
  _RAND_3072 = {1{`RANDOM}};
  amplifier_1_3_data_8 = _RAND_3072[7:0];
  _RAND_3073 = {1{`RANDOM}};
  amplifier_1_3_data_9 = _RAND_3073[7:0];
  _RAND_3074 = {1{`RANDOM}};
  amplifier_1_3_data_10 = _RAND_3074[7:0];
  _RAND_3075 = {1{`RANDOM}};
  amplifier_1_3_data_11 = _RAND_3075[7:0];
  _RAND_3076 = {1{`RANDOM}};
  amplifier_1_3_data_12 = _RAND_3076[7:0];
  _RAND_3077 = {1{`RANDOM}};
  amplifier_1_3_data_13 = _RAND_3077[7:0];
  _RAND_3078 = {1{`RANDOM}};
  amplifier_1_3_data_14 = _RAND_3078[7:0];
  _RAND_3079 = {1{`RANDOM}};
  amplifier_1_3_data_15 = _RAND_3079[7:0];
  _RAND_3080 = {1{`RANDOM}};
  amplifier_1_3_data_16 = _RAND_3080[7:0];
  _RAND_3081 = {1{`RANDOM}};
  amplifier_1_3_data_17 = _RAND_3081[7:0];
  _RAND_3082 = {1{`RANDOM}};
  amplifier_1_3_data_18 = _RAND_3082[7:0];
  _RAND_3083 = {1{`RANDOM}};
  amplifier_1_3_data_19 = _RAND_3083[7:0];
  _RAND_3084 = {1{`RANDOM}};
  amplifier_1_3_data_20 = _RAND_3084[7:0];
  _RAND_3085 = {1{`RANDOM}};
  amplifier_1_3_data_21 = _RAND_3085[7:0];
  _RAND_3086 = {1{`RANDOM}};
  amplifier_1_3_data_22 = _RAND_3086[7:0];
  _RAND_3087 = {1{`RANDOM}};
  amplifier_1_3_data_23 = _RAND_3087[7:0];
  _RAND_3088 = {1{`RANDOM}};
  amplifier_1_3_data_24 = _RAND_3088[7:0];
  _RAND_3089 = {1{`RANDOM}};
  amplifier_1_3_data_25 = _RAND_3089[7:0];
  _RAND_3090 = {1{`RANDOM}};
  amplifier_1_3_data_26 = _RAND_3090[7:0];
  _RAND_3091 = {1{`RANDOM}};
  amplifier_1_3_data_27 = _RAND_3091[7:0];
  _RAND_3092 = {1{`RANDOM}};
  amplifier_1_3_data_28 = _RAND_3092[7:0];
  _RAND_3093 = {1{`RANDOM}};
  amplifier_1_3_data_29 = _RAND_3093[7:0];
  _RAND_3094 = {1{`RANDOM}};
  amplifier_1_3_data_30 = _RAND_3094[7:0];
  _RAND_3095 = {1{`RANDOM}};
  amplifier_1_3_data_31 = _RAND_3095[7:0];
  _RAND_3096 = {1{`RANDOM}};
  amplifier_1_3_data_32 = _RAND_3096[7:0];
  _RAND_3097 = {1{`RANDOM}};
  amplifier_1_3_data_33 = _RAND_3097[7:0];
  _RAND_3098 = {1{`RANDOM}};
  amplifier_1_3_data_34 = _RAND_3098[7:0];
  _RAND_3099 = {1{`RANDOM}};
  amplifier_1_3_data_35 = _RAND_3099[7:0];
  _RAND_3100 = {1{`RANDOM}};
  amplifier_1_3_data_36 = _RAND_3100[7:0];
  _RAND_3101 = {1{`RANDOM}};
  amplifier_1_3_data_37 = _RAND_3101[7:0];
  _RAND_3102 = {1{`RANDOM}};
  amplifier_1_3_data_38 = _RAND_3102[7:0];
  _RAND_3103 = {1{`RANDOM}};
  amplifier_1_3_data_39 = _RAND_3103[7:0];
  _RAND_3104 = {1{`RANDOM}};
  amplifier_1_3_data_40 = _RAND_3104[7:0];
  _RAND_3105 = {1{`RANDOM}};
  amplifier_1_3_data_41 = _RAND_3105[7:0];
  _RAND_3106 = {1{`RANDOM}};
  amplifier_1_3_data_42 = _RAND_3106[7:0];
  _RAND_3107 = {1{`RANDOM}};
  amplifier_1_3_data_43 = _RAND_3107[7:0];
  _RAND_3108 = {1{`RANDOM}};
  amplifier_1_3_data_44 = _RAND_3108[7:0];
  _RAND_3109 = {1{`RANDOM}};
  amplifier_1_3_data_45 = _RAND_3109[7:0];
  _RAND_3110 = {1{`RANDOM}};
  amplifier_1_3_data_46 = _RAND_3110[7:0];
  _RAND_3111 = {1{`RANDOM}};
  amplifier_1_3_data_47 = _RAND_3111[7:0];
  _RAND_3112 = {1{`RANDOM}};
  amplifier_1_3_data_48 = _RAND_3112[7:0];
  _RAND_3113 = {1{`RANDOM}};
  amplifier_1_3_data_49 = _RAND_3113[7:0];
  _RAND_3114 = {1{`RANDOM}};
  amplifier_1_3_data_50 = _RAND_3114[7:0];
  _RAND_3115 = {1{`RANDOM}};
  amplifier_1_3_data_51 = _RAND_3115[7:0];
  _RAND_3116 = {1{`RANDOM}};
  amplifier_1_3_data_52 = _RAND_3116[7:0];
  _RAND_3117 = {1{`RANDOM}};
  amplifier_1_3_data_53 = _RAND_3117[7:0];
  _RAND_3118 = {1{`RANDOM}};
  amplifier_1_3_data_54 = _RAND_3118[7:0];
  _RAND_3119 = {1{`RANDOM}};
  amplifier_1_3_data_55 = _RAND_3119[7:0];
  _RAND_3120 = {1{`RANDOM}};
  amplifier_1_3_data_56 = _RAND_3120[7:0];
  _RAND_3121 = {1{`RANDOM}};
  amplifier_1_3_data_57 = _RAND_3121[7:0];
  _RAND_3122 = {1{`RANDOM}};
  amplifier_1_3_data_58 = _RAND_3122[7:0];
  _RAND_3123 = {1{`RANDOM}};
  amplifier_1_3_data_59 = _RAND_3123[7:0];
  _RAND_3124 = {1{`RANDOM}};
  amplifier_1_3_data_60 = _RAND_3124[7:0];
  _RAND_3125 = {1{`RANDOM}};
  amplifier_1_3_data_61 = _RAND_3125[7:0];
  _RAND_3126 = {1{`RANDOM}};
  amplifier_1_3_data_62 = _RAND_3126[7:0];
  _RAND_3127 = {1{`RANDOM}};
  amplifier_1_3_data_63 = _RAND_3127[7:0];
  _RAND_3128 = {1{`RANDOM}};
  amplifier_1_3_data_64 = _RAND_3128[7:0];
  _RAND_3129 = {1{`RANDOM}};
  amplifier_1_3_data_65 = _RAND_3129[7:0];
  _RAND_3130 = {1{`RANDOM}};
  amplifier_1_3_data_66 = _RAND_3130[7:0];
  _RAND_3131 = {1{`RANDOM}};
  amplifier_1_3_data_67 = _RAND_3131[7:0];
  _RAND_3132 = {1{`RANDOM}};
  amplifier_1_3_data_68 = _RAND_3132[7:0];
  _RAND_3133 = {1{`RANDOM}};
  amplifier_1_3_data_69 = _RAND_3133[7:0];
  _RAND_3134 = {1{`RANDOM}};
  amplifier_1_3_data_70 = _RAND_3134[7:0];
  _RAND_3135 = {1{`RANDOM}};
  amplifier_1_3_data_71 = _RAND_3135[7:0];
  _RAND_3136 = {1{`RANDOM}};
  amplifier_1_3_data_72 = _RAND_3136[7:0];
  _RAND_3137 = {1{`RANDOM}};
  amplifier_1_3_data_73 = _RAND_3137[7:0];
  _RAND_3138 = {1{`RANDOM}};
  amplifier_1_3_data_74 = _RAND_3138[7:0];
  _RAND_3139 = {1{`RANDOM}};
  amplifier_1_3_data_75 = _RAND_3139[7:0];
  _RAND_3140 = {1{`RANDOM}};
  amplifier_1_3_data_76 = _RAND_3140[7:0];
  _RAND_3141 = {1{`RANDOM}};
  amplifier_1_3_data_77 = _RAND_3141[7:0];
  _RAND_3142 = {1{`RANDOM}};
  amplifier_1_3_data_78 = _RAND_3142[7:0];
  _RAND_3143 = {1{`RANDOM}};
  amplifier_1_3_data_79 = _RAND_3143[7:0];
  _RAND_3144 = {1{`RANDOM}};
  amplifier_1_3_data_80 = _RAND_3144[7:0];
  _RAND_3145 = {1{`RANDOM}};
  amplifier_1_3_data_81 = _RAND_3145[7:0];
  _RAND_3146 = {1{`RANDOM}};
  amplifier_1_3_data_82 = _RAND_3146[7:0];
  _RAND_3147 = {1{`RANDOM}};
  amplifier_1_3_data_83 = _RAND_3147[7:0];
  _RAND_3148 = {1{`RANDOM}};
  amplifier_1_3_data_84 = _RAND_3148[7:0];
  _RAND_3149 = {1{`RANDOM}};
  amplifier_1_3_data_85 = _RAND_3149[7:0];
  _RAND_3150 = {1{`RANDOM}};
  amplifier_1_3_data_86 = _RAND_3150[7:0];
  _RAND_3151 = {1{`RANDOM}};
  amplifier_1_3_data_87 = _RAND_3151[7:0];
  _RAND_3152 = {1{`RANDOM}};
  amplifier_1_3_data_88 = _RAND_3152[7:0];
  _RAND_3153 = {1{`RANDOM}};
  amplifier_1_3_data_89 = _RAND_3153[7:0];
  _RAND_3154 = {1{`RANDOM}};
  amplifier_1_3_data_90 = _RAND_3154[7:0];
  _RAND_3155 = {1{`RANDOM}};
  amplifier_1_3_data_91 = _RAND_3155[7:0];
  _RAND_3156 = {1{`RANDOM}};
  amplifier_1_3_data_92 = _RAND_3156[7:0];
  _RAND_3157 = {1{`RANDOM}};
  amplifier_1_3_data_93 = _RAND_3157[7:0];
  _RAND_3158 = {1{`RANDOM}};
  amplifier_1_3_data_94 = _RAND_3158[7:0];
  _RAND_3159 = {1{`RANDOM}};
  amplifier_1_3_data_95 = _RAND_3159[7:0];
  _RAND_3160 = {1{`RANDOM}};
  amplifier_1_3_data_96 = _RAND_3160[7:0];
  _RAND_3161 = {1{`RANDOM}};
  amplifier_1_3_data_97 = _RAND_3161[7:0];
  _RAND_3162 = {1{`RANDOM}};
  amplifier_1_3_data_98 = _RAND_3162[7:0];
  _RAND_3163 = {1{`RANDOM}};
  amplifier_1_3_data_99 = _RAND_3163[7:0];
  _RAND_3164 = {1{`RANDOM}};
  amplifier_1_3_data_100 = _RAND_3164[7:0];
  _RAND_3165 = {1{`RANDOM}};
  amplifier_1_3_data_101 = _RAND_3165[7:0];
  _RAND_3166 = {1{`RANDOM}};
  amplifier_1_3_data_102 = _RAND_3166[7:0];
  _RAND_3167 = {1{`RANDOM}};
  amplifier_1_3_data_103 = _RAND_3167[7:0];
  _RAND_3168 = {1{`RANDOM}};
  amplifier_1_3_data_104 = _RAND_3168[7:0];
  _RAND_3169 = {1{`RANDOM}};
  amplifier_1_3_data_105 = _RAND_3169[7:0];
  _RAND_3170 = {1{`RANDOM}};
  amplifier_1_3_data_106 = _RAND_3170[7:0];
  _RAND_3171 = {1{`RANDOM}};
  amplifier_1_3_data_107 = _RAND_3171[7:0];
  _RAND_3172 = {1{`RANDOM}};
  amplifier_1_3_data_108 = _RAND_3172[7:0];
  _RAND_3173 = {1{`RANDOM}};
  amplifier_1_3_data_109 = _RAND_3173[7:0];
  _RAND_3174 = {1{`RANDOM}};
  amplifier_1_3_data_110 = _RAND_3174[7:0];
  _RAND_3175 = {1{`RANDOM}};
  amplifier_1_3_data_111 = _RAND_3175[7:0];
  _RAND_3176 = {1{`RANDOM}};
  amplifier_1_3_data_112 = _RAND_3176[7:0];
  _RAND_3177 = {1{`RANDOM}};
  amplifier_1_3_data_113 = _RAND_3177[7:0];
  _RAND_3178 = {1{`RANDOM}};
  amplifier_1_3_data_114 = _RAND_3178[7:0];
  _RAND_3179 = {1{`RANDOM}};
  amplifier_1_3_data_115 = _RAND_3179[7:0];
  _RAND_3180 = {1{`RANDOM}};
  amplifier_1_3_data_116 = _RAND_3180[7:0];
  _RAND_3181 = {1{`RANDOM}};
  amplifier_1_3_data_117 = _RAND_3181[7:0];
  _RAND_3182 = {1{`RANDOM}};
  amplifier_1_3_data_118 = _RAND_3182[7:0];
  _RAND_3183 = {1{`RANDOM}};
  amplifier_1_3_data_119 = _RAND_3183[7:0];
  _RAND_3184 = {1{`RANDOM}};
  amplifier_1_3_data_120 = _RAND_3184[7:0];
  _RAND_3185 = {1{`RANDOM}};
  amplifier_1_3_data_121 = _RAND_3185[7:0];
  _RAND_3186 = {1{`RANDOM}};
  amplifier_1_3_data_122 = _RAND_3186[7:0];
  _RAND_3187 = {1{`RANDOM}};
  amplifier_1_3_data_123 = _RAND_3187[7:0];
  _RAND_3188 = {1{`RANDOM}};
  amplifier_1_3_data_124 = _RAND_3188[7:0];
  _RAND_3189 = {1{`RANDOM}};
  amplifier_1_3_data_125 = _RAND_3189[7:0];
  _RAND_3190 = {1{`RANDOM}};
  amplifier_1_3_data_126 = _RAND_3190[7:0];
  _RAND_3191 = {1{`RANDOM}};
  amplifier_1_3_data_127 = _RAND_3191[7:0];
  _RAND_3192 = {1{`RANDOM}};
  amplifier_1_3_data_128 = _RAND_3192[7:0];
  _RAND_3193 = {1{`RANDOM}};
  amplifier_1_3_data_129 = _RAND_3193[7:0];
  _RAND_3194 = {1{`RANDOM}};
  amplifier_1_3_data_130 = _RAND_3194[7:0];
  _RAND_3195 = {1{`RANDOM}};
  amplifier_1_3_data_131 = _RAND_3195[7:0];
  _RAND_3196 = {1{`RANDOM}};
  amplifier_1_3_data_132 = _RAND_3196[7:0];
  _RAND_3197 = {1{`RANDOM}};
  amplifier_1_3_data_133 = _RAND_3197[7:0];
  _RAND_3198 = {1{`RANDOM}};
  amplifier_1_3_data_134 = _RAND_3198[7:0];
  _RAND_3199 = {1{`RANDOM}};
  amplifier_1_3_data_135 = _RAND_3199[7:0];
  _RAND_3200 = {1{`RANDOM}};
  amplifier_1_3_data_136 = _RAND_3200[7:0];
  _RAND_3201 = {1{`RANDOM}};
  amplifier_1_3_data_137 = _RAND_3201[7:0];
  _RAND_3202 = {1{`RANDOM}};
  amplifier_1_3_data_138 = _RAND_3202[7:0];
  _RAND_3203 = {1{`RANDOM}};
  amplifier_1_3_data_139 = _RAND_3203[7:0];
  _RAND_3204 = {1{`RANDOM}};
  amplifier_1_3_data_140 = _RAND_3204[7:0];
  _RAND_3205 = {1{`RANDOM}};
  amplifier_1_3_data_141 = _RAND_3205[7:0];
  _RAND_3206 = {1{`RANDOM}};
  amplifier_1_3_data_142 = _RAND_3206[7:0];
  _RAND_3207 = {1{`RANDOM}};
  amplifier_1_3_data_143 = _RAND_3207[7:0];
  _RAND_3208 = {1{`RANDOM}};
  amplifier_1_3_data_144 = _RAND_3208[7:0];
  _RAND_3209 = {1{`RANDOM}};
  amplifier_1_3_data_145 = _RAND_3209[7:0];
  _RAND_3210 = {1{`RANDOM}};
  amplifier_1_3_data_146 = _RAND_3210[7:0];
  _RAND_3211 = {1{`RANDOM}};
  amplifier_1_3_data_147 = _RAND_3211[7:0];
  _RAND_3212 = {1{`RANDOM}};
  amplifier_1_3_data_148 = _RAND_3212[7:0];
  _RAND_3213 = {1{`RANDOM}};
  amplifier_1_3_data_149 = _RAND_3213[7:0];
  _RAND_3214 = {1{`RANDOM}};
  amplifier_1_3_data_150 = _RAND_3214[7:0];
  _RAND_3215 = {1{`RANDOM}};
  amplifier_1_3_data_151 = _RAND_3215[7:0];
  _RAND_3216 = {1{`RANDOM}};
  amplifier_1_3_data_152 = _RAND_3216[7:0];
  _RAND_3217 = {1{`RANDOM}};
  amplifier_1_3_data_153 = _RAND_3217[7:0];
  _RAND_3218 = {1{`RANDOM}};
  amplifier_1_3_data_154 = _RAND_3218[7:0];
  _RAND_3219 = {1{`RANDOM}};
  amplifier_1_3_data_155 = _RAND_3219[7:0];
  _RAND_3220 = {1{`RANDOM}};
  amplifier_1_3_data_156 = _RAND_3220[7:0];
  _RAND_3221 = {1{`RANDOM}};
  amplifier_1_3_data_157 = _RAND_3221[7:0];
  _RAND_3222 = {1{`RANDOM}};
  amplifier_1_3_data_158 = _RAND_3222[7:0];
  _RAND_3223 = {1{`RANDOM}};
  amplifier_1_3_data_159 = _RAND_3223[7:0];
  _RAND_3224 = {1{`RANDOM}};
  amplifier_1_3_data_160 = _RAND_3224[7:0];
  _RAND_3225 = {1{`RANDOM}};
  amplifier_1_3_data_161 = _RAND_3225[7:0];
  _RAND_3226 = {1{`RANDOM}};
  amplifier_1_3_data_162 = _RAND_3226[7:0];
  _RAND_3227 = {1{`RANDOM}};
  amplifier_1_3_data_163 = _RAND_3227[7:0];
  _RAND_3228 = {1{`RANDOM}};
  amplifier_1_3_data_164 = _RAND_3228[7:0];
  _RAND_3229 = {1{`RANDOM}};
  amplifier_1_3_data_165 = _RAND_3229[7:0];
  _RAND_3230 = {1{`RANDOM}};
  amplifier_1_3_data_166 = _RAND_3230[7:0];
  _RAND_3231 = {1{`RANDOM}};
  amplifier_1_3_data_167 = _RAND_3231[7:0];
  _RAND_3232 = {1{`RANDOM}};
  amplifier_1_3_data_168 = _RAND_3232[7:0];
  _RAND_3233 = {1{`RANDOM}};
  amplifier_1_3_data_169 = _RAND_3233[7:0];
  _RAND_3234 = {1{`RANDOM}};
  amplifier_1_3_data_170 = _RAND_3234[7:0];
  _RAND_3235 = {1{`RANDOM}};
  amplifier_1_3_data_171 = _RAND_3235[7:0];
  _RAND_3236 = {1{`RANDOM}};
  amplifier_1_3_data_172 = _RAND_3236[7:0];
  _RAND_3237 = {1{`RANDOM}};
  amplifier_1_3_data_173 = _RAND_3237[7:0];
  _RAND_3238 = {1{`RANDOM}};
  amplifier_1_3_data_174 = _RAND_3238[7:0];
  _RAND_3239 = {1{`RANDOM}};
  amplifier_1_3_data_175 = _RAND_3239[7:0];
  _RAND_3240 = {1{`RANDOM}};
  amplifier_1_3_data_176 = _RAND_3240[7:0];
  _RAND_3241 = {1{`RANDOM}};
  amplifier_1_3_data_177 = _RAND_3241[7:0];
  _RAND_3242 = {1{`RANDOM}};
  amplifier_1_3_data_178 = _RAND_3242[7:0];
  _RAND_3243 = {1{`RANDOM}};
  amplifier_1_3_data_179 = _RAND_3243[7:0];
  _RAND_3244 = {1{`RANDOM}};
  amplifier_1_3_data_180 = _RAND_3244[7:0];
  _RAND_3245 = {1{`RANDOM}};
  amplifier_1_3_data_181 = _RAND_3245[7:0];
  _RAND_3246 = {1{`RANDOM}};
  amplifier_1_3_data_182 = _RAND_3246[7:0];
  _RAND_3247 = {1{`RANDOM}};
  amplifier_1_3_data_183 = _RAND_3247[7:0];
  _RAND_3248 = {1{`RANDOM}};
  amplifier_1_3_data_184 = _RAND_3248[7:0];
  _RAND_3249 = {1{`RANDOM}};
  amplifier_1_3_data_185 = _RAND_3249[7:0];
  _RAND_3250 = {1{`RANDOM}};
  amplifier_1_3_data_186 = _RAND_3250[7:0];
  _RAND_3251 = {1{`RANDOM}};
  amplifier_1_3_data_187 = _RAND_3251[7:0];
  _RAND_3252 = {1{`RANDOM}};
  amplifier_1_3_data_188 = _RAND_3252[7:0];
  _RAND_3253 = {1{`RANDOM}};
  amplifier_1_3_data_189 = _RAND_3253[7:0];
  _RAND_3254 = {1{`RANDOM}};
  amplifier_1_3_data_190 = _RAND_3254[7:0];
  _RAND_3255 = {1{`RANDOM}};
  amplifier_1_3_data_191 = _RAND_3255[7:0];
  _RAND_3256 = {1{`RANDOM}};
  amplifier_1_3_data_192 = _RAND_3256[7:0];
  _RAND_3257 = {1{`RANDOM}};
  amplifier_1_3_data_193 = _RAND_3257[7:0];
  _RAND_3258 = {1{`RANDOM}};
  amplifier_1_3_data_194 = _RAND_3258[7:0];
  _RAND_3259 = {1{`RANDOM}};
  amplifier_1_3_data_195 = _RAND_3259[7:0];
  _RAND_3260 = {1{`RANDOM}};
  amplifier_1_3_data_196 = _RAND_3260[7:0];
  _RAND_3261 = {1{`RANDOM}};
  amplifier_1_3_data_197 = _RAND_3261[7:0];
  _RAND_3262 = {1{`RANDOM}};
  amplifier_1_3_data_198 = _RAND_3262[7:0];
  _RAND_3263 = {1{`RANDOM}};
  amplifier_1_3_data_199 = _RAND_3263[7:0];
  _RAND_3264 = {1{`RANDOM}};
  amplifier_1_3_data_200 = _RAND_3264[7:0];
  _RAND_3265 = {1{`RANDOM}};
  amplifier_1_3_data_201 = _RAND_3265[7:0];
  _RAND_3266 = {1{`RANDOM}};
  amplifier_1_3_data_202 = _RAND_3266[7:0];
  _RAND_3267 = {1{`RANDOM}};
  amplifier_1_3_data_203 = _RAND_3267[7:0];
  _RAND_3268 = {1{`RANDOM}};
  amplifier_1_3_data_204 = _RAND_3268[7:0];
  _RAND_3269 = {1{`RANDOM}};
  amplifier_1_3_data_205 = _RAND_3269[7:0];
  _RAND_3270 = {1{`RANDOM}};
  amplifier_1_3_data_206 = _RAND_3270[7:0];
  _RAND_3271 = {1{`RANDOM}};
  amplifier_1_3_data_207 = _RAND_3271[7:0];
  _RAND_3272 = {1{`RANDOM}};
  amplifier_1_3_data_208 = _RAND_3272[7:0];
  _RAND_3273 = {1{`RANDOM}};
  amplifier_1_3_data_209 = _RAND_3273[7:0];
  _RAND_3274 = {1{`RANDOM}};
  amplifier_1_3_data_210 = _RAND_3274[7:0];
  _RAND_3275 = {1{`RANDOM}};
  amplifier_1_3_data_211 = _RAND_3275[7:0];
  _RAND_3276 = {1{`RANDOM}};
  amplifier_1_3_data_212 = _RAND_3276[7:0];
  _RAND_3277 = {1{`RANDOM}};
  amplifier_1_3_data_213 = _RAND_3277[7:0];
  _RAND_3278 = {1{`RANDOM}};
  amplifier_1_3_data_214 = _RAND_3278[7:0];
  _RAND_3279 = {1{`RANDOM}};
  amplifier_1_3_data_215 = _RAND_3279[7:0];
  _RAND_3280 = {1{`RANDOM}};
  amplifier_1_3_data_216 = _RAND_3280[7:0];
  _RAND_3281 = {1{`RANDOM}};
  amplifier_1_3_data_217 = _RAND_3281[7:0];
  _RAND_3282 = {1{`RANDOM}};
  amplifier_1_3_data_218 = _RAND_3282[7:0];
  _RAND_3283 = {1{`RANDOM}};
  amplifier_1_3_data_219 = _RAND_3283[7:0];
  _RAND_3284 = {1{`RANDOM}};
  amplifier_1_3_data_220 = _RAND_3284[7:0];
  _RAND_3285 = {1{`RANDOM}};
  amplifier_1_3_data_221 = _RAND_3285[7:0];
  _RAND_3286 = {1{`RANDOM}};
  amplifier_1_3_data_222 = _RAND_3286[7:0];
  _RAND_3287 = {1{`RANDOM}};
  amplifier_1_3_data_223 = _RAND_3287[7:0];
  _RAND_3288 = {1{`RANDOM}};
  amplifier_1_3_data_224 = _RAND_3288[7:0];
  _RAND_3289 = {1{`RANDOM}};
  amplifier_1_3_data_225 = _RAND_3289[7:0];
  _RAND_3290 = {1{`RANDOM}};
  amplifier_1_3_data_226 = _RAND_3290[7:0];
  _RAND_3291 = {1{`RANDOM}};
  amplifier_1_3_data_227 = _RAND_3291[7:0];
  _RAND_3292 = {1{`RANDOM}};
  amplifier_1_3_data_228 = _RAND_3292[7:0];
  _RAND_3293 = {1{`RANDOM}};
  amplifier_1_3_data_229 = _RAND_3293[7:0];
  _RAND_3294 = {1{`RANDOM}};
  amplifier_1_3_data_230 = _RAND_3294[7:0];
  _RAND_3295 = {1{`RANDOM}};
  amplifier_1_3_data_231 = _RAND_3295[7:0];
  _RAND_3296 = {1{`RANDOM}};
  amplifier_1_3_data_232 = _RAND_3296[7:0];
  _RAND_3297 = {1{`RANDOM}};
  amplifier_1_3_data_233 = _RAND_3297[7:0];
  _RAND_3298 = {1{`RANDOM}};
  amplifier_1_3_data_234 = _RAND_3298[7:0];
  _RAND_3299 = {1{`RANDOM}};
  amplifier_1_3_data_235 = _RAND_3299[7:0];
  _RAND_3300 = {1{`RANDOM}};
  amplifier_1_3_data_236 = _RAND_3300[7:0];
  _RAND_3301 = {1{`RANDOM}};
  amplifier_1_3_data_237 = _RAND_3301[7:0];
  _RAND_3302 = {1{`RANDOM}};
  amplifier_1_3_data_238 = _RAND_3302[7:0];
  _RAND_3303 = {1{`RANDOM}};
  amplifier_1_3_data_239 = _RAND_3303[7:0];
  _RAND_3304 = {1{`RANDOM}};
  amplifier_1_3_data_240 = _RAND_3304[7:0];
  _RAND_3305 = {1{`RANDOM}};
  amplifier_1_3_data_241 = _RAND_3305[7:0];
  _RAND_3306 = {1{`RANDOM}};
  amplifier_1_3_data_242 = _RAND_3306[7:0];
  _RAND_3307 = {1{`RANDOM}};
  amplifier_1_3_data_243 = _RAND_3307[7:0];
  _RAND_3308 = {1{`RANDOM}};
  amplifier_1_3_data_244 = _RAND_3308[7:0];
  _RAND_3309 = {1{`RANDOM}};
  amplifier_1_3_data_245 = _RAND_3309[7:0];
  _RAND_3310 = {1{`RANDOM}};
  amplifier_1_3_data_246 = _RAND_3310[7:0];
  _RAND_3311 = {1{`RANDOM}};
  amplifier_1_3_data_247 = _RAND_3311[7:0];
  _RAND_3312 = {1{`RANDOM}};
  amplifier_1_3_data_248 = _RAND_3312[7:0];
  _RAND_3313 = {1{`RANDOM}};
  amplifier_1_3_data_249 = _RAND_3313[7:0];
  _RAND_3314 = {1{`RANDOM}};
  amplifier_1_3_data_250 = _RAND_3314[7:0];
  _RAND_3315 = {1{`RANDOM}};
  amplifier_1_3_data_251 = _RAND_3315[7:0];
  _RAND_3316 = {1{`RANDOM}};
  amplifier_1_3_data_252 = _RAND_3316[7:0];
  _RAND_3317 = {1{`RANDOM}};
  amplifier_1_3_data_253 = _RAND_3317[7:0];
  _RAND_3318 = {1{`RANDOM}};
  amplifier_1_3_data_254 = _RAND_3318[7:0];
  _RAND_3319 = {1{`RANDOM}};
  amplifier_1_3_data_255 = _RAND_3319[7:0];
  _RAND_3320 = {1{`RANDOM}};
  amplifier_1_3_header_0 = _RAND_3320[15:0];
  _RAND_3321 = {1{`RANDOM}};
  amplifier_1_3_header_1 = _RAND_3321[15:0];
  _RAND_3322 = {1{`RANDOM}};
  amplifier_1_3_header_2 = _RAND_3322[15:0];
  _RAND_3323 = {1{`RANDOM}};
  amplifier_1_3_header_3 = _RAND_3323[15:0];
  _RAND_3324 = {1{`RANDOM}};
  amplifier_1_3_header_4 = _RAND_3324[15:0];
  _RAND_3325 = {1{`RANDOM}};
  amplifier_1_3_header_5 = _RAND_3325[15:0];
  _RAND_3326 = {1{`RANDOM}};
  amplifier_1_3_header_6 = _RAND_3326[15:0];
  _RAND_3327 = {1{`RANDOM}};
  amplifier_1_3_header_7 = _RAND_3327[15:0];
  _RAND_3328 = {1{`RANDOM}};
  amplifier_1_3_header_8 = _RAND_3328[15:0];
  _RAND_3329 = {1{`RANDOM}};
  amplifier_1_3_header_9 = _RAND_3329[15:0];
  _RAND_3330 = {1{`RANDOM}};
  amplifier_1_3_header_10 = _RAND_3330[15:0];
  _RAND_3331 = {1{`RANDOM}};
  amplifier_1_3_header_11 = _RAND_3331[15:0];
  _RAND_3332 = {1{`RANDOM}};
  amplifier_1_3_header_12 = _RAND_3332[15:0];
  _RAND_3333 = {1{`RANDOM}};
  amplifier_1_3_header_13 = _RAND_3333[15:0];
  _RAND_3334 = {1{`RANDOM}};
  amplifier_1_3_header_14 = _RAND_3334[15:0];
  _RAND_3335 = {1{`RANDOM}};
  amplifier_1_3_header_15 = _RAND_3335[15:0];
  _RAND_3336 = {1{`RANDOM}};
  amplifier_1_3_parse_current_state = _RAND_3336[7:0];
  _RAND_3337 = {1{`RANDOM}};
  amplifier_1_3_parse_current_offset = _RAND_3337[7:0];
  _RAND_3338 = {1{`RANDOM}};
  amplifier_1_3_parse_transition_field = _RAND_3338[15:0];
  _RAND_3339 = {1{`RANDOM}};
  amplifier_1_3_next_processor_id = _RAND_3339[1:0];
  _RAND_3340 = {1{`RANDOM}};
  amplifier_1_3_next_config_id = _RAND_3340[0:0];
  _RAND_3341 = {1{`RANDOM}};
  amplifier_1_3_is_valid_processor = _RAND_3341[0:0];
  _RAND_3342 = {1{`RANDOM}};
  next_proc_id_buf_0_0 = _RAND_3342[1:0];
  _RAND_3343 = {1{`RANDOM}};
  next_proc_id_buf_0_1 = _RAND_3343[1:0];
  _RAND_3344 = {1{`RANDOM}};
  next_proc_id_buf_0_2 = _RAND_3344[1:0];
  _RAND_3345 = {1{`RANDOM}};
  next_proc_id_buf_0_3 = _RAND_3345[1:0];
  _RAND_3346 = {1{`RANDOM}};
  next_proc_id_buf_1_0 = _RAND_3346[1:0];
  _RAND_3347 = {1{`RANDOM}};
  next_proc_id_buf_1_1 = _RAND_3347[1:0];
  _RAND_3348 = {1{`RANDOM}};
  next_proc_id_buf_1_2 = _RAND_3348[1:0];
  _RAND_3349 = {1{`RANDOM}};
  next_proc_id_buf_1_3 = _RAND_3349[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
