module Executor(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input         io_hit,
  input  [63:0] io_match_value,
  input         io_action_mod_en,
  input  [7:0]  io_action_mod_addr,
  input  [63:0] io_action_mod_data_0,
  input  [63:0] io_action_mod_data_1
);
  wire  pipe1_clock; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_0; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_1; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_2; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_3; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_4; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_5; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_6; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_7; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_8; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_9; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_10; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_11; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_12; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_13; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_14; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_15; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_16; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_17; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_18; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_19; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_20; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_21; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_22; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_23; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_24; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_25; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_26; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_27; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_28; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_29; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_30; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_31; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_32; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_33; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_34; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_35; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_36; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_37; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_38; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_39; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_40; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_41; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_42; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_43; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_44; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_45; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_46; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_47; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_48; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_49; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_50; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_51; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_52; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_53; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_54; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_55; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_56; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_57; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_58; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_59; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_60; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_61; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_62; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_63; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_64; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_65; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_66; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_67; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_68; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_69; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_70; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_71; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_72; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_73; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_74; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_75; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_76; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_77; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_78; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_79; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_80; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_81; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_82; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_83; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_84; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_85; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_86; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_87; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_88; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_89; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_90; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_91; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_92; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_93; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_94; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_95; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_0; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_1; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_2; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_3; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_4; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_5; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_6; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_7; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_8; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_9; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_10; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_11; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_12; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_13; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_14; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_15; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_state; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_offset; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_in_parse_transition_field; // @[executor.scala 317:23]
  wire [1:0] pipe1_io_pipe_phv_in_next_processor_id; // @[executor.scala 317:23]
  wire  pipe1_io_pipe_phv_in_next_config_id; // @[executor.scala 317:23]
  wire  pipe1_io_pipe_phv_in_is_valid_processor; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_0; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_1; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_2; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_3; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_4; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_5; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_6; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_7; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_8; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_9; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_10; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_11; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_12; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_13; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_14; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_15; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_16; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_17; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_18; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_19; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_20; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_21; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_22; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_23; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_24; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_25; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_26; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_27; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_28; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_29; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_30; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_31; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_32; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_33; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_34; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_35; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_36; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_37; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_38; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_39; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_40; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_41; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_42; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_43; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_44; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_45; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_46; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_47; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_48; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_49; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_50; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_51; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_52; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_53; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_54; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_55; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_56; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_57; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_58; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_59; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_60; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_61; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_62; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_63; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_64; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_65; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_66; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_67; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_68; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_69; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_70; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_71; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_72; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_73; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_74; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_75; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_76; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_77; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_78; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_79; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_80; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_81; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_82; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_83; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_84; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_85; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_86; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_87; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_88; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_89; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_90; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_91; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_92; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_93; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_94; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_95; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_0; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_1; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_2; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_3; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_4; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_5; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_6; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_7; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_8; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_9; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_10; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_11; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_12; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_13; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_14; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_15; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_state; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_offset; // @[executor.scala 317:23]
  wire [15:0] pipe1_io_pipe_phv_out_parse_transition_field; // @[executor.scala 317:23]
  wire [1:0] pipe1_io_pipe_phv_out_next_processor_id; // @[executor.scala 317:23]
  wire  pipe1_io_pipe_phv_out_next_config_id; // @[executor.scala 317:23]
  wire  pipe1_io_pipe_phv_out_is_valid_processor; // @[executor.scala 317:23]
  wire  pipe1_io_hit; // @[executor.scala 317:23]
  wire [63:0] pipe1_io_match_value; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_args_out_0; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_args_out_1; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_args_out_2; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_args_out_3; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_args_out_4; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_args_out_5; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_args_out_6; // @[executor.scala 317:23]
  wire [31:0] pipe1_io_vliw_out_0; // @[executor.scala 317:23]
  wire [31:0] pipe1_io_vliw_out_1; // @[executor.scala 317:23]
  wire [31:0] pipe1_io_vliw_out_2; // @[executor.scala 317:23]
  wire [31:0] pipe1_io_vliw_out_3; // @[executor.scala 317:23]
  wire  pipe1_io_action_mod_en; // @[executor.scala 317:23]
  wire [7:0] pipe1_io_action_mod_addr; // @[executor.scala 317:23]
  wire [63:0] pipe1_io_action_mod_data_0; // @[executor.scala 317:23]
  wire [63:0] pipe1_io_action_mod_data_1; // @[executor.scala 317:23]
  wire  pipe2_clock; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_0; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_1; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_2; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_3; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_4; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_5; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_6; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_7; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_8; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_9; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_10; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_11; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_12; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_13; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_14; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_15; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_16; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_17; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_18; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_19; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_20; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_21; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_22; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_23; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_24; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_25; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_26; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_27; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_28; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_29; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_30; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_31; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_32; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_33; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_34; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_35; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_36; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_37; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_38; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_39; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_40; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_41; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_42; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_43; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_44; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_45; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_46; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_47; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_48; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_49; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_50; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_51; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_52; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_53; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_54; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_55; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_56; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_57; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_58; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_59; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_60; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_61; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_62; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_63; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_64; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_65; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_66; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_67; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_68; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_69; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_70; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_71; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_72; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_73; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_74; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_75; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_76; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_77; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_78; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_79; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_80; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_81; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_82; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_83; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_84; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_85; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_86; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_87; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_88; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_89; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_90; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_91; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_92; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_93; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_94; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_95; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_0; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_1; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_2; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_3; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_4; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_5; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_6; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_7; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_8; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_9; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_10; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_11; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_12; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_13; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_14; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_15; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_state; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_offset; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_in_parse_transition_field; // @[executor.scala 318:23]
  wire [1:0] pipe2_io_pipe_phv_in_next_processor_id; // @[executor.scala 318:23]
  wire  pipe2_io_pipe_phv_in_next_config_id; // @[executor.scala 318:23]
  wire  pipe2_io_pipe_phv_in_is_valid_processor; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_0; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_1; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_2; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_3; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_4; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_5; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_6; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_7; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_8; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_9; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_10; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_11; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_12; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_13; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_14; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_15; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_16; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_17; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_18; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_19; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_20; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_21; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_22; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_23; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_24; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_25; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_26; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_27; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_28; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_29; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_30; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_31; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_32; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_33; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_34; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_35; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_36; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_37; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_38; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_39; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_40; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_41; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_42; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_43; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_44; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_45; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_46; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_47; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_48; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_49; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_50; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_51; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_52; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_53; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_54; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_55; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_56; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_57; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_58; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_59; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_60; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_61; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_62; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_63; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_64; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_65; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_66; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_67; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_68; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_69; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_70; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_71; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_72; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_73; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_74; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_75; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_76; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_77; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_78; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_79; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_80; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_81; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_82; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_83; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_84; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_85; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_86; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_87; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_88; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_89; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_90; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_91; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_92; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_93; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_94; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_95; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_0; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_1; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_2; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_3; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_4; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_5; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_6; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_7; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_8; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_9; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_10; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_11; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_12; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_13; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_14; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_15; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_state; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_offset; // @[executor.scala 318:23]
  wire [15:0] pipe2_io_pipe_phv_out_parse_transition_field; // @[executor.scala 318:23]
  wire [1:0] pipe2_io_pipe_phv_out_next_processor_id; // @[executor.scala 318:23]
  wire  pipe2_io_pipe_phv_out_next_config_id; // @[executor.scala 318:23]
  wire  pipe2_io_pipe_phv_out_is_valid_processor; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_args_in_0; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_args_in_1; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_args_in_2; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_args_in_3; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_args_in_4; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_args_in_5; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_args_in_6; // @[executor.scala 318:23]
  wire [31:0] pipe2_io_vliw_in_0; // @[executor.scala 318:23]
  wire [31:0] pipe2_io_vliw_in_1; // @[executor.scala 318:23]
  wire [31:0] pipe2_io_vliw_in_2; // @[executor.scala 318:23]
  wire [31:0] pipe2_io_vliw_in_3; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_args_out_0; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_args_out_1; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_args_out_2; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_args_out_3; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_args_out_4; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_args_out_5; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_args_out_6; // @[executor.scala 318:23]
  wire [31:0] pipe2_io_vliw_out_0; // @[executor.scala 318:23]
  wire [31:0] pipe2_io_vliw_out_1; // @[executor.scala 318:23]
  wire [31:0] pipe2_io_vliw_out_2; // @[executor.scala 318:23]
  wire [31:0] pipe2_io_vliw_out_3; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_offset_out_0; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_offset_out_1; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_offset_out_2; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_offset_out_3; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_length_out_0; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_length_out_1; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_length_out_2; // @[executor.scala 318:23]
  wire [7:0] pipe2_io_length_out_3; // @[executor.scala 318:23]
  wire  pipe3_clock; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_0; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_1; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_2; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_3; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_4; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_5; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_6; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_7; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_8; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_9; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_10; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_11; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_12; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_13; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_14; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_15; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_16; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_17; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_18; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_19; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_20; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_21; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_22; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_23; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_24; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_25; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_26; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_27; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_28; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_29; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_30; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_31; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_32; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_33; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_34; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_35; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_36; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_37; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_38; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_39; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_40; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_41; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_42; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_43; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_44; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_45; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_46; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_47; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_48; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_49; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_50; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_51; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_52; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_53; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_54; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_55; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_56; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_57; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_58; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_59; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_60; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_61; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_62; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_63; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_64; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_65; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_66; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_67; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_68; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_69; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_70; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_71; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_72; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_73; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_74; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_75; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_76; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_77; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_78; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_79; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_80; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_81; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_82; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_83; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_84; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_85; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_86; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_87; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_88; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_89; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_90; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_91; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_92; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_93; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_94; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_95; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_0; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_1; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_2; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_3; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_4; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_5; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_6; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_7; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_8; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_9; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_10; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_11; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_12; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_13; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_14; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_15; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_parse_current_state; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_in_parse_current_offset; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_in_parse_transition_field; // @[executor.scala 319:23]
  wire [1:0] pipe3_io_pipe_phv_in_next_processor_id; // @[executor.scala 319:23]
  wire  pipe3_io_pipe_phv_in_next_config_id; // @[executor.scala 319:23]
  wire  pipe3_io_pipe_phv_in_is_valid_processor; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_0; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_1; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_2; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_3; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_4; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_5; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_6; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_7; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_8; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_9; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_10; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_11; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_12; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_13; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_14; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_15; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_16; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_17; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_18; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_19; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_20; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_21; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_22; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_23; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_24; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_25; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_26; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_27; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_28; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_29; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_30; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_31; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_32; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_33; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_34; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_35; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_36; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_37; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_38; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_39; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_40; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_41; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_42; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_43; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_44; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_45; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_46; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_47; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_48; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_49; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_50; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_51; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_52; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_53; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_54; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_55; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_56; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_57; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_58; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_59; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_60; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_61; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_62; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_63; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_64; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_65; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_66; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_67; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_68; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_69; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_70; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_71; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_72; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_73; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_74; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_75; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_76; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_77; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_78; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_79; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_80; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_81; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_82; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_83; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_84; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_85; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_86; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_87; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_88; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_89; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_90; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_91; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_92; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_93; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_94; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_95; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_0; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_1; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_2; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_3; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_4; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_5; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_6; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_7; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_8; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_9; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_10; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_11; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_12; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_13; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_14; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_15; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_parse_current_state; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_pipe_phv_out_parse_current_offset; // @[executor.scala 319:23]
  wire [15:0] pipe3_io_pipe_phv_out_parse_transition_field; // @[executor.scala 319:23]
  wire [1:0] pipe3_io_pipe_phv_out_next_processor_id; // @[executor.scala 319:23]
  wire  pipe3_io_pipe_phv_out_next_config_id; // @[executor.scala 319:23]
  wire  pipe3_io_pipe_phv_out_is_valid_processor; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_args_in_0; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_args_in_1; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_args_in_2; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_args_in_3; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_args_in_4; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_args_in_5; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_args_in_6; // @[executor.scala 319:23]
  wire [31:0] pipe3_io_vliw_in_0; // @[executor.scala 319:23]
  wire [31:0] pipe3_io_vliw_in_1; // @[executor.scala 319:23]
  wire [31:0] pipe3_io_vliw_in_2; // @[executor.scala 319:23]
  wire [31:0] pipe3_io_vliw_in_3; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_offset_in_0; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_offset_in_1; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_offset_in_2; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_offset_in_3; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_length_in_0; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_length_in_1; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_length_in_2; // @[executor.scala 319:23]
  wire [7:0] pipe3_io_length_in_3; // @[executor.scala 319:23]
  wire [31:0] pipe3_io_vliw_out_0; // @[executor.scala 319:23]
  wire [31:0] pipe3_io_vliw_out_1; // @[executor.scala 319:23]
  wire [31:0] pipe3_io_vliw_out_2; // @[executor.scala 319:23]
  wire [31:0] pipe3_io_vliw_out_3; // @[executor.scala 319:23]
  wire [63:0] pipe3_io_field_out_0; // @[executor.scala 319:23]
  wire [63:0] pipe3_io_field_out_1; // @[executor.scala 319:23]
  wire [63:0] pipe3_io_field_out_2; // @[executor.scala 319:23]
  wire [63:0] pipe3_io_field_out_3; // @[executor.scala 319:23]
  wire  pipe4_clock; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_0; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_1; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_2; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_3; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_4; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_5; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_6; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_7; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_8; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_9; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_10; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_11; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_12; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_13; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_14; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_15; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_16; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_17; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_18; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_19; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_20; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_21; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_22; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_23; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_24; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_25; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_26; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_27; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_28; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_29; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_30; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_31; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_32; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_33; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_34; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_35; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_36; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_37; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_38; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_39; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_40; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_41; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_42; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_43; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_44; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_45; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_46; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_47; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_48; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_49; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_50; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_51; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_52; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_53; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_54; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_55; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_56; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_57; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_58; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_59; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_60; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_61; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_62; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_63; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_64; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_65; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_66; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_67; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_68; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_69; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_70; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_71; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_72; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_73; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_74; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_75; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_76; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_77; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_78; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_79; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_80; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_81; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_82; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_83; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_84; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_85; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_86; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_87; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_88; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_89; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_90; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_91; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_92; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_93; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_94; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_95; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_0; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_1; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_2; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_3; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_4; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_5; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_6; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_7; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_8; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_9; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_10; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_11; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_12; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_13; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_14; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_15; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_parse_current_state; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_in_parse_current_offset; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_in_parse_transition_field; // @[executor.scala 320:23]
  wire [1:0] pipe4_io_pipe_phv_in_next_processor_id; // @[executor.scala 320:23]
  wire  pipe4_io_pipe_phv_in_next_config_id; // @[executor.scala 320:23]
  wire  pipe4_io_pipe_phv_in_is_valid_processor; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_0; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_1; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_2; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_3; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_4; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_5; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_6; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_7; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_8; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_9; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_10; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_11; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_12; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_13; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_14; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_15; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_16; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_17; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_18; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_19; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_20; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_21; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_22; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_23; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_24; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_25; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_26; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_27; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_28; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_29; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_30; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_31; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_32; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_33; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_34; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_35; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_36; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_37; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_38; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_39; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_40; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_41; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_42; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_43; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_44; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_45; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_46; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_47; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_48; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_49; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_50; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_51; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_52; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_53; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_54; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_55; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_56; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_57; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_58; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_59; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_60; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_61; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_62; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_63; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_64; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_65; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_66; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_67; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_68; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_69; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_70; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_71; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_72; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_73; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_74; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_75; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_76; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_77; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_78; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_79; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_80; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_81; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_82; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_83; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_84; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_85; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_86; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_87; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_88; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_89; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_90; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_91; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_92; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_93; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_94; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_95; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_0; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_1; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_2; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_3; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_4; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_5; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_6; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_7; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_8; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_9; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_10; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_11; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_12; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_13; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_14; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_15; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_parse_current_state; // @[executor.scala 320:23]
  wire [7:0] pipe4_io_pipe_phv_out_parse_current_offset; // @[executor.scala 320:23]
  wire [15:0] pipe4_io_pipe_phv_out_parse_transition_field; // @[executor.scala 320:23]
  wire [1:0] pipe4_io_pipe_phv_out_next_processor_id; // @[executor.scala 320:23]
  wire  pipe4_io_pipe_phv_out_next_config_id; // @[executor.scala 320:23]
  wire  pipe4_io_pipe_phv_out_is_valid_processor; // @[executor.scala 320:23]
  wire [31:0] pipe4_io_vliw_in_0; // @[executor.scala 320:23]
  wire [31:0] pipe4_io_vliw_in_1; // @[executor.scala 320:23]
  wire [31:0] pipe4_io_vliw_in_2; // @[executor.scala 320:23]
  wire [31:0] pipe4_io_vliw_in_3; // @[executor.scala 320:23]
  wire [63:0] pipe4_io_field_in_0; // @[executor.scala 320:23]
  wire [63:0] pipe4_io_field_in_1; // @[executor.scala 320:23]
  wire [63:0] pipe4_io_field_in_2; // @[executor.scala 320:23]
  wire [63:0] pipe4_io_field_in_3; // @[executor.scala 320:23]
  wire [31:0] pipe4_io_vliw_out_0; // @[executor.scala 320:23]
  wire [31:0] pipe4_io_vliw_out_1; // @[executor.scala 320:23]
  wire [31:0] pipe4_io_vliw_out_2; // @[executor.scala 320:23]
  wire [31:0] pipe4_io_vliw_out_3; // @[executor.scala 320:23]
  wire [63:0] pipe4_io_field_out_0; // @[executor.scala 320:23]
  wire [63:0] pipe4_io_field_out_1; // @[executor.scala 320:23]
  wire [63:0] pipe4_io_field_out_2; // @[executor.scala 320:23]
  wire [63:0] pipe4_io_field_out_3; // @[executor.scala 320:23]
  wire  pipe5_clock; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_0; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_1; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_2; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_3; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_4; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_5; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_6; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_7; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_8; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_9; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_10; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_11; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_12; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_13; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_14; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_15; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_16; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_17; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_18; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_19; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_20; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_21; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_22; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_23; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_24; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_25; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_26; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_27; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_28; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_29; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_30; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_31; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_32; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_33; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_34; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_35; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_36; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_37; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_38; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_39; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_40; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_41; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_42; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_43; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_44; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_45; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_46; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_47; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_48; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_49; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_50; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_51; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_52; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_53; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_54; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_55; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_56; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_57; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_58; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_59; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_60; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_61; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_62; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_63; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_64; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_65; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_66; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_67; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_68; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_69; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_70; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_71; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_72; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_73; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_74; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_75; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_76; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_77; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_78; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_79; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_80; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_81; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_82; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_83; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_84; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_85; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_86; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_87; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_88; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_89; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_90; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_91; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_92; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_93; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_94; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_95; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_0; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_1; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_2; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_3; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_4; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_5; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_6; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_7; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_8; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_9; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_10; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_11; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_12; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_13; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_14; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_15; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_parse_current_state; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_in_parse_current_offset; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_in_parse_transition_field; // @[executor.scala 321:23]
  wire [1:0] pipe5_io_pipe_phv_in_next_processor_id; // @[executor.scala 321:23]
  wire  pipe5_io_pipe_phv_in_next_config_id; // @[executor.scala 321:23]
  wire  pipe5_io_pipe_phv_in_is_valid_processor; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_0; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_1; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_2; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_3; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_4; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_5; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_6; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_7; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_8; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_9; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_10; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_11; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_12; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_13; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_14; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_15; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_16; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_17; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_18; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_19; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_20; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_21; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_22; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_23; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_24; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_25; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_26; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_27; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_28; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_29; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_30; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_31; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_32; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_33; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_34; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_35; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_36; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_37; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_38; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_39; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_40; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_41; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_42; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_43; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_44; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_45; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_46; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_47; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_48; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_49; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_50; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_51; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_52; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_53; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_54; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_55; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_56; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_57; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_58; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_59; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_60; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_61; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_62; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_63; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_64; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_65; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_66; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_67; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_68; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_69; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_70; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_71; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_72; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_73; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_74; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_75; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_76; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_77; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_78; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_79; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_80; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_81; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_82; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_83; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_84; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_85; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_86; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_87; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_88; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_89; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_90; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_91; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_92; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_93; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_94; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_95; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_0; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_1; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_2; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_3; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_4; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_5; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_6; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_7; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_8; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_9; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_10; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_11; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_12; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_13; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_14; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_15; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_parse_current_state; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_pipe_phv_out_parse_current_offset; // @[executor.scala 321:23]
  wire [15:0] pipe5_io_pipe_phv_out_parse_transition_field; // @[executor.scala 321:23]
  wire [1:0] pipe5_io_pipe_phv_out_next_processor_id; // @[executor.scala 321:23]
  wire  pipe5_io_pipe_phv_out_next_config_id; // @[executor.scala 321:23]
  wire  pipe5_io_pipe_phv_out_is_valid_processor; // @[executor.scala 321:23]
  wire [31:0] pipe5_io_vliw_in_0; // @[executor.scala 321:23]
  wire [31:0] pipe5_io_vliw_in_1; // @[executor.scala 321:23]
  wire [31:0] pipe5_io_vliw_in_2; // @[executor.scala 321:23]
  wire [31:0] pipe5_io_vliw_in_3; // @[executor.scala 321:23]
  wire [63:0] pipe5_io_field_in_0; // @[executor.scala 321:23]
  wire [63:0] pipe5_io_field_in_1; // @[executor.scala 321:23]
  wire [63:0] pipe5_io_field_in_2; // @[executor.scala 321:23]
  wire [63:0] pipe5_io_field_in_3; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_offset_out_0; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_offset_out_1; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_offset_out_2; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_offset_out_3; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_length_out_0; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_length_out_1; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_length_out_2; // @[executor.scala 321:23]
  wire [7:0] pipe5_io_length_out_3; // @[executor.scala 321:23]
  wire [63:0] pipe5_io_field_out_0; // @[executor.scala 321:23]
  wire [63:0] pipe5_io_field_out_1; // @[executor.scala 321:23]
  wire [63:0] pipe5_io_field_out_2; // @[executor.scala 321:23]
  wire [63:0] pipe5_io_field_out_3; // @[executor.scala 321:23]
  wire  pipe6_clock; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_0; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_1; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_2; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_3; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_4; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_5; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_6; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_7; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_8; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_9; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_10; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_11; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_12; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_13; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_14; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_15; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_16; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_17; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_18; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_19; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_20; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_21; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_22; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_23; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_24; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_25; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_26; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_27; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_28; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_29; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_30; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_31; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_32; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_33; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_34; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_35; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_36; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_37; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_38; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_39; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_40; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_41; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_42; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_43; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_44; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_45; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_46; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_47; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_48; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_49; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_50; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_51; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_52; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_53; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_54; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_55; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_56; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_57; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_58; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_59; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_60; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_61; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_62; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_63; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_64; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_65; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_66; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_67; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_68; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_69; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_70; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_71; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_72; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_73; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_74; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_75; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_76; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_77; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_78; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_79; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_80; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_81; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_82; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_83; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_84; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_85; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_86; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_87; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_88; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_89; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_90; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_91; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_92; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_93; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_94; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_95; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_0; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_1; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_2; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_3; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_4; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_5; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_6; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_7; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_8; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_9; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_10; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_11; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_12; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_13; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_14; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_15; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_parse_current_state; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_in_parse_current_offset; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_in_parse_transition_field; // @[executor.scala 322:23]
  wire [1:0] pipe6_io_pipe_phv_in_next_processor_id; // @[executor.scala 322:23]
  wire  pipe6_io_pipe_phv_in_next_config_id; // @[executor.scala 322:23]
  wire  pipe6_io_pipe_phv_in_is_valid_processor; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_0; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_1; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_2; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_3; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_4; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_5; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_6; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_7; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_8; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_9; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_10; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_11; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_12; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_13; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_14; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_15; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_16; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_17; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_18; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_19; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_20; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_21; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_22; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_23; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_24; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_25; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_26; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_27; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_28; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_29; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_30; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_31; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_32; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_33; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_34; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_35; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_36; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_37; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_38; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_39; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_40; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_41; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_42; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_43; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_44; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_45; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_46; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_47; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_48; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_49; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_50; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_51; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_52; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_53; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_54; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_55; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_56; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_57; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_58; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_59; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_60; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_61; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_62; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_63; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_64; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_65; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_66; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_67; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_68; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_69; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_70; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_71; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_72; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_73; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_74; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_75; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_76; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_77; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_78; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_79; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_80; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_81; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_82; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_83; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_84; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_85; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_86; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_87; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_88; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_89; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_90; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_91; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_92; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_93; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_94; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_95; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_0; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_1; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_2; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_3; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_4; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_5; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_6; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_7; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_8; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_9; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_10; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_11; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_12; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_13; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_14; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_15; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_parse_current_state; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_pipe_phv_out_parse_current_offset; // @[executor.scala 322:23]
  wire [15:0] pipe6_io_pipe_phv_out_parse_transition_field; // @[executor.scala 322:23]
  wire [1:0] pipe6_io_pipe_phv_out_next_processor_id; // @[executor.scala 322:23]
  wire  pipe6_io_pipe_phv_out_next_config_id; // @[executor.scala 322:23]
  wire  pipe6_io_pipe_phv_out_is_valid_processor; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_offset_in_0; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_offset_in_1; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_offset_in_2; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_offset_in_3; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_length_in_0; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_length_in_1; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_length_in_2; // @[executor.scala 322:23]
  wire [7:0] pipe6_io_length_in_3; // @[executor.scala 322:23]
  wire [63:0] pipe6_io_field_in_0; // @[executor.scala 322:23]
  wire [63:0] pipe6_io_field_in_1; // @[executor.scala 322:23]
  wire [63:0] pipe6_io_field_in_2; // @[executor.scala 322:23]
  wire [63:0] pipe6_io_field_in_3; // @[executor.scala 322:23]
  ActionReader pipe1 ( // @[executor.scala 317:23]
    .clock(pipe1_clock),
    .io_pipe_phv_in_data_0(pipe1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe1_io_pipe_phv_out_is_valid_processor),
    .io_hit(pipe1_io_hit),
    .io_match_value(pipe1_io_match_value),
    .io_args_out_0(pipe1_io_args_out_0),
    .io_args_out_1(pipe1_io_args_out_1),
    .io_args_out_2(pipe1_io_args_out_2),
    .io_args_out_3(pipe1_io_args_out_3),
    .io_args_out_4(pipe1_io_args_out_4),
    .io_args_out_5(pipe1_io_args_out_5),
    .io_args_out_6(pipe1_io_args_out_6),
    .io_vliw_out_0(pipe1_io_vliw_out_0),
    .io_vliw_out_1(pipe1_io_vliw_out_1),
    .io_vliw_out_2(pipe1_io_vliw_out_2),
    .io_vliw_out_3(pipe1_io_vliw_out_3),
    .io_action_mod_en(pipe1_io_action_mod_en),
    .io_action_mod_addr(pipe1_io_action_mod_addr),
    .io_action_mod_data_0(pipe1_io_action_mod_data_0),
    .io_action_mod_data_1(pipe1_io_action_mod_data_1)
  );
  PrimitiveGetOffset pipe2 ( // @[executor.scala 318:23]
    .clock(pipe2_clock),
    .io_pipe_phv_in_data_0(pipe2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe2_io_pipe_phv_out_is_valid_processor),
    .io_args_in_0(pipe2_io_args_in_0),
    .io_args_in_1(pipe2_io_args_in_1),
    .io_args_in_2(pipe2_io_args_in_2),
    .io_args_in_3(pipe2_io_args_in_3),
    .io_args_in_4(pipe2_io_args_in_4),
    .io_args_in_5(pipe2_io_args_in_5),
    .io_args_in_6(pipe2_io_args_in_6),
    .io_vliw_in_0(pipe2_io_vliw_in_0),
    .io_vliw_in_1(pipe2_io_vliw_in_1),
    .io_vliw_in_2(pipe2_io_vliw_in_2),
    .io_vliw_in_3(pipe2_io_vliw_in_3),
    .io_args_out_0(pipe2_io_args_out_0),
    .io_args_out_1(pipe2_io_args_out_1),
    .io_args_out_2(pipe2_io_args_out_2),
    .io_args_out_3(pipe2_io_args_out_3),
    .io_args_out_4(pipe2_io_args_out_4),
    .io_args_out_5(pipe2_io_args_out_5),
    .io_args_out_6(pipe2_io_args_out_6),
    .io_vliw_out_0(pipe2_io_vliw_out_0),
    .io_vliw_out_1(pipe2_io_vliw_out_1),
    .io_vliw_out_2(pipe2_io_vliw_out_2),
    .io_vliw_out_3(pipe2_io_vliw_out_3),
    .io_offset_out_0(pipe2_io_offset_out_0),
    .io_offset_out_1(pipe2_io_offset_out_1),
    .io_offset_out_2(pipe2_io_offset_out_2),
    .io_offset_out_3(pipe2_io_offset_out_3),
    .io_length_out_0(pipe2_io_length_out_0),
    .io_length_out_1(pipe2_io_length_out_1),
    .io_length_out_2(pipe2_io_length_out_2),
    .io_length_out_3(pipe2_io_length_out_3)
  );
  PrimitiveGetSource pipe3 ( // @[executor.scala 319:23]
    .clock(pipe3_clock),
    .io_pipe_phv_in_data_0(pipe3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe3_io_pipe_phv_out_is_valid_processor),
    .io_args_in_0(pipe3_io_args_in_0),
    .io_args_in_1(pipe3_io_args_in_1),
    .io_args_in_2(pipe3_io_args_in_2),
    .io_args_in_3(pipe3_io_args_in_3),
    .io_args_in_4(pipe3_io_args_in_4),
    .io_args_in_5(pipe3_io_args_in_5),
    .io_args_in_6(pipe3_io_args_in_6),
    .io_vliw_in_0(pipe3_io_vliw_in_0),
    .io_vliw_in_1(pipe3_io_vliw_in_1),
    .io_vliw_in_2(pipe3_io_vliw_in_2),
    .io_vliw_in_3(pipe3_io_vliw_in_3),
    .io_offset_in_0(pipe3_io_offset_in_0),
    .io_offset_in_1(pipe3_io_offset_in_1),
    .io_offset_in_2(pipe3_io_offset_in_2),
    .io_offset_in_3(pipe3_io_offset_in_3),
    .io_length_in_0(pipe3_io_length_in_0),
    .io_length_in_1(pipe3_io_length_in_1),
    .io_length_in_2(pipe3_io_length_in_2),
    .io_length_in_3(pipe3_io_length_in_3),
    .io_vliw_out_0(pipe3_io_vliw_out_0),
    .io_vliw_out_1(pipe3_io_vliw_out_1),
    .io_vliw_out_2(pipe3_io_vliw_out_2),
    .io_vliw_out_3(pipe3_io_vliw_out_3),
    .io_field_out_0(pipe3_io_field_out_0),
    .io_field_out_1(pipe3_io_field_out_1),
    .io_field_out_2(pipe3_io_field_out_2),
    .io_field_out_3(pipe3_io_field_out_3)
  );
  PrimitiveALU pipe4 ( // @[executor.scala 320:23]
    .clock(pipe4_clock),
    .io_pipe_phv_in_data_0(pipe4_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe4_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe4_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe4_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe4_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe4_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe4_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe4_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe4_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe4_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe4_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe4_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe4_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe4_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe4_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe4_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe4_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe4_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe4_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe4_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe4_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe4_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe4_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe4_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe4_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe4_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe4_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe4_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe4_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe4_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe4_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe4_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe4_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe4_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe4_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe4_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe4_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe4_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe4_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe4_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe4_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe4_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe4_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe4_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe4_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe4_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe4_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe4_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe4_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe4_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe4_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe4_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe4_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe4_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe4_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe4_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe4_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe4_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe4_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe4_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe4_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe4_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe4_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe4_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe4_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe4_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe4_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe4_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe4_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe4_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe4_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe4_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe4_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe4_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe4_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe4_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe4_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe4_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe4_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe4_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe4_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe4_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe4_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe4_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe4_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe4_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe4_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe4_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe4_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe4_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe4_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe4_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe4_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe4_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe4_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe4_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe4_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe4_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe4_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe4_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe4_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe4_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe4_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe4_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe4_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe4_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe4_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe4_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe4_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe4_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe4_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe4_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe4_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe4_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe4_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe4_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe4_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe4_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe4_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe4_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe4_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe4_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe4_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe4_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe4_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe4_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe4_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe4_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe4_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe4_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe4_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe4_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe4_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe4_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe4_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe4_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe4_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe4_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe4_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe4_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe4_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe4_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe4_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe4_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe4_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe4_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe4_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe4_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe4_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe4_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe4_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe4_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe4_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe4_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe4_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe4_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe4_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe4_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe4_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe4_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe4_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe4_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe4_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe4_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe4_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe4_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe4_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe4_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe4_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe4_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe4_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe4_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe4_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe4_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe4_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe4_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe4_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe4_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe4_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe4_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe4_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe4_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe4_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe4_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe4_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe4_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe4_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe4_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe4_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe4_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe4_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe4_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe4_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe4_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe4_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe4_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe4_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe4_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe4_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe4_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe4_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe4_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe4_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe4_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe4_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe4_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe4_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe4_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe4_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe4_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe4_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe4_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe4_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe4_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe4_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe4_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe4_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe4_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe4_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe4_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe4_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe4_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe4_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe4_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe4_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe4_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe4_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe4_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe4_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe4_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe4_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe4_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe4_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe4_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe4_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe4_io_pipe_phv_out_is_valid_processor),
    .io_vliw_in_0(pipe4_io_vliw_in_0),
    .io_vliw_in_1(pipe4_io_vliw_in_1),
    .io_vliw_in_2(pipe4_io_vliw_in_2),
    .io_vliw_in_3(pipe4_io_vliw_in_3),
    .io_field_in_0(pipe4_io_field_in_0),
    .io_field_in_1(pipe4_io_field_in_1),
    .io_field_in_2(pipe4_io_field_in_2),
    .io_field_in_3(pipe4_io_field_in_3),
    .io_vliw_out_0(pipe4_io_vliw_out_0),
    .io_vliw_out_1(pipe4_io_vliw_out_1),
    .io_vliw_out_2(pipe4_io_vliw_out_2),
    .io_vliw_out_3(pipe4_io_vliw_out_3),
    .io_field_out_0(pipe4_io_field_out_0),
    .io_field_out_1(pipe4_io_field_out_1),
    .io_field_out_2(pipe4_io_field_out_2),
    .io_field_out_3(pipe4_io_field_out_3)
  );
  PrimitiveGetWriteBackOffset pipe5 ( // @[executor.scala 321:23]
    .clock(pipe5_clock),
    .io_pipe_phv_in_data_0(pipe5_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe5_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe5_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe5_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe5_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe5_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe5_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe5_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe5_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe5_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe5_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe5_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe5_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe5_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe5_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe5_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe5_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe5_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe5_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe5_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe5_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe5_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe5_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe5_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe5_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe5_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe5_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe5_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe5_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe5_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe5_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe5_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe5_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe5_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe5_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe5_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe5_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe5_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe5_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe5_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe5_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe5_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe5_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe5_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe5_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe5_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe5_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe5_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe5_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe5_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe5_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe5_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe5_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe5_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe5_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe5_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe5_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe5_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe5_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe5_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe5_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe5_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe5_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe5_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe5_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe5_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe5_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe5_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe5_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe5_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe5_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe5_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe5_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe5_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe5_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe5_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe5_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe5_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe5_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe5_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe5_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe5_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe5_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe5_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe5_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe5_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe5_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe5_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe5_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe5_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe5_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe5_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe5_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe5_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe5_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe5_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe5_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe5_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe5_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe5_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe5_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe5_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe5_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe5_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe5_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe5_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe5_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe5_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe5_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe5_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe5_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe5_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe5_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe5_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe5_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe5_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe5_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe5_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe5_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe5_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe5_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe5_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe5_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe5_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe5_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe5_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe5_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe5_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe5_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe5_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe5_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe5_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe5_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe5_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe5_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe5_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe5_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe5_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe5_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe5_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe5_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe5_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe5_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe5_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe5_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe5_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe5_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe5_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe5_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe5_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe5_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe5_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe5_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe5_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe5_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe5_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe5_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe5_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe5_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe5_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe5_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe5_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe5_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe5_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe5_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe5_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe5_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe5_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe5_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe5_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe5_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe5_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe5_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe5_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe5_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe5_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe5_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe5_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe5_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe5_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe5_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe5_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe5_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe5_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe5_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe5_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe5_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe5_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe5_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe5_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe5_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe5_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe5_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe5_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe5_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe5_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe5_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe5_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe5_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe5_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe5_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe5_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe5_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe5_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe5_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe5_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe5_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe5_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe5_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe5_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe5_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe5_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe5_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe5_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe5_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe5_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe5_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe5_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe5_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe5_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe5_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe5_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe5_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe5_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe5_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe5_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe5_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe5_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe5_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe5_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe5_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe5_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe5_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe5_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe5_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe5_io_pipe_phv_out_is_valid_processor),
    .io_vliw_in_0(pipe5_io_vliw_in_0),
    .io_vliw_in_1(pipe5_io_vliw_in_1),
    .io_vliw_in_2(pipe5_io_vliw_in_2),
    .io_vliw_in_3(pipe5_io_vliw_in_3),
    .io_field_in_0(pipe5_io_field_in_0),
    .io_field_in_1(pipe5_io_field_in_1),
    .io_field_in_2(pipe5_io_field_in_2),
    .io_field_in_3(pipe5_io_field_in_3),
    .io_offset_out_0(pipe5_io_offset_out_0),
    .io_offset_out_1(pipe5_io_offset_out_1),
    .io_offset_out_2(pipe5_io_offset_out_2),
    .io_offset_out_3(pipe5_io_offset_out_3),
    .io_length_out_0(pipe5_io_length_out_0),
    .io_length_out_1(pipe5_io_length_out_1),
    .io_length_out_2(pipe5_io_length_out_2),
    .io_length_out_3(pipe5_io_length_out_3),
    .io_field_out_0(pipe5_io_field_out_0),
    .io_field_out_1(pipe5_io_field_out_1),
    .io_field_out_2(pipe5_io_field_out_2),
    .io_field_out_3(pipe5_io_field_out_3)
  );
  PrimitiveWriteBack pipe6 ( // @[executor.scala 322:23]
    .clock(pipe6_clock),
    .io_pipe_phv_in_data_0(pipe6_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe6_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe6_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe6_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe6_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe6_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe6_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe6_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe6_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe6_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe6_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe6_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe6_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe6_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe6_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe6_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe6_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe6_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe6_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe6_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe6_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe6_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe6_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe6_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe6_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe6_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe6_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe6_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe6_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe6_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe6_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe6_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe6_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe6_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe6_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe6_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe6_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe6_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe6_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe6_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe6_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe6_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe6_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe6_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe6_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe6_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe6_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe6_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe6_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe6_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe6_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe6_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe6_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe6_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe6_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe6_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe6_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe6_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe6_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe6_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe6_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe6_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe6_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe6_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe6_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe6_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe6_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe6_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe6_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe6_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe6_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe6_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe6_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe6_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe6_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe6_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe6_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe6_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe6_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe6_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe6_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe6_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe6_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe6_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe6_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe6_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe6_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe6_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe6_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe6_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe6_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe6_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe6_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe6_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe6_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe6_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe6_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe6_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe6_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe6_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe6_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe6_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe6_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe6_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe6_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe6_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe6_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe6_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe6_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe6_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe6_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe6_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe6_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe6_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe6_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe6_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe6_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe6_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe6_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe6_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe6_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe6_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe6_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe6_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe6_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe6_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe6_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe6_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe6_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe6_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe6_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe6_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe6_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe6_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe6_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe6_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe6_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe6_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe6_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe6_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe6_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe6_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe6_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe6_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe6_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe6_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe6_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe6_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe6_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe6_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe6_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe6_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe6_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe6_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe6_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe6_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe6_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe6_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe6_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe6_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe6_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe6_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe6_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe6_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe6_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe6_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe6_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe6_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe6_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe6_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe6_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe6_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe6_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe6_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe6_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe6_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe6_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe6_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe6_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe6_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe6_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe6_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe6_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe6_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe6_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe6_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe6_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe6_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe6_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe6_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe6_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe6_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe6_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe6_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe6_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe6_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe6_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe6_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe6_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe6_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe6_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe6_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe6_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe6_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe6_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe6_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe6_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe6_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe6_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe6_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe6_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe6_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe6_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe6_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe6_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe6_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe6_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe6_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe6_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe6_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe6_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe6_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe6_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe6_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe6_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe6_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe6_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe6_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe6_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe6_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe6_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe6_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe6_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe6_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe6_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe6_io_pipe_phv_out_is_valid_processor),
    .io_offset_in_0(pipe6_io_offset_in_0),
    .io_offset_in_1(pipe6_io_offset_in_1),
    .io_offset_in_2(pipe6_io_offset_in_2),
    .io_offset_in_3(pipe6_io_offset_in_3),
    .io_length_in_0(pipe6_io_length_in_0),
    .io_length_in_1(pipe6_io_length_in_1),
    .io_length_in_2(pipe6_io_length_in_2),
    .io_length_in_3(pipe6_io_length_in_3),
    .io_field_in_0(pipe6_io_field_in_0),
    .io_field_in_1(pipe6_io_field_in_1),
    .io_field_in_2(pipe6_io_field_in_2),
    .io_field_in_3(pipe6_io_field_in_3)
  );
  assign io_pipe_phv_out_data_0 = pipe6_io_pipe_phv_out_data_0; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_1 = pipe6_io_pipe_phv_out_data_1; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_2 = pipe6_io_pipe_phv_out_data_2; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_3 = pipe6_io_pipe_phv_out_data_3; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_4 = pipe6_io_pipe_phv_out_data_4; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_5 = pipe6_io_pipe_phv_out_data_5; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_6 = pipe6_io_pipe_phv_out_data_6; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_7 = pipe6_io_pipe_phv_out_data_7; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_8 = pipe6_io_pipe_phv_out_data_8; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_9 = pipe6_io_pipe_phv_out_data_9; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_10 = pipe6_io_pipe_phv_out_data_10; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_11 = pipe6_io_pipe_phv_out_data_11; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_12 = pipe6_io_pipe_phv_out_data_12; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_13 = pipe6_io_pipe_phv_out_data_13; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_14 = pipe6_io_pipe_phv_out_data_14; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_15 = pipe6_io_pipe_phv_out_data_15; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_16 = pipe6_io_pipe_phv_out_data_16; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_17 = pipe6_io_pipe_phv_out_data_17; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_18 = pipe6_io_pipe_phv_out_data_18; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_19 = pipe6_io_pipe_phv_out_data_19; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_20 = pipe6_io_pipe_phv_out_data_20; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_21 = pipe6_io_pipe_phv_out_data_21; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_22 = pipe6_io_pipe_phv_out_data_22; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_23 = pipe6_io_pipe_phv_out_data_23; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_24 = pipe6_io_pipe_phv_out_data_24; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_25 = pipe6_io_pipe_phv_out_data_25; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_26 = pipe6_io_pipe_phv_out_data_26; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_27 = pipe6_io_pipe_phv_out_data_27; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_28 = pipe6_io_pipe_phv_out_data_28; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_29 = pipe6_io_pipe_phv_out_data_29; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_30 = pipe6_io_pipe_phv_out_data_30; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_31 = pipe6_io_pipe_phv_out_data_31; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_32 = pipe6_io_pipe_phv_out_data_32; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_33 = pipe6_io_pipe_phv_out_data_33; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_34 = pipe6_io_pipe_phv_out_data_34; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_35 = pipe6_io_pipe_phv_out_data_35; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_36 = pipe6_io_pipe_phv_out_data_36; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_37 = pipe6_io_pipe_phv_out_data_37; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_38 = pipe6_io_pipe_phv_out_data_38; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_39 = pipe6_io_pipe_phv_out_data_39; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_40 = pipe6_io_pipe_phv_out_data_40; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_41 = pipe6_io_pipe_phv_out_data_41; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_42 = pipe6_io_pipe_phv_out_data_42; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_43 = pipe6_io_pipe_phv_out_data_43; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_44 = pipe6_io_pipe_phv_out_data_44; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_45 = pipe6_io_pipe_phv_out_data_45; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_46 = pipe6_io_pipe_phv_out_data_46; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_47 = pipe6_io_pipe_phv_out_data_47; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_48 = pipe6_io_pipe_phv_out_data_48; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_49 = pipe6_io_pipe_phv_out_data_49; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_50 = pipe6_io_pipe_phv_out_data_50; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_51 = pipe6_io_pipe_phv_out_data_51; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_52 = pipe6_io_pipe_phv_out_data_52; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_53 = pipe6_io_pipe_phv_out_data_53; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_54 = pipe6_io_pipe_phv_out_data_54; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_55 = pipe6_io_pipe_phv_out_data_55; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_56 = pipe6_io_pipe_phv_out_data_56; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_57 = pipe6_io_pipe_phv_out_data_57; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_58 = pipe6_io_pipe_phv_out_data_58; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_59 = pipe6_io_pipe_phv_out_data_59; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_60 = pipe6_io_pipe_phv_out_data_60; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_61 = pipe6_io_pipe_phv_out_data_61; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_62 = pipe6_io_pipe_phv_out_data_62; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_63 = pipe6_io_pipe_phv_out_data_63; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_64 = pipe6_io_pipe_phv_out_data_64; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_65 = pipe6_io_pipe_phv_out_data_65; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_66 = pipe6_io_pipe_phv_out_data_66; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_67 = pipe6_io_pipe_phv_out_data_67; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_68 = pipe6_io_pipe_phv_out_data_68; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_69 = pipe6_io_pipe_phv_out_data_69; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_70 = pipe6_io_pipe_phv_out_data_70; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_71 = pipe6_io_pipe_phv_out_data_71; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_72 = pipe6_io_pipe_phv_out_data_72; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_73 = pipe6_io_pipe_phv_out_data_73; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_74 = pipe6_io_pipe_phv_out_data_74; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_75 = pipe6_io_pipe_phv_out_data_75; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_76 = pipe6_io_pipe_phv_out_data_76; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_77 = pipe6_io_pipe_phv_out_data_77; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_78 = pipe6_io_pipe_phv_out_data_78; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_79 = pipe6_io_pipe_phv_out_data_79; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_80 = pipe6_io_pipe_phv_out_data_80; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_81 = pipe6_io_pipe_phv_out_data_81; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_82 = pipe6_io_pipe_phv_out_data_82; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_83 = pipe6_io_pipe_phv_out_data_83; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_84 = pipe6_io_pipe_phv_out_data_84; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_85 = pipe6_io_pipe_phv_out_data_85; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_86 = pipe6_io_pipe_phv_out_data_86; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_87 = pipe6_io_pipe_phv_out_data_87; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_88 = pipe6_io_pipe_phv_out_data_88; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_89 = pipe6_io_pipe_phv_out_data_89; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_90 = pipe6_io_pipe_phv_out_data_90; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_91 = pipe6_io_pipe_phv_out_data_91; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_92 = pipe6_io_pipe_phv_out_data_92; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_93 = pipe6_io_pipe_phv_out_data_93; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_94 = pipe6_io_pipe_phv_out_data_94; // @[executor.scala 352:27]
  assign io_pipe_phv_out_data_95 = pipe6_io_pipe_phv_out_data_95; // @[executor.scala 352:27]
  assign io_pipe_phv_out_header_0 = pipe6_io_pipe_phv_out_header_0; // @[executor.scala 352:27]
  assign io_pipe_phv_out_header_1 = pipe6_io_pipe_phv_out_header_1; // @[executor.scala 352:27]
  assign io_pipe_phv_out_header_2 = pipe6_io_pipe_phv_out_header_2; // @[executor.scala 352:27]
  assign io_pipe_phv_out_header_3 = pipe6_io_pipe_phv_out_header_3; // @[executor.scala 352:27]
  assign io_pipe_phv_out_header_4 = pipe6_io_pipe_phv_out_header_4; // @[executor.scala 352:27]
  assign io_pipe_phv_out_header_5 = pipe6_io_pipe_phv_out_header_5; // @[executor.scala 352:27]
  assign io_pipe_phv_out_header_6 = pipe6_io_pipe_phv_out_header_6; // @[executor.scala 352:27]
  assign io_pipe_phv_out_header_7 = pipe6_io_pipe_phv_out_header_7; // @[executor.scala 352:27]
  assign io_pipe_phv_out_header_8 = pipe6_io_pipe_phv_out_header_8; // @[executor.scala 352:27]
  assign io_pipe_phv_out_header_9 = pipe6_io_pipe_phv_out_header_9; // @[executor.scala 352:27]
  assign io_pipe_phv_out_header_10 = pipe6_io_pipe_phv_out_header_10; // @[executor.scala 352:27]
  assign io_pipe_phv_out_header_11 = pipe6_io_pipe_phv_out_header_11; // @[executor.scala 352:27]
  assign io_pipe_phv_out_header_12 = pipe6_io_pipe_phv_out_header_12; // @[executor.scala 352:27]
  assign io_pipe_phv_out_header_13 = pipe6_io_pipe_phv_out_header_13; // @[executor.scala 352:27]
  assign io_pipe_phv_out_header_14 = pipe6_io_pipe_phv_out_header_14; // @[executor.scala 352:27]
  assign io_pipe_phv_out_header_15 = pipe6_io_pipe_phv_out_header_15; // @[executor.scala 352:27]
  assign io_pipe_phv_out_parse_current_state = pipe6_io_pipe_phv_out_parse_current_state; // @[executor.scala 352:27]
  assign io_pipe_phv_out_parse_current_offset = pipe6_io_pipe_phv_out_parse_current_offset; // @[executor.scala 352:27]
  assign io_pipe_phv_out_parse_transition_field = pipe6_io_pipe_phv_out_parse_transition_field; // @[executor.scala 352:27]
  assign io_pipe_phv_out_next_processor_id = pipe6_io_pipe_phv_out_next_processor_id; // @[executor.scala 352:27]
  assign io_pipe_phv_out_next_config_id = pipe6_io_pipe_phv_out_next_config_id; // @[executor.scala 352:27]
  assign io_pipe_phv_out_is_valid_processor = pipe6_io_pipe_phv_out_is_valid_processor; // @[executor.scala 352:27]
  assign pipe1_clock = clock;
  assign pipe1_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[executor.scala 324:26]
  assign pipe1_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[executor.scala 324:26]
  assign pipe1_io_hit = io_hit; // @[executor.scala 325:26]
  assign pipe1_io_match_value = io_match_value; // @[executor.scala 326:26]
  assign pipe1_io_action_mod_en = io_action_mod_en; // @[executor.scala 327:26]
  assign pipe1_io_action_mod_addr = io_action_mod_addr; // @[executor.scala 327:26]
  assign pipe1_io_action_mod_data_0 = io_action_mod_data_0; // @[executor.scala 327:26]
  assign pipe1_io_action_mod_data_1 = io_action_mod_data_1; // @[executor.scala 327:26]
  assign pipe2_clock = clock;
  assign pipe2_io_pipe_phv_in_data_0 = pipe1_io_pipe_phv_out_data_0; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_1 = pipe1_io_pipe_phv_out_data_1; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_2 = pipe1_io_pipe_phv_out_data_2; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_3 = pipe1_io_pipe_phv_out_data_3; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_4 = pipe1_io_pipe_phv_out_data_4; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_5 = pipe1_io_pipe_phv_out_data_5; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_6 = pipe1_io_pipe_phv_out_data_6; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_7 = pipe1_io_pipe_phv_out_data_7; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_8 = pipe1_io_pipe_phv_out_data_8; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_9 = pipe1_io_pipe_phv_out_data_9; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_10 = pipe1_io_pipe_phv_out_data_10; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_11 = pipe1_io_pipe_phv_out_data_11; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_12 = pipe1_io_pipe_phv_out_data_12; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_13 = pipe1_io_pipe_phv_out_data_13; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_14 = pipe1_io_pipe_phv_out_data_14; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_15 = pipe1_io_pipe_phv_out_data_15; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_16 = pipe1_io_pipe_phv_out_data_16; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_17 = pipe1_io_pipe_phv_out_data_17; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_18 = pipe1_io_pipe_phv_out_data_18; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_19 = pipe1_io_pipe_phv_out_data_19; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_20 = pipe1_io_pipe_phv_out_data_20; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_21 = pipe1_io_pipe_phv_out_data_21; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_22 = pipe1_io_pipe_phv_out_data_22; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_23 = pipe1_io_pipe_phv_out_data_23; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_24 = pipe1_io_pipe_phv_out_data_24; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_25 = pipe1_io_pipe_phv_out_data_25; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_26 = pipe1_io_pipe_phv_out_data_26; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_27 = pipe1_io_pipe_phv_out_data_27; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_28 = pipe1_io_pipe_phv_out_data_28; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_29 = pipe1_io_pipe_phv_out_data_29; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_30 = pipe1_io_pipe_phv_out_data_30; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_31 = pipe1_io_pipe_phv_out_data_31; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_32 = pipe1_io_pipe_phv_out_data_32; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_33 = pipe1_io_pipe_phv_out_data_33; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_34 = pipe1_io_pipe_phv_out_data_34; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_35 = pipe1_io_pipe_phv_out_data_35; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_36 = pipe1_io_pipe_phv_out_data_36; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_37 = pipe1_io_pipe_phv_out_data_37; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_38 = pipe1_io_pipe_phv_out_data_38; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_39 = pipe1_io_pipe_phv_out_data_39; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_40 = pipe1_io_pipe_phv_out_data_40; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_41 = pipe1_io_pipe_phv_out_data_41; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_42 = pipe1_io_pipe_phv_out_data_42; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_43 = pipe1_io_pipe_phv_out_data_43; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_44 = pipe1_io_pipe_phv_out_data_44; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_45 = pipe1_io_pipe_phv_out_data_45; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_46 = pipe1_io_pipe_phv_out_data_46; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_47 = pipe1_io_pipe_phv_out_data_47; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_48 = pipe1_io_pipe_phv_out_data_48; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_49 = pipe1_io_pipe_phv_out_data_49; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_50 = pipe1_io_pipe_phv_out_data_50; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_51 = pipe1_io_pipe_phv_out_data_51; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_52 = pipe1_io_pipe_phv_out_data_52; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_53 = pipe1_io_pipe_phv_out_data_53; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_54 = pipe1_io_pipe_phv_out_data_54; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_55 = pipe1_io_pipe_phv_out_data_55; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_56 = pipe1_io_pipe_phv_out_data_56; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_57 = pipe1_io_pipe_phv_out_data_57; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_58 = pipe1_io_pipe_phv_out_data_58; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_59 = pipe1_io_pipe_phv_out_data_59; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_60 = pipe1_io_pipe_phv_out_data_60; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_61 = pipe1_io_pipe_phv_out_data_61; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_62 = pipe1_io_pipe_phv_out_data_62; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_63 = pipe1_io_pipe_phv_out_data_63; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_64 = pipe1_io_pipe_phv_out_data_64; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_65 = pipe1_io_pipe_phv_out_data_65; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_66 = pipe1_io_pipe_phv_out_data_66; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_67 = pipe1_io_pipe_phv_out_data_67; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_68 = pipe1_io_pipe_phv_out_data_68; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_69 = pipe1_io_pipe_phv_out_data_69; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_70 = pipe1_io_pipe_phv_out_data_70; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_71 = pipe1_io_pipe_phv_out_data_71; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_72 = pipe1_io_pipe_phv_out_data_72; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_73 = pipe1_io_pipe_phv_out_data_73; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_74 = pipe1_io_pipe_phv_out_data_74; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_75 = pipe1_io_pipe_phv_out_data_75; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_76 = pipe1_io_pipe_phv_out_data_76; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_77 = pipe1_io_pipe_phv_out_data_77; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_78 = pipe1_io_pipe_phv_out_data_78; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_79 = pipe1_io_pipe_phv_out_data_79; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_80 = pipe1_io_pipe_phv_out_data_80; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_81 = pipe1_io_pipe_phv_out_data_81; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_82 = pipe1_io_pipe_phv_out_data_82; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_83 = pipe1_io_pipe_phv_out_data_83; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_84 = pipe1_io_pipe_phv_out_data_84; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_85 = pipe1_io_pipe_phv_out_data_85; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_86 = pipe1_io_pipe_phv_out_data_86; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_87 = pipe1_io_pipe_phv_out_data_87; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_88 = pipe1_io_pipe_phv_out_data_88; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_89 = pipe1_io_pipe_phv_out_data_89; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_90 = pipe1_io_pipe_phv_out_data_90; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_91 = pipe1_io_pipe_phv_out_data_91; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_92 = pipe1_io_pipe_phv_out_data_92; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_93 = pipe1_io_pipe_phv_out_data_93; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_94 = pipe1_io_pipe_phv_out_data_94; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_data_95 = pipe1_io_pipe_phv_out_data_95; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_header_0 = pipe1_io_pipe_phv_out_header_0; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_header_1 = pipe1_io_pipe_phv_out_header_1; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_header_2 = pipe1_io_pipe_phv_out_header_2; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_header_3 = pipe1_io_pipe_phv_out_header_3; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_header_4 = pipe1_io_pipe_phv_out_header_4; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_header_5 = pipe1_io_pipe_phv_out_header_5; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_header_6 = pipe1_io_pipe_phv_out_header_6; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_header_7 = pipe1_io_pipe_phv_out_header_7; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_header_8 = pipe1_io_pipe_phv_out_header_8; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_header_9 = pipe1_io_pipe_phv_out_header_9; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_header_10 = pipe1_io_pipe_phv_out_header_10; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_header_11 = pipe1_io_pipe_phv_out_header_11; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_header_12 = pipe1_io_pipe_phv_out_header_12; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_header_13 = pipe1_io_pipe_phv_out_header_13; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_header_14 = pipe1_io_pipe_phv_out_header_14; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_header_15 = pipe1_io_pipe_phv_out_header_15; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_parse_current_state = pipe1_io_pipe_phv_out_parse_current_state; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_parse_current_offset = pipe1_io_pipe_phv_out_parse_current_offset; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_parse_transition_field = pipe1_io_pipe_phv_out_parse_transition_field; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_next_processor_id = pipe1_io_pipe_phv_out_next_processor_id; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_next_config_id = pipe1_io_pipe_phv_out_next_config_id; // @[executor.scala 329:26]
  assign pipe2_io_pipe_phv_in_is_valid_processor = pipe1_io_pipe_phv_out_is_valid_processor; // @[executor.scala 329:26]
  assign pipe2_io_args_in_0 = pipe1_io_args_out_0; // @[executor.scala 330:26]
  assign pipe2_io_args_in_1 = pipe1_io_args_out_1; // @[executor.scala 330:26]
  assign pipe2_io_args_in_2 = pipe1_io_args_out_2; // @[executor.scala 330:26]
  assign pipe2_io_args_in_3 = pipe1_io_args_out_3; // @[executor.scala 330:26]
  assign pipe2_io_args_in_4 = pipe1_io_args_out_4; // @[executor.scala 330:26]
  assign pipe2_io_args_in_5 = pipe1_io_args_out_5; // @[executor.scala 330:26]
  assign pipe2_io_args_in_6 = pipe1_io_args_out_6; // @[executor.scala 330:26]
  assign pipe2_io_vliw_in_0 = pipe1_io_vliw_out_0; // @[executor.scala 331:26]
  assign pipe2_io_vliw_in_1 = pipe1_io_vliw_out_1; // @[executor.scala 331:26]
  assign pipe2_io_vliw_in_2 = pipe1_io_vliw_out_2; // @[executor.scala 331:26]
  assign pipe2_io_vliw_in_3 = pipe1_io_vliw_out_3; // @[executor.scala 331:26]
  assign pipe3_clock = clock;
  assign pipe3_io_pipe_phv_in_data_0 = pipe2_io_pipe_phv_out_data_0; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_1 = pipe2_io_pipe_phv_out_data_1; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_2 = pipe2_io_pipe_phv_out_data_2; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_3 = pipe2_io_pipe_phv_out_data_3; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_4 = pipe2_io_pipe_phv_out_data_4; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_5 = pipe2_io_pipe_phv_out_data_5; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_6 = pipe2_io_pipe_phv_out_data_6; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_7 = pipe2_io_pipe_phv_out_data_7; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_8 = pipe2_io_pipe_phv_out_data_8; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_9 = pipe2_io_pipe_phv_out_data_9; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_10 = pipe2_io_pipe_phv_out_data_10; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_11 = pipe2_io_pipe_phv_out_data_11; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_12 = pipe2_io_pipe_phv_out_data_12; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_13 = pipe2_io_pipe_phv_out_data_13; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_14 = pipe2_io_pipe_phv_out_data_14; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_15 = pipe2_io_pipe_phv_out_data_15; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_16 = pipe2_io_pipe_phv_out_data_16; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_17 = pipe2_io_pipe_phv_out_data_17; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_18 = pipe2_io_pipe_phv_out_data_18; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_19 = pipe2_io_pipe_phv_out_data_19; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_20 = pipe2_io_pipe_phv_out_data_20; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_21 = pipe2_io_pipe_phv_out_data_21; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_22 = pipe2_io_pipe_phv_out_data_22; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_23 = pipe2_io_pipe_phv_out_data_23; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_24 = pipe2_io_pipe_phv_out_data_24; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_25 = pipe2_io_pipe_phv_out_data_25; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_26 = pipe2_io_pipe_phv_out_data_26; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_27 = pipe2_io_pipe_phv_out_data_27; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_28 = pipe2_io_pipe_phv_out_data_28; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_29 = pipe2_io_pipe_phv_out_data_29; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_30 = pipe2_io_pipe_phv_out_data_30; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_31 = pipe2_io_pipe_phv_out_data_31; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_32 = pipe2_io_pipe_phv_out_data_32; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_33 = pipe2_io_pipe_phv_out_data_33; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_34 = pipe2_io_pipe_phv_out_data_34; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_35 = pipe2_io_pipe_phv_out_data_35; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_36 = pipe2_io_pipe_phv_out_data_36; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_37 = pipe2_io_pipe_phv_out_data_37; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_38 = pipe2_io_pipe_phv_out_data_38; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_39 = pipe2_io_pipe_phv_out_data_39; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_40 = pipe2_io_pipe_phv_out_data_40; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_41 = pipe2_io_pipe_phv_out_data_41; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_42 = pipe2_io_pipe_phv_out_data_42; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_43 = pipe2_io_pipe_phv_out_data_43; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_44 = pipe2_io_pipe_phv_out_data_44; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_45 = pipe2_io_pipe_phv_out_data_45; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_46 = pipe2_io_pipe_phv_out_data_46; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_47 = pipe2_io_pipe_phv_out_data_47; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_48 = pipe2_io_pipe_phv_out_data_48; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_49 = pipe2_io_pipe_phv_out_data_49; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_50 = pipe2_io_pipe_phv_out_data_50; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_51 = pipe2_io_pipe_phv_out_data_51; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_52 = pipe2_io_pipe_phv_out_data_52; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_53 = pipe2_io_pipe_phv_out_data_53; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_54 = pipe2_io_pipe_phv_out_data_54; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_55 = pipe2_io_pipe_phv_out_data_55; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_56 = pipe2_io_pipe_phv_out_data_56; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_57 = pipe2_io_pipe_phv_out_data_57; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_58 = pipe2_io_pipe_phv_out_data_58; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_59 = pipe2_io_pipe_phv_out_data_59; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_60 = pipe2_io_pipe_phv_out_data_60; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_61 = pipe2_io_pipe_phv_out_data_61; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_62 = pipe2_io_pipe_phv_out_data_62; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_63 = pipe2_io_pipe_phv_out_data_63; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_64 = pipe2_io_pipe_phv_out_data_64; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_65 = pipe2_io_pipe_phv_out_data_65; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_66 = pipe2_io_pipe_phv_out_data_66; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_67 = pipe2_io_pipe_phv_out_data_67; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_68 = pipe2_io_pipe_phv_out_data_68; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_69 = pipe2_io_pipe_phv_out_data_69; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_70 = pipe2_io_pipe_phv_out_data_70; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_71 = pipe2_io_pipe_phv_out_data_71; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_72 = pipe2_io_pipe_phv_out_data_72; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_73 = pipe2_io_pipe_phv_out_data_73; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_74 = pipe2_io_pipe_phv_out_data_74; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_75 = pipe2_io_pipe_phv_out_data_75; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_76 = pipe2_io_pipe_phv_out_data_76; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_77 = pipe2_io_pipe_phv_out_data_77; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_78 = pipe2_io_pipe_phv_out_data_78; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_79 = pipe2_io_pipe_phv_out_data_79; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_80 = pipe2_io_pipe_phv_out_data_80; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_81 = pipe2_io_pipe_phv_out_data_81; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_82 = pipe2_io_pipe_phv_out_data_82; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_83 = pipe2_io_pipe_phv_out_data_83; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_84 = pipe2_io_pipe_phv_out_data_84; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_85 = pipe2_io_pipe_phv_out_data_85; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_86 = pipe2_io_pipe_phv_out_data_86; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_87 = pipe2_io_pipe_phv_out_data_87; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_88 = pipe2_io_pipe_phv_out_data_88; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_89 = pipe2_io_pipe_phv_out_data_89; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_90 = pipe2_io_pipe_phv_out_data_90; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_91 = pipe2_io_pipe_phv_out_data_91; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_92 = pipe2_io_pipe_phv_out_data_92; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_93 = pipe2_io_pipe_phv_out_data_93; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_94 = pipe2_io_pipe_phv_out_data_94; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_data_95 = pipe2_io_pipe_phv_out_data_95; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_header_0 = pipe2_io_pipe_phv_out_header_0; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_header_1 = pipe2_io_pipe_phv_out_header_1; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_header_2 = pipe2_io_pipe_phv_out_header_2; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_header_3 = pipe2_io_pipe_phv_out_header_3; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_header_4 = pipe2_io_pipe_phv_out_header_4; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_header_5 = pipe2_io_pipe_phv_out_header_5; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_header_6 = pipe2_io_pipe_phv_out_header_6; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_header_7 = pipe2_io_pipe_phv_out_header_7; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_header_8 = pipe2_io_pipe_phv_out_header_8; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_header_9 = pipe2_io_pipe_phv_out_header_9; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_header_10 = pipe2_io_pipe_phv_out_header_10; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_header_11 = pipe2_io_pipe_phv_out_header_11; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_header_12 = pipe2_io_pipe_phv_out_header_12; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_header_13 = pipe2_io_pipe_phv_out_header_13; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_header_14 = pipe2_io_pipe_phv_out_header_14; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_header_15 = pipe2_io_pipe_phv_out_header_15; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_parse_current_state = pipe2_io_pipe_phv_out_parse_current_state; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_parse_current_offset = pipe2_io_pipe_phv_out_parse_current_offset; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_parse_transition_field = pipe2_io_pipe_phv_out_parse_transition_field; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_next_processor_id = pipe2_io_pipe_phv_out_next_processor_id; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_next_config_id = pipe2_io_pipe_phv_out_next_config_id; // @[executor.scala 333:26]
  assign pipe3_io_pipe_phv_in_is_valid_processor = pipe2_io_pipe_phv_out_is_valid_processor; // @[executor.scala 333:26]
  assign pipe3_io_args_in_0 = pipe2_io_args_out_0; // @[executor.scala 334:26]
  assign pipe3_io_args_in_1 = pipe2_io_args_out_1; // @[executor.scala 334:26]
  assign pipe3_io_args_in_2 = pipe2_io_args_out_2; // @[executor.scala 334:26]
  assign pipe3_io_args_in_3 = pipe2_io_args_out_3; // @[executor.scala 334:26]
  assign pipe3_io_args_in_4 = pipe2_io_args_out_4; // @[executor.scala 334:26]
  assign pipe3_io_args_in_5 = pipe2_io_args_out_5; // @[executor.scala 334:26]
  assign pipe3_io_args_in_6 = pipe2_io_args_out_6; // @[executor.scala 334:26]
  assign pipe3_io_vliw_in_0 = pipe2_io_vliw_out_0; // @[executor.scala 335:26]
  assign pipe3_io_vliw_in_1 = pipe2_io_vliw_out_1; // @[executor.scala 335:26]
  assign pipe3_io_vliw_in_2 = pipe2_io_vliw_out_2; // @[executor.scala 335:26]
  assign pipe3_io_vliw_in_3 = pipe2_io_vliw_out_3; // @[executor.scala 335:26]
  assign pipe3_io_offset_in_0 = pipe2_io_offset_out_0; // @[executor.scala 336:26]
  assign pipe3_io_offset_in_1 = pipe2_io_offset_out_1; // @[executor.scala 336:26]
  assign pipe3_io_offset_in_2 = pipe2_io_offset_out_2; // @[executor.scala 336:26]
  assign pipe3_io_offset_in_3 = pipe2_io_offset_out_3; // @[executor.scala 336:26]
  assign pipe3_io_length_in_0 = pipe2_io_length_out_0; // @[executor.scala 337:26]
  assign pipe3_io_length_in_1 = pipe2_io_length_out_1; // @[executor.scala 337:26]
  assign pipe3_io_length_in_2 = pipe2_io_length_out_2; // @[executor.scala 337:26]
  assign pipe3_io_length_in_3 = pipe2_io_length_out_3; // @[executor.scala 337:26]
  assign pipe4_clock = clock;
  assign pipe4_io_pipe_phv_in_data_0 = pipe3_io_pipe_phv_out_data_0; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_1 = pipe3_io_pipe_phv_out_data_1; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_2 = pipe3_io_pipe_phv_out_data_2; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_3 = pipe3_io_pipe_phv_out_data_3; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_4 = pipe3_io_pipe_phv_out_data_4; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_5 = pipe3_io_pipe_phv_out_data_5; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_6 = pipe3_io_pipe_phv_out_data_6; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_7 = pipe3_io_pipe_phv_out_data_7; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_8 = pipe3_io_pipe_phv_out_data_8; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_9 = pipe3_io_pipe_phv_out_data_9; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_10 = pipe3_io_pipe_phv_out_data_10; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_11 = pipe3_io_pipe_phv_out_data_11; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_12 = pipe3_io_pipe_phv_out_data_12; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_13 = pipe3_io_pipe_phv_out_data_13; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_14 = pipe3_io_pipe_phv_out_data_14; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_15 = pipe3_io_pipe_phv_out_data_15; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_16 = pipe3_io_pipe_phv_out_data_16; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_17 = pipe3_io_pipe_phv_out_data_17; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_18 = pipe3_io_pipe_phv_out_data_18; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_19 = pipe3_io_pipe_phv_out_data_19; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_20 = pipe3_io_pipe_phv_out_data_20; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_21 = pipe3_io_pipe_phv_out_data_21; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_22 = pipe3_io_pipe_phv_out_data_22; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_23 = pipe3_io_pipe_phv_out_data_23; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_24 = pipe3_io_pipe_phv_out_data_24; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_25 = pipe3_io_pipe_phv_out_data_25; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_26 = pipe3_io_pipe_phv_out_data_26; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_27 = pipe3_io_pipe_phv_out_data_27; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_28 = pipe3_io_pipe_phv_out_data_28; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_29 = pipe3_io_pipe_phv_out_data_29; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_30 = pipe3_io_pipe_phv_out_data_30; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_31 = pipe3_io_pipe_phv_out_data_31; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_32 = pipe3_io_pipe_phv_out_data_32; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_33 = pipe3_io_pipe_phv_out_data_33; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_34 = pipe3_io_pipe_phv_out_data_34; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_35 = pipe3_io_pipe_phv_out_data_35; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_36 = pipe3_io_pipe_phv_out_data_36; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_37 = pipe3_io_pipe_phv_out_data_37; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_38 = pipe3_io_pipe_phv_out_data_38; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_39 = pipe3_io_pipe_phv_out_data_39; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_40 = pipe3_io_pipe_phv_out_data_40; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_41 = pipe3_io_pipe_phv_out_data_41; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_42 = pipe3_io_pipe_phv_out_data_42; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_43 = pipe3_io_pipe_phv_out_data_43; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_44 = pipe3_io_pipe_phv_out_data_44; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_45 = pipe3_io_pipe_phv_out_data_45; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_46 = pipe3_io_pipe_phv_out_data_46; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_47 = pipe3_io_pipe_phv_out_data_47; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_48 = pipe3_io_pipe_phv_out_data_48; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_49 = pipe3_io_pipe_phv_out_data_49; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_50 = pipe3_io_pipe_phv_out_data_50; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_51 = pipe3_io_pipe_phv_out_data_51; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_52 = pipe3_io_pipe_phv_out_data_52; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_53 = pipe3_io_pipe_phv_out_data_53; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_54 = pipe3_io_pipe_phv_out_data_54; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_55 = pipe3_io_pipe_phv_out_data_55; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_56 = pipe3_io_pipe_phv_out_data_56; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_57 = pipe3_io_pipe_phv_out_data_57; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_58 = pipe3_io_pipe_phv_out_data_58; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_59 = pipe3_io_pipe_phv_out_data_59; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_60 = pipe3_io_pipe_phv_out_data_60; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_61 = pipe3_io_pipe_phv_out_data_61; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_62 = pipe3_io_pipe_phv_out_data_62; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_63 = pipe3_io_pipe_phv_out_data_63; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_64 = pipe3_io_pipe_phv_out_data_64; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_65 = pipe3_io_pipe_phv_out_data_65; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_66 = pipe3_io_pipe_phv_out_data_66; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_67 = pipe3_io_pipe_phv_out_data_67; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_68 = pipe3_io_pipe_phv_out_data_68; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_69 = pipe3_io_pipe_phv_out_data_69; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_70 = pipe3_io_pipe_phv_out_data_70; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_71 = pipe3_io_pipe_phv_out_data_71; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_72 = pipe3_io_pipe_phv_out_data_72; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_73 = pipe3_io_pipe_phv_out_data_73; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_74 = pipe3_io_pipe_phv_out_data_74; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_75 = pipe3_io_pipe_phv_out_data_75; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_76 = pipe3_io_pipe_phv_out_data_76; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_77 = pipe3_io_pipe_phv_out_data_77; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_78 = pipe3_io_pipe_phv_out_data_78; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_79 = pipe3_io_pipe_phv_out_data_79; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_80 = pipe3_io_pipe_phv_out_data_80; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_81 = pipe3_io_pipe_phv_out_data_81; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_82 = pipe3_io_pipe_phv_out_data_82; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_83 = pipe3_io_pipe_phv_out_data_83; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_84 = pipe3_io_pipe_phv_out_data_84; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_85 = pipe3_io_pipe_phv_out_data_85; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_86 = pipe3_io_pipe_phv_out_data_86; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_87 = pipe3_io_pipe_phv_out_data_87; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_88 = pipe3_io_pipe_phv_out_data_88; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_89 = pipe3_io_pipe_phv_out_data_89; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_90 = pipe3_io_pipe_phv_out_data_90; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_91 = pipe3_io_pipe_phv_out_data_91; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_92 = pipe3_io_pipe_phv_out_data_92; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_93 = pipe3_io_pipe_phv_out_data_93; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_94 = pipe3_io_pipe_phv_out_data_94; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_data_95 = pipe3_io_pipe_phv_out_data_95; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_header_0 = pipe3_io_pipe_phv_out_header_0; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_header_1 = pipe3_io_pipe_phv_out_header_1; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_header_2 = pipe3_io_pipe_phv_out_header_2; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_header_3 = pipe3_io_pipe_phv_out_header_3; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_header_4 = pipe3_io_pipe_phv_out_header_4; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_header_5 = pipe3_io_pipe_phv_out_header_5; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_header_6 = pipe3_io_pipe_phv_out_header_6; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_header_7 = pipe3_io_pipe_phv_out_header_7; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_header_8 = pipe3_io_pipe_phv_out_header_8; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_header_9 = pipe3_io_pipe_phv_out_header_9; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_header_10 = pipe3_io_pipe_phv_out_header_10; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_header_11 = pipe3_io_pipe_phv_out_header_11; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_header_12 = pipe3_io_pipe_phv_out_header_12; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_header_13 = pipe3_io_pipe_phv_out_header_13; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_header_14 = pipe3_io_pipe_phv_out_header_14; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_header_15 = pipe3_io_pipe_phv_out_header_15; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_parse_current_state = pipe3_io_pipe_phv_out_parse_current_state; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_parse_current_offset = pipe3_io_pipe_phv_out_parse_current_offset; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_parse_transition_field = pipe3_io_pipe_phv_out_parse_transition_field; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_next_processor_id = pipe3_io_pipe_phv_out_next_processor_id; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_next_config_id = pipe3_io_pipe_phv_out_next_config_id; // @[executor.scala 339:26]
  assign pipe4_io_pipe_phv_in_is_valid_processor = pipe3_io_pipe_phv_out_is_valid_processor; // @[executor.scala 339:26]
  assign pipe4_io_vliw_in_0 = pipe3_io_vliw_out_0; // @[executor.scala 340:26]
  assign pipe4_io_vliw_in_1 = pipe3_io_vliw_out_1; // @[executor.scala 340:26]
  assign pipe4_io_vliw_in_2 = pipe3_io_vliw_out_2; // @[executor.scala 340:26]
  assign pipe4_io_vliw_in_3 = pipe3_io_vliw_out_3; // @[executor.scala 340:26]
  assign pipe4_io_field_in_0 = pipe3_io_field_out_0; // @[executor.scala 341:26]
  assign pipe4_io_field_in_1 = pipe3_io_field_out_1; // @[executor.scala 341:26]
  assign pipe4_io_field_in_2 = pipe3_io_field_out_2; // @[executor.scala 341:26]
  assign pipe4_io_field_in_3 = pipe3_io_field_out_3; // @[executor.scala 341:26]
  assign pipe5_clock = clock;
  assign pipe5_io_pipe_phv_in_data_0 = pipe4_io_pipe_phv_out_data_0; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_1 = pipe4_io_pipe_phv_out_data_1; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_2 = pipe4_io_pipe_phv_out_data_2; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_3 = pipe4_io_pipe_phv_out_data_3; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_4 = pipe4_io_pipe_phv_out_data_4; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_5 = pipe4_io_pipe_phv_out_data_5; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_6 = pipe4_io_pipe_phv_out_data_6; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_7 = pipe4_io_pipe_phv_out_data_7; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_8 = pipe4_io_pipe_phv_out_data_8; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_9 = pipe4_io_pipe_phv_out_data_9; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_10 = pipe4_io_pipe_phv_out_data_10; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_11 = pipe4_io_pipe_phv_out_data_11; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_12 = pipe4_io_pipe_phv_out_data_12; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_13 = pipe4_io_pipe_phv_out_data_13; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_14 = pipe4_io_pipe_phv_out_data_14; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_15 = pipe4_io_pipe_phv_out_data_15; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_16 = pipe4_io_pipe_phv_out_data_16; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_17 = pipe4_io_pipe_phv_out_data_17; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_18 = pipe4_io_pipe_phv_out_data_18; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_19 = pipe4_io_pipe_phv_out_data_19; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_20 = pipe4_io_pipe_phv_out_data_20; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_21 = pipe4_io_pipe_phv_out_data_21; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_22 = pipe4_io_pipe_phv_out_data_22; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_23 = pipe4_io_pipe_phv_out_data_23; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_24 = pipe4_io_pipe_phv_out_data_24; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_25 = pipe4_io_pipe_phv_out_data_25; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_26 = pipe4_io_pipe_phv_out_data_26; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_27 = pipe4_io_pipe_phv_out_data_27; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_28 = pipe4_io_pipe_phv_out_data_28; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_29 = pipe4_io_pipe_phv_out_data_29; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_30 = pipe4_io_pipe_phv_out_data_30; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_31 = pipe4_io_pipe_phv_out_data_31; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_32 = pipe4_io_pipe_phv_out_data_32; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_33 = pipe4_io_pipe_phv_out_data_33; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_34 = pipe4_io_pipe_phv_out_data_34; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_35 = pipe4_io_pipe_phv_out_data_35; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_36 = pipe4_io_pipe_phv_out_data_36; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_37 = pipe4_io_pipe_phv_out_data_37; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_38 = pipe4_io_pipe_phv_out_data_38; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_39 = pipe4_io_pipe_phv_out_data_39; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_40 = pipe4_io_pipe_phv_out_data_40; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_41 = pipe4_io_pipe_phv_out_data_41; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_42 = pipe4_io_pipe_phv_out_data_42; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_43 = pipe4_io_pipe_phv_out_data_43; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_44 = pipe4_io_pipe_phv_out_data_44; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_45 = pipe4_io_pipe_phv_out_data_45; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_46 = pipe4_io_pipe_phv_out_data_46; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_47 = pipe4_io_pipe_phv_out_data_47; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_48 = pipe4_io_pipe_phv_out_data_48; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_49 = pipe4_io_pipe_phv_out_data_49; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_50 = pipe4_io_pipe_phv_out_data_50; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_51 = pipe4_io_pipe_phv_out_data_51; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_52 = pipe4_io_pipe_phv_out_data_52; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_53 = pipe4_io_pipe_phv_out_data_53; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_54 = pipe4_io_pipe_phv_out_data_54; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_55 = pipe4_io_pipe_phv_out_data_55; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_56 = pipe4_io_pipe_phv_out_data_56; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_57 = pipe4_io_pipe_phv_out_data_57; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_58 = pipe4_io_pipe_phv_out_data_58; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_59 = pipe4_io_pipe_phv_out_data_59; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_60 = pipe4_io_pipe_phv_out_data_60; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_61 = pipe4_io_pipe_phv_out_data_61; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_62 = pipe4_io_pipe_phv_out_data_62; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_63 = pipe4_io_pipe_phv_out_data_63; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_64 = pipe4_io_pipe_phv_out_data_64; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_65 = pipe4_io_pipe_phv_out_data_65; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_66 = pipe4_io_pipe_phv_out_data_66; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_67 = pipe4_io_pipe_phv_out_data_67; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_68 = pipe4_io_pipe_phv_out_data_68; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_69 = pipe4_io_pipe_phv_out_data_69; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_70 = pipe4_io_pipe_phv_out_data_70; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_71 = pipe4_io_pipe_phv_out_data_71; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_72 = pipe4_io_pipe_phv_out_data_72; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_73 = pipe4_io_pipe_phv_out_data_73; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_74 = pipe4_io_pipe_phv_out_data_74; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_75 = pipe4_io_pipe_phv_out_data_75; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_76 = pipe4_io_pipe_phv_out_data_76; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_77 = pipe4_io_pipe_phv_out_data_77; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_78 = pipe4_io_pipe_phv_out_data_78; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_79 = pipe4_io_pipe_phv_out_data_79; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_80 = pipe4_io_pipe_phv_out_data_80; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_81 = pipe4_io_pipe_phv_out_data_81; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_82 = pipe4_io_pipe_phv_out_data_82; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_83 = pipe4_io_pipe_phv_out_data_83; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_84 = pipe4_io_pipe_phv_out_data_84; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_85 = pipe4_io_pipe_phv_out_data_85; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_86 = pipe4_io_pipe_phv_out_data_86; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_87 = pipe4_io_pipe_phv_out_data_87; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_88 = pipe4_io_pipe_phv_out_data_88; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_89 = pipe4_io_pipe_phv_out_data_89; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_90 = pipe4_io_pipe_phv_out_data_90; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_91 = pipe4_io_pipe_phv_out_data_91; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_92 = pipe4_io_pipe_phv_out_data_92; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_93 = pipe4_io_pipe_phv_out_data_93; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_94 = pipe4_io_pipe_phv_out_data_94; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_data_95 = pipe4_io_pipe_phv_out_data_95; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_header_0 = pipe4_io_pipe_phv_out_header_0; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_header_1 = pipe4_io_pipe_phv_out_header_1; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_header_2 = pipe4_io_pipe_phv_out_header_2; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_header_3 = pipe4_io_pipe_phv_out_header_3; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_header_4 = pipe4_io_pipe_phv_out_header_4; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_header_5 = pipe4_io_pipe_phv_out_header_5; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_header_6 = pipe4_io_pipe_phv_out_header_6; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_header_7 = pipe4_io_pipe_phv_out_header_7; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_header_8 = pipe4_io_pipe_phv_out_header_8; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_header_9 = pipe4_io_pipe_phv_out_header_9; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_header_10 = pipe4_io_pipe_phv_out_header_10; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_header_11 = pipe4_io_pipe_phv_out_header_11; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_header_12 = pipe4_io_pipe_phv_out_header_12; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_header_13 = pipe4_io_pipe_phv_out_header_13; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_header_14 = pipe4_io_pipe_phv_out_header_14; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_header_15 = pipe4_io_pipe_phv_out_header_15; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_parse_current_state = pipe4_io_pipe_phv_out_parse_current_state; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_parse_current_offset = pipe4_io_pipe_phv_out_parse_current_offset; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_parse_transition_field = pipe4_io_pipe_phv_out_parse_transition_field; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_next_processor_id = pipe4_io_pipe_phv_out_next_processor_id; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_next_config_id = pipe4_io_pipe_phv_out_next_config_id; // @[executor.scala 343:26]
  assign pipe5_io_pipe_phv_in_is_valid_processor = pipe4_io_pipe_phv_out_is_valid_processor; // @[executor.scala 343:26]
  assign pipe5_io_vliw_in_0 = pipe4_io_vliw_out_0; // @[executor.scala 344:26]
  assign pipe5_io_vliw_in_1 = pipe4_io_vliw_out_1; // @[executor.scala 344:26]
  assign pipe5_io_vliw_in_2 = pipe4_io_vliw_out_2; // @[executor.scala 344:26]
  assign pipe5_io_vliw_in_3 = pipe4_io_vliw_out_3; // @[executor.scala 344:26]
  assign pipe5_io_field_in_0 = pipe4_io_field_out_0; // @[executor.scala 345:26]
  assign pipe5_io_field_in_1 = pipe4_io_field_out_1; // @[executor.scala 345:26]
  assign pipe5_io_field_in_2 = pipe4_io_field_out_2; // @[executor.scala 345:26]
  assign pipe5_io_field_in_3 = pipe4_io_field_out_3; // @[executor.scala 345:26]
  assign pipe6_clock = clock;
  assign pipe6_io_pipe_phv_in_data_0 = pipe5_io_pipe_phv_out_data_0; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_1 = pipe5_io_pipe_phv_out_data_1; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_2 = pipe5_io_pipe_phv_out_data_2; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_3 = pipe5_io_pipe_phv_out_data_3; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_4 = pipe5_io_pipe_phv_out_data_4; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_5 = pipe5_io_pipe_phv_out_data_5; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_6 = pipe5_io_pipe_phv_out_data_6; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_7 = pipe5_io_pipe_phv_out_data_7; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_8 = pipe5_io_pipe_phv_out_data_8; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_9 = pipe5_io_pipe_phv_out_data_9; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_10 = pipe5_io_pipe_phv_out_data_10; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_11 = pipe5_io_pipe_phv_out_data_11; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_12 = pipe5_io_pipe_phv_out_data_12; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_13 = pipe5_io_pipe_phv_out_data_13; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_14 = pipe5_io_pipe_phv_out_data_14; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_15 = pipe5_io_pipe_phv_out_data_15; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_16 = pipe5_io_pipe_phv_out_data_16; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_17 = pipe5_io_pipe_phv_out_data_17; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_18 = pipe5_io_pipe_phv_out_data_18; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_19 = pipe5_io_pipe_phv_out_data_19; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_20 = pipe5_io_pipe_phv_out_data_20; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_21 = pipe5_io_pipe_phv_out_data_21; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_22 = pipe5_io_pipe_phv_out_data_22; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_23 = pipe5_io_pipe_phv_out_data_23; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_24 = pipe5_io_pipe_phv_out_data_24; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_25 = pipe5_io_pipe_phv_out_data_25; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_26 = pipe5_io_pipe_phv_out_data_26; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_27 = pipe5_io_pipe_phv_out_data_27; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_28 = pipe5_io_pipe_phv_out_data_28; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_29 = pipe5_io_pipe_phv_out_data_29; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_30 = pipe5_io_pipe_phv_out_data_30; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_31 = pipe5_io_pipe_phv_out_data_31; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_32 = pipe5_io_pipe_phv_out_data_32; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_33 = pipe5_io_pipe_phv_out_data_33; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_34 = pipe5_io_pipe_phv_out_data_34; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_35 = pipe5_io_pipe_phv_out_data_35; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_36 = pipe5_io_pipe_phv_out_data_36; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_37 = pipe5_io_pipe_phv_out_data_37; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_38 = pipe5_io_pipe_phv_out_data_38; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_39 = pipe5_io_pipe_phv_out_data_39; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_40 = pipe5_io_pipe_phv_out_data_40; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_41 = pipe5_io_pipe_phv_out_data_41; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_42 = pipe5_io_pipe_phv_out_data_42; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_43 = pipe5_io_pipe_phv_out_data_43; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_44 = pipe5_io_pipe_phv_out_data_44; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_45 = pipe5_io_pipe_phv_out_data_45; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_46 = pipe5_io_pipe_phv_out_data_46; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_47 = pipe5_io_pipe_phv_out_data_47; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_48 = pipe5_io_pipe_phv_out_data_48; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_49 = pipe5_io_pipe_phv_out_data_49; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_50 = pipe5_io_pipe_phv_out_data_50; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_51 = pipe5_io_pipe_phv_out_data_51; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_52 = pipe5_io_pipe_phv_out_data_52; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_53 = pipe5_io_pipe_phv_out_data_53; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_54 = pipe5_io_pipe_phv_out_data_54; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_55 = pipe5_io_pipe_phv_out_data_55; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_56 = pipe5_io_pipe_phv_out_data_56; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_57 = pipe5_io_pipe_phv_out_data_57; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_58 = pipe5_io_pipe_phv_out_data_58; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_59 = pipe5_io_pipe_phv_out_data_59; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_60 = pipe5_io_pipe_phv_out_data_60; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_61 = pipe5_io_pipe_phv_out_data_61; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_62 = pipe5_io_pipe_phv_out_data_62; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_63 = pipe5_io_pipe_phv_out_data_63; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_64 = pipe5_io_pipe_phv_out_data_64; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_65 = pipe5_io_pipe_phv_out_data_65; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_66 = pipe5_io_pipe_phv_out_data_66; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_67 = pipe5_io_pipe_phv_out_data_67; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_68 = pipe5_io_pipe_phv_out_data_68; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_69 = pipe5_io_pipe_phv_out_data_69; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_70 = pipe5_io_pipe_phv_out_data_70; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_71 = pipe5_io_pipe_phv_out_data_71; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_72 = pipe5_io_pipe_phv_out_data_72; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_73 = pipe5_io_pipe_phv_out_data_73; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_74 = pipe5_io_pipe_phv_out_data_74; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_75 = pipe5_io_pipe_phv_out_data_75; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_76 = pipe5_io_pipe_phv_out_data_76; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_77 = pipe5_io_pipe_phv_out_data_77; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_78 = pipe5_io_pipe_phv_out_data_78; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_79 = pipe5_io_pipe_phv_out_data_79; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_80 = pipe5_io_pipe_phv_out_data_80; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_81 = pipe5_io_pipe_phv_out_data_81; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_82 = pipe5_io_pipe_phv_out_data_82; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_83 = pipe5_io_pipe_phv_out_data_83; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_84 = pipe5_io_pipe_phv_out_data_84; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_85 = pipe5_io_pipe_phv_out_data_85; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_86 = pipe5_io_pipe_phv_out_data_86; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_87 = pipe5_io_pipe_phv_out_data_87; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_88 = pipe5_io_pipe_phv_out_data_88; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_89 = pipe5_io_pipe_phv_out_data_89; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_90 = pipe5_io_pipe_phv_out_data_90; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_91 = pipe5_io_pipe_phv_out_data_91; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_92 = pipe5_io_pipe_phv_out_data_92; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_93 = pipe5_io_pipe_phv_out_data_93; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_94 = pipe5_io_pipe_phv_out_data_94; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_data_95 = pipe5_io_pipe_phv_out_data_95; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_header_0 = pipe5_io_pipe_phv_out_header_0; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_header_1 = pipe5_io_pipe_phv_out_header_1; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_header_2 = pipe5_io_pipe_phv_out_header_2; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_header_3 = pipe5_io_pipe_phv_out_header_3; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_header_4 = pipe5_io_pipe_phv_out_header_4; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_header_5 = pipe5_io_pipe_phv_out_header_5; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_header_6 = pipe5_io_pipe_phv_out_header_6; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_header_7 = pipe5_io_pipe_phv_out_header_7; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_header_8 = pipe5_io_pipe_phv_out_header_8; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_header_9 = pipe5_io_pipe_phv_out_header_9; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_header_10 = pipe5_io_pipe_phv_out_header_10; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_header_11 = pipe5_io_pipe_phv_out_header_11; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_header_12 = pipe5_io_pipe_phv_out_header_12; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_header_13 = pipe5_io_pipe_phv_out_header_13; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_header_14 = pipe5_io_pipe_phv_out_header_14; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_header_15 = pipe5_io_pipe_phv_out_header_15; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_parse_current_state = pipe5_io_pipe_phv_out_parse_current_state; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_parse_current_offset = pipe5_io_pipe_phv_out_parse_current_offset; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_parse_transition_field = pipe5_io_pipe_phv_out_parse_transition_field; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_next_processor_id = pipe5_io_pipe_phv_out_next_processor_id; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_next_config_id = pipe5_io_pipe_phv_out_next_config_id; // @[executor.scala 347:26]
  assign pipe6_io_pipe_phv_in_is_valid_processor = pipe5_io_pipe_phv_out_is_valid_processor; // @[executor.scala 347:26]
  assign pipe6_io_offset_in_0 = pipe5_io_offset_out_0; // @[executor.scala 349:26]
  assign pipe6_io_offset_in_1 = pipe5_io_offset_out_1; // @[executor.scala 349:26]
  assign pipe6_io_offset_in_2 = pipe5_io_offset_out_2; // @[executor.scala 349:26]
  assign pipe6_io_offset_in_3 = pipe5_io_offset_out_3; // @[executor.scala 349:26]
  assign pipe6_io_length_in_0 = pipe5_io_length_out_0; // @[executor.scala 350:26]
  assign pipe6_io_length_in_1 = pipe5_io_length_out_1; // @[executor.scala 350:26]
  assign pipe6_io_length_in_2 = pipe5_io_length_out_2; // @[executor.scala 350:26]
  assign pipe6_io_length_in_3 = pipe5_io_length_out_3; // @[executor.scala 350:26]
  assign pipe6_io_field_in_0 = pipe5_io_field_out_0; // @[executor.scala 348:26]
  assign pipe6_io_field_in_1 = pipe5_io_field_out_1; // @[executor.scala 348:26]
  assign pipe6_io_field_in_2 = pipe5_io_field_out_2; // @[executor.scala 348:26]
  assign pipe6_io_field_in_3 = pipe5_io_field_out_3; // @[executor.scala 348:26]
endmodule
