module MatchGetOffset(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input  [7:0]  io_key_config_0_header_id,
  input  [7:0]  io_key_config_0_internal_offset,
  input  [7:0]  io_key_config_1_header_id,
  input  [7:0]  io_key_config_1_internal_offset,
  output [7:0]  io_key_offset
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[matcher.scala 34:22]
  reg [7:0] phv_data_1; // @[matcher.scala 34:22]
  reg [7:0] phv_data_2; // @[matcher.scala 34:22]
  reg [7:0] phv_data_3; // @[matcher.scala 34:22]
  reg [7:0] phv_data_4; // @[matcher.scala 34:22]
  reg [7:0] phv_data_5; // @[matcher.scala 34:22]
  reg [7:0] phv_data_6; // @[matcher.scala 34:22]
  reg [7:0] phv_data_7; // @[matcher.scala 34:22]
  reg [7:0] phv_data_8; // @[matcher.scala 34:22]
  reg [7:0] phv_data_9; // @[matcher.scala 34:22]
  reg [7:0] phv_data_10; // @[matcher.scala 34:22]
  reg [7:0] phv_data_11; // @[matcher.scala 34:22]
  reg [7:0] phv_data_12; // @[matcher.scala 34:22]
  reg [7:0] phv_data_13; // @[matcher.scala 34:22]
  reg [7:0] phv_data_14; // @[matcher.scala 34:22]
  reg [7:0] phv_data_15; // @[matcher.scala 34:22]
  reg [7:0] phv_data_16; // @[matcher.scala 34:22]
  reg [7:0] phv_data_17; // @[matcher.scala 34:22]
  reg [7:0] phv_data_18; // @[matcher.scala 34:22]
  reg [7:0] phv_data_19; // @[matcher.scala 34:22]
  reg [7:0] phv_data_20; // @[matcher.scala 34:22]
  reg [7:0] phv_data_21; // @[matcher.scala 34:22]
  reg [7:0] phv_data_22; // @[matcher.scala 34:22]
  reg [7:0] phv_data_23; // @[matcher.scala 34:22]
  reg [7:0] phv_data_24; // @[matcher.scala 34:22]
  reg [7:0] phv_data_25; // @[matcher.scala 34:22]
  reg [7:0] phv_data_26; // @[matcher.scala 34:22]
  reg [7:0] phv_data_27; // @[matcher.scala 34:22]
  reg [7:0] phv_data_28; // @[matcher.scala 34:22]
  reg [7:0] phv_data_29; // @[matcher.scala 34:22]
  reg [7:0] phv_data_30; // @[matcher.scala 34:22]
  reg [7:0] phv_data_31; // @[matcher.scala 34:22]
  reg [7:0] phv_data_32; // @[matcher.scala 34:22]
  reg [7:0] phv_data_33; // @[matcher.scala 34:22]
  reg [7:0] phv_data_34; // @[matcher.scala 34:22]
  reg [7:0] phv_data_35; // @[matcher.scala 34:22]
  reg [7:0] phv_data_36; // @[matcher.scala 34:22]
  reg [7:0] phv_data_37; // @[matcher.scala 34:22]
  reg [7:0] phv_data_38; // @[matcher.scala 34:22]
  reg [7:0] phv_data_39; // @[matcher.scala 34:22]
  reg [7:0] phv_data_40; // @[matcher.scala 34:22]
  reg [7:0] phv_data_41; // @[matcher.scala 34:22]
  reg [7:0] phv_data_42; // @[matcher.scala 34:22]
  reg [7:0] phv_data_43; // @[matcher.scala 34:22]
  reg [7:0] phv_data_44; // @[matcher.scala 34:22]
  reg [7:0] phv_data_45; // @[matcher.scala 34:22]
  reg [7:0] phv_data_46; // @[matcher.scala 34:22]
  reg [7:0] phv_data_47; // @[matcher.scala 34:22]
  reg [7:0] phv_data_48; // @[matcher.scala 34:22]
  reg [7:0] phv_data_49; // @[matcher.scala 34:22]
  reg [7:0] phv_data_50; // @[matcher.scala 34:22]
  reg [7:0] phv_data_51; // @[matcher.scala 34:22]
  reg [7:0] phv_data_52; // @[matcher.scala 34:22]
  reg [7:0] phv_data_53; // @[matcher.scala 34:22]
  reg [7:0] phv_data_54; // @[matcher.scala 34:22]
  reg [7:0] phv_data_55; // @[matcher.scala 34:22]
  reg [7:0] phv_data_56; // @[matcher.scala 34:22]
  reg [7:0] phv_data_57; // @[matcher.scala 34:22]
  reg [7:0] phv_data_58; // @[matcher.scala 34:22]
  reg [7:0] phv_data_59; // @[matcher.scala 34:22]
  reg [7:0] phv_data_60; // @[matcher.scala 34:22]
  reg [7:0] phv_data_61; // @[matcher.scala 34:22]
  reg [7:0] phv_data_62; // @[matcher.scala 34:22]
  reg [7:0] phv_data_63; // @[matcher.scala 34:22]
  reg [7:0] phv_data_64; // @[matcher.scala 34:22]
  reg [7:0] phv_data_65; // @[matcher.scala 34:22]
  reg [7:0] phv_data_66; // @[matcher.scala 34:22]
  reg [7:0] phv_data_67; // @[matcher.scala 34:22]
  reg [7:0] phv_data_68; // @[matcher.scala 34:22]
  reg [7:0] phv_data_69; // @[matcher.scala 34:22]
  reg [7:0] phv_data_70; // @[matcher.scala 34:22]
  reg [7:0] phv_data_71; // @[matcher.scala 34:22]
  reg [7:0] phv_data_72; // @[matcher.scala 34:22]
  reg [7:0] phv_data_73; // @[matcher.scala 34:22]
  reg [7:0] phv_data_74; // @[matcher.scala 34:22]
  reg [7:0] phv_data_75; // @[matcher.scala 34:22]
  reg [7:0] phv_data_76; // @[matcher.scala 34:22]
  reg [7:0] phv_data_77; // @[matcher.scala 34:22]
  reg [7:0] phv_data_78; // @[matcher.scala 34:22]
  reg [7:0] phv_data_79; // @[matcher.scala 34:22]
  reg [7:0] phv_data_80; // @[matcher.scala 34:22]
  reg [7:0] phv_data_81; // @[matcher.scala 34:22]
  reg [7:0] phv_data_82; // @[matcher.scala 34:22]
  reg [7:0] phv_data_83; // @[matcher.scala 34:22]
  reg [7:0] phv_data_84; // @[matcher.scala 34:22]
  reg [7:0] phv_data_85; // @[matcher.scala 34:22]
  reg [7:0] phv_data_86; // @[matcher.scala 34:22]
  reg [7:0] phv_data_87; // @[matcher.scala 34:22]
  reg [7:0] phv_data_88; // @[matcher.scala 34:22]
  reg [7:0] phv_data_89; // @[matcher.scala 34:22]
  reg [7:0] phv_data_90; // @[matcher.scala 34:22]
  reg [7:0] phv_data_91; // @[matcher.scala 34:22]
  reg [7:0] phv_data_92; // @[matcher.scala 34:22]
  reg [7:0] phv_data_93; // @[matcher.scala 34:22]
  reg [7:0] phv_data_94; // @[matcher.scala 34:22]
  reg [7:0] phv_data_95; // @[matcher.scala 34:22]
  reg [15:0] phv_header_0; // @[matcher.scala 34:22]
  reg [15:0] phv_header_1; // @[matcher.scala 34:22]
  reg [15:0] phv_header_2; // @[matcher.scala 34:22]
  reg [15:0] phv_header_3; // @[matcher.scala 34:22]
  reg [15:0] phv_header_4; // @[matcher.scala 34:22]
  reg [15:0] phv_header_5; // @[matcher.scala 34:22]
  reg [15:0] phv_header_6; // @[matcher.scala 34:22]
  reg [15:0] phv_header_7; // @[matcher.scala 34:22]
  reg [15:0] phv_header_8; // @[matcher.scala 34:22]
  reg [15:0] phv_header_9; // @[matcher.scala 34:22]
  reg [15:0] phv_header_10; // @[matcher.scala 34:22]
  reg [15:0] phv_header_11; // @[matcher.scala 34:22]
  reg [15:0] phv_header_12; // @[matcher.scala 34:22]
  reg [15:0] phv_header_13; // @[matcher.scala 34:22]
  reg [15:0] phv_header_14; // @[matcher.scala 34:22]
  reg [15:0] phv_header_15; // @[matcher.scala 34:22]
  reg [7:0] phv_parse_current_state; // @[matcher.scala 34:22]
  reg [7:0] phv_parse_current_offset; // @[matcher.scala 34:22]
  reg [15:0] phv_parse_transition_field; // @[matcher.scala 34:22]
  reg [1:0] phv_next_processor_id; // @[matcher.scala 34:22]
  reg  phv_next_config_id; // @[matcher.scala 34:22]
  reg  phv_is_valid_processor; // @[matcher.scala 34:22]
  wire [7:0] _GEN_4 = phv_next_config_id ? io_key_config_1_header_id : io_key_config_0_header_id; // @[]
  wire [7:0] _GEN_5 = phv_next_config_id ? io_key_config_1_internal_offset : io_key_config_0_internal_offset; // @[]
  wire [15:0] _GEN_9 = 4'h1 == _GEN_4[3:0] ? phv_header_1 : phv_header_0; // @[const.scala 32:43 const.scala 32:43]
  wire [15:0] _GEN_10 = 4'h2 == _GEN_4[3:0] ? phv_header_2 : _GEN_9; // @[const.scala 32:43 const.scala 32:43]
  wire [15:0] _GEN_11 = 4'h3 == _GEN_4[3:0] ? phv_header_3 : _GEN_10; // @[const.scala 32:43 const.scala 32:43]
  wire [15:0] _GEN_12 = 4'h4 == _GEN_4[3:0] ? phv_header_4 : _GEN_11; // @[const.scala 32:43 const.scala 32:43]
  wire [15:0] _GEN_13 = 4'h5 == _GEN_4[3:0] ? phv_header_5 : _GEN_12; // @[const.scala 32:43 const.scala 32:43]
  wire [15:0] _GEN_14 = 4'h6 == _GEN_4[3:0] ? phv_header_6 : _GEN_13; // @[const.scala 32:43 const.scala 32:43]
  wire [15:0] _GEN_15 = 4'h7 == _GEN_4[3:0] ? phv_header_7 : _GEN_14; // @[const.scala 32:43 const.scala 32:43]
  wire [15:0] _GEN_16 = 4'h8 == _GEN_4[3:0] ? phv_header_8 : _GEN_15; // @[const.scala 32:43 const.scala 32:43]
  wire [15:0] _GEN_17 = 4'h9 == _GEN_4[3:0] ? phv_header_9 : _GEN_16; // @[const.scala 32:43 const.scala 32:43]
  wire [15:0] _GEN_18 = 4'ha == _GEN_4[3:0] ? phv_header_10 : _GEN_17; // @[const.scala 32:43 const.scala 32:43]
  wire [15:0] _GEN_19 = 4'hb == _GEN_4[3:0] ? phv_header_11 : _GEN_18; // @[const.scala 32:43 const.scala 32:43]
  wire [15:0] _GEN_20 = 4'hc == _GEN_4[3:0] ? phv_header_12 : _GEN_19; // @[const.scala 32:43 const.scala 32:43]
  wire [15:0] _GEN_21 = 4'hd == _GEN_4[3:0] ? phv_header_13 : _GEN_20; // @[const.scala 32:43 const.scala 32:43]
  wire [15:0] _GEN_22 = 4'he == _GEN_4[3:0] ? phv_header_14 : _GEN_21; // @[const.scala 32:43 const.scala 32:43]
  wire [15:0] _GEN_23 = 4'hf == _GEN_4[3:0] ? phv_header_15 : _GEN_22; // @[const.scala 32:43 const.scala 32:43]
  wire [7:0] header_offset = _GEN_23[15:8]; // @[const.scala 32:43]
  wire [7:0] key_offset = header_offset + _GEN_5; // @[matcher.scala 41:44]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[matcher.scala 36:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[matcher.scala 36:25]
  assign io_key_offset = phv_is_valid_processor ? key_offset : 8'h0; // @[matcher.scala 38:39 matcher.scala 42:27 matcher.scala 44:27]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[matcher.scala 35:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[matcher.scala 35:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[matcher.scala 35:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[matcher.scala 35:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[matcher.scala 35:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[matcher.scala 35:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[matcher.scala 35:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[matcher.scala 35:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[matcher.scala 35:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[matcher.scala 35:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[matcher.scala 35:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[matcher.scala 35:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[matcher.scala 35:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[matcher.scala 35:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[matcher.scala 35:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[matcher.scala 35:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[matcher.scala 35:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[matcher.scala 35:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[matcher.scala 35:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[matcher.scala 35:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[matcher.scala 35:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[matcher.scala 35:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[matcher.scala 35:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[matcher.scala 35:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[matcher.scala 35:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[matcher.scala 35:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[matcher.scala 35:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[matcher.scala 35:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[matcher.scala 35:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[matcher.scala 35:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[matcher.scala 35:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[matcher.scala 35:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[matcher.scala 35:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[matcher.scala 35:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[matcher.scala 35:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[matcher.scala 35:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[matcher.scala 35:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[matcher.scala 35:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[matcher.scala 35:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[matcher.scala 35:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[matcher.scala 35:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[matcher.scala 35:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[matcher.scala 35:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[matcher.scala 35:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[matcher.scala 35:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[matcher.scala 35:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[matcher.scala 35:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[matcher.scala 35:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[matcher.scala 35:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[matcher.scala 35:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[matcher.scala 35:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[matcher.scala 35:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[matcher.scala 35:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[matcher.scala 35:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[matcher.scala 35:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[matcher.scala 35:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[matcher.scala 35:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[matcher.scala 35:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[matcher.scala 35:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[matcher.scala 35:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[matcher.scala 35:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[matcher.scala 35:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[matcher.scala 35:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[matcher.scala 35:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[matcher.scala 35:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[matcher.scala 35:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[matcher.scala 35:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[matcher.scala 35:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[matcher.scala 35:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[matcher.scala 35:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[matcher.scala 35:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[matcher.scala 35:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[matcher.scala 35:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[matcher.scala 35:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[matcher.scala 35:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[matcher.scala 35:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[matcher.scala 35:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[matcher.scala 35:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[matcher.scala 35:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[matcher.scala 35:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[matcher.scala 35:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[matcher.scala 35:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[matcher.scala 35:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[matcher.scala 35:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[matcher.scala 35:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[matcher.scala 35:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[matcher.scala 35:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[matcher.scala 35:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[matcher.scala 35:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[matcher.scala 35:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[matcher.scala 35:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[matcher.scala 35:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[matcher.scala 35:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[matcher.scala 35:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[matcher.scala 35:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[matcher.scala 35:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[matcher.scala 35:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[matcher.scala 35:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[matcher.scala 35:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[matcher.scala 35:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[matcher.scala 35:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[matcher.scala 35:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[matcher.scala 35:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[matcher.scala 35:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[matcher.scala 35:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[matcher.scala 35:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[matcher.scala 35:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[matcher.scala 35:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[matcher.scala 35:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[matcher.scala 35:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[matcher.scala 35:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[matcher.scala 35:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[matcher.scala 35:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[matcher.scala 35:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[matcher.scala 35:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[matcher.scala 35:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[matcher.scala 35:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[matcher.scala 35:13]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  phv_next_config_id = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_117[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MatchGetKey(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input  [3:0]  io_key_config_0_key_length,
  input  [3:0]  io_key_config_1_key_length,
  input  [7:0]  io_key_offset,
  output [63:0] io_match_key
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[matcher.scala 58:22]
  reg [7:0] phv_data_1; // @[matcher.scala 58:22]
  reg [7:0] phv_data_2; // @[matcher.scala 58:22]
  reg [7:0] phv_data_3; // @[matcher.scala 58:22]
  reg [7:0] phv_data_4; // @[matcher.scala 58:22]
  reg [7:0] phv_data_5; // @[matcher.scala 58:22]
  reg [7:0] phv_data_6; // @[matcher.scala 58:22]
  reg [7:0] phv_data_7; // @[matcher.scala 58:22]
  reg [7:0] phv_data_8; // @[matcher.scala 58:22]
  reg [7:0] phv_data_9; // @[matcher.scala 58:22]
  reg [7:0] phv_data_10; // @[matcher.scala 58:22]
  reg [7:0] phv_data_11; // @[matcher.scala 58:22]
  reg [7:0] phv_data_12; // @[matcher.scala 58:22]
  reg [7:0] phv_data_13; // @[matcher.scala 58:22]
  reg [7:0] phv_data_14; // @[matcher.scala 58:22]
  reg [7:0] phv_data_15; // @[matcher.scala 58:22]
  reg [7:0] phv_data_16; // @[matcher.scala 58:22]
  reg [7:0] phv_data_17; // @[matcher.scala 58:22]
  reg [7:0] phv_data_18; // @[matcher.scala 58:22]
  reg [7:0] phv_data_19; // @[matcher.scala 58:22]
  reg [7:0] phv_data_20; // @[matcher.scala 58:22]
  reg [7:0] phv_data_21; // @[matcher.scala 58:22]
  reg [7:0] phv_data_22; // @[matcher.scala 58:22]
  reg [7:0] phv_data_23; // @[matcher.scala 58:22]
  reg [7:0] phv_data_24; // @[matcher.scala 58:22]
  reg [7:0] phv_data_25; // @[matcher.scala 58:22]
  reg [7:0] phv_data_26; // @[matcher.scala 58:22]
  reg [7:0] phv_data_27; // @[matcher.scala 58:22]
  reg [7:0] phv_data_28; // @[matcher.scala 58:22]
  reg [7:0] phv_data_29; // @[matcher.scala 58:22]
  reg [7:0] phv_data_30; // @[matcher.scala 58:22]
  reg [7:0] phv_data_31; // @[matcher.scala 58:22]
  reg [7:0] phv_data_32; // @[matcher.scala 58:22]
  reg [7:0] phv_data_33; // @[matcher.scala 58:22]
  reg [7:0] phv_data_34; // @[matcher.scala 58:22]
  reg [7:0] phv_data_35; // @[matcher.scala 58:22]
  reg [7:0] phv_data_36; // @[matcher.scala 58:22]
  reg [7:0] phv_data_37; // @[matcher.scala 58:22]
  reg [7:0] phv_data_38; // @[matcher.scala 58:22]
  reg [7:0] phv_data_39; // @[matcher.scala 58:22]
  reg [7:0] phv_data_40; // @[matcher.scala 58:22]
  reg [7:0] phv_data_41; // @[matcher.scala 58:22]
  reg [7:0] phv_data_42; // @[matcher.scala 58:22]
  reg [7:0] phv_data_43; // @[matcher.scala 58:22]
  reg [7:0] phv_data_44; // @[matcher.scala 58:22]
  reg [7:0] phv_data_45; // @[matcher.scala 58:22]
  reg [7:0] phv_data_46; // @[matcher.scala 58:22]
  reg [7:0] phv_data_47; // @[matcher.scala 58:22]
  reg [7:0] phv_data_48; // @[matcher.scala 58:22]
  reg [7:0] phv_data_49; // @[matcher.scala 58:22]
  reg [7:0] phv_data_50; // @[matcher.scala 58:22]
  reg [7:0] phv_data_51; // @[matcher.scala 58:22]
  reg [7:0] phv_data_52; // @[matcher.scala 58:22]
  reg [7:0] phv_data_53; // @[matcher.scala 58:22]
  reg [7:0] phv_data_54; // @[matcher.scala 58:22]
  reg [7:0] phv_data_55; // @[matcher.scala 58:22]
  reg [7:0] phv_data_56; // @[matcher.scala 58:22]
  reg [7:0] phv_data_57; // @[matcher.scala 58:22]
  reg [7:0] phv_data_58; // @[matcher.scala 58:22]
  reg [7:0] phv_data_59; // @[matcher.scala 58:22]
  reg [7:0] phv_data_60; // @[matcher.scala 58:22]
  reg [7:0] phv_data_61; // @[matcher.scala 58:22]
  reg [7:0] phv_data_62; // @[matcher.scala 58:22]
  reg [7:0] phv_data_63; // @[matcher.scala 58:22]
  reg [7:0] phv_data_64; // @[matcher.scala 58:22]
  reg [7:0] phv_data_65; // @[matcher.scala 58:22]
  reg [7:0] phv_data_66; // @[matcher.scala 58:22]
  reg [7:0] phv_data_67; // @[matcher.scala 58:22]
  reg [7:0] phv_data_68; // @[matcher.scala 58:22]
  reg [7:0] phv_data_69; // @[matcher.scala 58:22]
  reg [7:0] phv_data_70; // @[matcher.scala 58:22]
  reg [7:0] phv_data_71; // @[matcher.scala 58:22]
  reg [7:0] phv_data_72; // @[matcher.scala 58:22]
  reg [7:0] phv_data_73; // @[matcher.scala 58:22]
  reg [7:0] phv_data_74; // @[matcher.scala 58:22]
  reg [7:0] phv_data_75; // @[matcher.scala 58:22]
  reg [7:0] phv_data_76; // @[matcher.scala 58:22]
  reg [7:0] phv_data_77; // @[matcher.scala 58:22]
  reg [7:0] phv_data_78; // @[matcher.scala 58:22]
  reg [7:0] phv_data_79; // @[matcher.scala 58:22]
  reg [7:0] phv_data_80; // @[matcher.scala 58:22]
  reg [7:0] phv_data_81; // @[matcher.scala 58:22]
  reg [7:0] phv_data_82; // @[matcher.scala 58:22]
  reg [7:0] phv_data_83; // @[matcher.scala 58:22]
  reg [7:0] phv_data_84; // @[matcher.scala 58:22]
  reg [7:0] phv_data_85; // @[matcher.scala 58:22]
  reg [7:0] phv_data_86; // @[matcher.scala 58:22]
  reg [7:0] phv_data_87; // @[matcher.scala 58:22]
  reg [7:0] phv_data_88; // @[matcher.scala 58:22]
  reg [7:0] phv_data_89; // @[matcher.scala 58:22]
  reg [7:0] phv_data_90; // @[matcher.scala 58:22]
  reg [7:0] phv_data_91; // @[matcher.scala 58:22]
  reg [7:0] phv_data_92; // @[matcher.scala 58:22]
  reg [7:0] phv_data_93; // @[matcher.scala 58:22]
  reg [7:0] phv_data_94; // @[matcher.scala 58:22]
  reg [7:0] phv_data_95; // @[matcher.scala 58:22]
  reg [15:0] phv_header_0; // @[matcher.scala 58:22]
  reg [15:0] phv_header_1; // @[matcher.scala 58:22]
  reg [15:0] phv_header_2; // @[matcher.scala 58:22]
  reg [15:0] phv_header_3; // @[matcher.scala 58:22]
  reg [15:0] phv_header_4; // @[matcher.scala 58:22]
  reg [15:0] phv_header_5; // @[matcher.scala 58:22]
  reg [15:0] phv_header_6; // @[matcher.scala 58:22]
  reg [15:0] phv_header_7; // @[matcher.scala 58:22]
  reg [15:0] phv_header_8; // @[matcher.scala 58:22]
  reg [15:0] phv_header_9; // @[matcher.scala 58:22]
  reg [15:0] phv_header_10; // @[matcher.scala 58:22]
  reg [15:0] phv_header_11; // @[matcher.scala 58:22]
  reg [15:0] phv_header_12; // @[matcher.scala 58:22]
  reg [15:0] phv_header_13; // @[matcher.scala 58:22]
  reg [15:0] phv_header_14; // @[matcher.scala 58:22]
  reg [15:0] phv_header_15; // @[matcher.scala 58:22]
  reg [7:0] phv_parse_current_state; // @[matcher.scala 58:22]
  reg [7:0] phv_parse_current_offset; // @[matcher.scala 58:22]
  reg [15:0] phv_parse_transition_field; // @[matcher.scala 58:22]
  reg [1:0] phv_next_processor_id; // @[matcher.scala 58:22]
  reg  phv_next_config_id; // @[matcher.scala 58:22]
  reg  phv_is_valid_processor; // @[matcher.scala 58:22]
  reg [7:0] key_offset; // @[matcher.scala 62:29]
  wire [3:0] _GEN_6 = phv_next_config_id ? io_key_config_1_key_length : io_key_config_0_key_length; // @[matcher.scala 71:36 matcher.scala 71:36]
  wire [8:0] _match_key_bytes_7_T = {{1'd0}, key_offset}; // @[matcher.scala 72:98]
  wire [7:0] _GEN_9 = 7'h1 == _match_key_bytes_7_T[6:0] ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_10 = 7'h2 == _match_key_bytes_7_T[6:0] ? phv_data_2 : _GEN_9; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_11 = 7'h3 == _match_key_bytes_7_T[6:0] ? phv_data_3 : _GEN_10; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_12 = 7'h4 == _match_key_bytes_7_T[6:0] ? phv_data_4 : _GEN_11; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_13 = 7'h5 == _match_key_bytes_7_T[6:0] ? phv_data_5 : _GEN_12; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_14 = 7'h6 == _match_key_bytes_7_T[6:0] ? phv_data_6 : _GEN_13; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_15 = 7'h7 == _match_key_bytes_7_T[6:0] ? phv_data_7 : _GEN_14; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_16 = 7'h8 == _match_key_bytes_7_T[6:0] ? phv_data_8 : _GEN_15; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_17 = 7'h9 == _match_key_bytes_7_T[6:0] ? phv_data_9 : _GEN_16; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_18 = 7'ha == _match_key_bytes_7_T[6:0] ? phv_data_10 : _GEN_17; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_19 = 7'hb == _match_key_bytes_7_T[6:0] ? phv_data_11 : _GEN_18; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_20 = 7'hc == _match_key_bytes_7_T[6:0] ? phv_data_12 : _GEN_19; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_21 = 7'hd == _match_key_bytes_7_T[6:0] ? phv_data_13 : _GEN_20; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_22 = 7'he == _match_key_bytes_7_T[6:0] ? phv_data_14 : _GEN_21; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_23 = 7'hf == _match_key_bytes_7_T[6:0] ? phv_data_15 : _GEN_22; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_24 = 7'h10 == _match_key_bytes_7_T[6:0] ? phv_data_16 : _GEN_23; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_25 = 7'h11 == _match_key_bytes_7_T[6:0] ? phv_data_17 : _GEN_24; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_26 = 7'h12 == _match_key_bytes_7_T[6:0] ? phv_data_18 : _GEN_25; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_27 = 7'h13 == _match_key_bytes_7_T[6:0] ? phv_data_19 : _GEN_26; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_28 = 7'h14 == _match_key_bytes_7_T[6:0] ? phv_data_20 : _GEN_27; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_29 = 7'h15 == _match_key_bytes_7_T[6:0] ? phv_data_21 : _GEN_28; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_30 = 7'h16 == _match_key_bytes_7_T[6:0] ? phv_data_22 : _GEN_29; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_31 = 7'h17 == _match_key_bytes_7_T[6:0] ? phv_data_23 : _GEN_30; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_32 = 7'h18 == _match_key_bytes_7_T[6:0] ? phv_data_24 : _GEN_31; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_33 = 7'h19 == _match_key_bytes_7_T[6:0] ? phv_data_25 : _GEN_32; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_34 = 7'h1a == _match_key_bytes_7_T[6:0] ? phv_data_26 : _GEN_33; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_35 = 7'h1b == _match_key_bytes_7_T[6:0] ? phv_data_27 : _GEN_34; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_36 = 7'h1c == _match_key_bytes_7_T[6:0] ? phv_data_28 : _GEN_35; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_37 = 7'h1d == _match_key_bytes_7_T[6:0] ? phv_data_29 : _GEN_36; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_38 = 7'h1e == _match_key_bytes_7_T[6:0] ? phv_data_30 : _GEN_37; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_39 = 7'h1f == _match_key_bytes_7_T[6:0] ? phv_data_31 : _GEN_38; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_40 = 7'h20 == _match_key_bytes_7_T[6:0] ? phv_data_32 : _GEN_39; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_41 = 7'h21 == _match_key_bytes_7_T[6:0] ? phv_data_33 : _GEN_40; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_42 = 7'h22 == _match_key_bytes_7_T[6:0] ? phv_data_34 : _GEN_41; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_43 = 7'h23 == _match_key_bytes_7_T[6:0] ? phv_data_35 : _GEN_42; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_44 = 7'h24 == _match_key_bytes_7_T[6:0] ? phv_data_36 : _GEN_43; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_45 = 7'h25 == _match_key_bytes_7_T[6:0] ? phv_data_37 : _GEN_44; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_46 = 7'h26 == _match_key_bytes_7_T[6:0] ? phv_data_38 : _GEN_45; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_47 = 7'h27 == _match_key_bytes_7_T[6:0] ? phv_data_39 : _GEN_46; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_48 = 7'h28 == _match_key_bytes_7_T[6:0] ? phv_data_40 : _GEN_47; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_49 = 7'h29 == _match_key_bytes_7_T[6:0] ? phv_data_41 : _GEN_48; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_50 = 7'h2a == _match_key_bytes_7_T[6:0] ? phv_data_42 : _GEN_49; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_51 = 7'h2b == _match_key_bytes_7_T[6:0] ? phv_data_43 : _GEN_50; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_52 = 7'h2c == _match_key_bytes_7_T[6:0] ? phv_data_44 : _GEN_51; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_53 = 7'h2d == _match_key_bytes_7_T[6:0] ? phv_data_45 : _GEN_52; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_54 = 7'h2e == _match_key_bytes_7_T[6:0] ? phv_data_46 : _GEN_53; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_55 = 7'h2f == _match_key_bytes_7_T[6:0] ? phv_data_47 : _GEN_54; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_56 = 7'h30 == _match_key_bytes_7_T[6:0] ? phv_data_48 : _GEN_55; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_57 = 7'h31 == _match_key_bytes_7_T[6:0] ? phv_data_49 : _GEN_56; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_58 = 7'h32 == _match_key_bytes_7_T[6:0] ? phv_data_50 : _GEN_57; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_59 = 7'h33 == _match_key_bytes_7_T[6:0] ? phv_data_51 : _GEN_58; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_60 = 7'h34 == _match_key_bytes_7_T[6:0] ? phv_data_52 : _GEN_59; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_61 = 7'h35 == _match_key_bytes_7_T[6:0] ? phv_data_53 : _GEN_60; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_62 = 7'h36 == _match_key_bytes_7_T[6:0] ? phv_data_54 : _GEN_61; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_63 = 7'h37 == _match_key_bytes_7_T[6:0] ? phv_data_55 : _GEN_62; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_64 = 7'h38 == _match_key_bytes_7_T[6:0] ? phv_data_56 : _GEN_63; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_65 = 7'h39 == _match_key_bytes_7_T[6:0] ? phv_data_57 : _GEN_64; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_66 = 7'h3a == _match_key_bytes_7_T[6:0] ? phv_data_58 : _GEN_65; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_67 = 7'h3b == _match_key_bytes_7_T[6:0] ? phv_data_59 : _GEN_66; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_68 = 7'h3c == _match_key_bytes_7_T[6:0] ? phv_data_60 : _GEN_67; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_69 = 7'h3d == _match_key_bytes_7_T[6:0] ? phv_data_61 : _GEN_68; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_70 = 7'h3e == _match_key_bytes_7_T[6:0] ? phv_data_62 : _GEN_69; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_71 = 7'h3f == _match_key_bytes_7_T[6:0] ? phv_data_63 : _GEN_70; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_72 = 7'h40 == _match_key_bytes_7_T[6:0] ? phv_data_64 : _GEN_71; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_73 = 7'h41 == _match_key_bytes_7_T[6:0] ? phv_data_65 : _GEN_72; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_74 = 7'h42 == _match_key_bytes_7_T[6:0] ? phv_data_66 : _GEN_73; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_75 = 7'h43 == _match_key_bytes_7_T[6:0] ? phv_data_67 : _GEN_74; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_76 = 7'h44 == _match_key_bytes_7_T[6:0] ? phv_data_68 : _GEN_75; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_77 = 7'h45 == _match_key_bytes_7_T[6:0] ? phv_data_69 : _GEN_76; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_78 = 7'h46 == _match_key_bytes_7_T[6:0] ? phv_data_70 : _GEN_77; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_79 = 7'h47 == _match_key_bytes_7_T[6:0] ? phv_data_71 : _GEN_78; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_80 = 7'h48 == _match_key_bytes_7_T[6:0] ? phv_data_72 : _GEN_79; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_81 = 7'h49 == _match_key_bytes_7_T[6:0] ? phv_data_73 : _GEN_80; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_82 = 7'h4a == _match_key_bytes_7_T[6:0] ? phv_data_74 : _GEN_81; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_83 = 7'h4b == _match_key_bytes_7_T[6:0] ? phv_data_75 : _GEN_82; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_84 = 7'h4c == _match_key_bytes_7_T[6:0] ? phv_data_76 : _GEN_83; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_85 = 7'h4d == _match_key_bytes_7_T[6:0] ? phv_data_77 : _GEN_84; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_86 = 7'h4e == _match_key_bytes_7_T[6:0] ? phv_data_78 : _GEN_85; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_87 = 7'h4f == _match_key_bytes_7_T[6:0] ? phv_data_79 : _GEN_86; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_88 = 7'h50 == _match_key_bytes_7_T[6:0] ? phv_data_80 : _GEN_87; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_89 = 7'h51 == _match_key_bytes_7_T[6:0] ? phv_data_81 : _GEN_88; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_90 = 7'h52 == _match_key_bytes_7_T[6:0] ? phv_data_82 : _GEN_89; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_91 = 7'h53 == _match_key_bytes_7_T[6:0] ? phv_data_83 : _GEN_90; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_92 = 7'h54 == _match_key_bytes_7_T[6:0] ? phv_data_84 : _GEN_91; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_93 = 7'h55 == _match_key_bytes_7_T[6:0] ? phv_data_85 : _GEN_92; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_94 = 7'h56 == _match_key_bytes_7_T[6:0] ? phv_data_86 : _GEN_93; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_95 = 7'h57 == _match_key_bytes_7_T[6:0] ? phv_data_87 : _GEN_94; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_96 = 7'h58 == _match_key_bytes_7_T[6:0] ? phv_data_88 : _GEN_95; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_97 = 7'h59 == _match_key_bytes_7_T[6:0] ? phv_data_89 : _GEN_96; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_98 = 7'h5a == _match_key_bytes_7_T[6:0] ? phv_data_90 : _GEN_97; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_99 = 7'h5b == _match_key_bytes_7_T[6:0] ? phv_data_91 : _GEN_98; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_100 = 7'h5c == _match_key_bytes_7_T[6:0] ? phv_data_92 : _GEN_99; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_101 = 7'h5d == _match_key_bytes_7_T[6:0] ? phv_data_93 : _GEN_100; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_102 = 7'h5e == _match_key_bytes_7_T[6:0] ? phv_data_94 : _GEN_101; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_103 = 7'h5f == _match_key_bytes_7_T[6:0] ? phv_data_95 : _GEN_102; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_7 = 4'h0 < _GEN_6 ? _GEN_103 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_6_T_1 = key_offset + 8'h1; // @[matcher.scala 72:98]
  wire [7:0] _GEN_106 = 7'h1 == _match_key_bytes_6_T_1[6:0] ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_107 = 7'h2 == _match_key_bytes_6_T_1[6:0] ? phv_data_2 : _GEN_106; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_108 = 7'h3 == _match_key_bytes_6_T_1[6:0] ? phv_data_3 : _GEN_107; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_109 = 7'h4 == _match_key_bytes_6_T_1[6:0] ? phv_data_4 : _GEN_108; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_110 = 7'h5 == _match_key_bytes_6_T_1[6:0] ? phv_data_5 : _GEN_109; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_111 = 7'h6 == _match_key_bytes_6_T_1[6:0] ? phv_data_6 : _GEN_110; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_112 = 7'h7 == _match_key_bytes_6_T_1[6:0] ? phv_data_7 : _GEN_111; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_113 = 7'h8 == _match_key_bytes_6_T_1[6:0] ? phv_data_8 : _GEN_112; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_114 = 7'h9 == _match_key_bytes_6_T_1[6:0] ? phv_data_9 : _GEN_113; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_115 = 7'ha == _match_key_bytes_6_T_1[6:0] ? phv_data_10 : _GEN_114; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_116 = 7'hb == _match_key_bytes_6_T_1[6:0] ? phv_data_11 : _GEN_115; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_117 = 7'hc == _match_key_bytes_6_T_1[6:0] ? phv_data_12 : _GEN_116; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_118 = 7'hd == _match_key_bytes_6_T_1[6:0] ? phv_data_13 : _GEN_117; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_119 = 7'he == _match_key_bytes_6_T_1[6:0] ? phv_data_14 : _GEN_118; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_120 = 7'hf == _match_key_bytes_6_T_1[6:0] ? phv_data_15 : _GEN_119; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_121 = 7'h10 == _match_key_bytes_6_T_1[6:0] ? phv_data_16 : _GEN_120; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_122 = 7'h11 == _match_key_bytes_6_T_1[6:0] ? phv_data_17 : _GEN_121; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_123 = 7'h12 == _match_key_bytes_6_T_1[6:0] ? phv_data_18 : _GEN_122; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_124 = 7'h13 == _match_key_bytes_6_T_1[6:0] ? phv_data_19 : _GEN_123; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_125 = 7'h14 == _match_key_bytes_6_T_1[6:0] ? phv_data_20 : _GEN_124; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_126 = 7'h15 == _match_key_bytes_6_T_1[6:0] ? phv_data_21 : _GEN_125; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_127 = 7'h16 == _match_key_bytes_6_T_1[6:0] ? phv_data_22 : _GEN_126; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_128 = 7'h17 == _match_key_bytes_6_T_1[6:0] ? phv_data_23 : _GEN_127; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_129 = 7'h18 == _match_key_bytes_6_T_1[6:0] ? phv_data_24 : _GEN_128; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_130 = 7'h19 == _match_key_bytes_6_T_1[6:0] ? phv_data_25 : _GEN_129; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_131 = 7'h1a == _match_key_bytes_6_T_1[6:0] ? phv_data_26 : _GEN_130; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_132 = 7'h1b == _match_key_bytes_6_T_1[6:0] ? phv_data_27 : _GEN_131; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_133 = 7'h1c == _match_key_bytes_6_T_1[6:0] ? phv_data_28 : _GEN_132; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_134 = 7'h1d == _match_key_bytes_6_T_1[6:0] ? phv_data_29 : _GEN_133; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_135 = 7'h1e == _match_key_bytes_6_T_1[6:0] ? phv_data_30 : _GEN_134; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_136 = 7'h1f == _match_key_bytes_6_T_1[6:0] ? phv_data_31 : _GEN_135; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_137 = 7'h20 == _match_key_bytes_6_T_1[6:0] ? phv_data_32 : _GEN_136; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_138 = 7'h21 == _match_key_bytes_6_T_1[6:0] ? phv_data_33 : _GEN_137; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_139 = 7'h22 == _match_key_bytes_6_T_1[6:0] ? phv_data_34 : _GEN_138; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_140 = 7'h23 == _match_key_bytes_6_T_1[6:0] ? phv_data_35 : _GEN_139; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_141 = 7'h24 == _match_key_bytes_6_T_1[6:0] ? phv_data_36 : _GEN_140; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_142 = 7'h25 == _match_key_bytes_6_T_1[6:0] ? phv_data_37 : _GEN_141; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_143 = 7'h26 == _match_key_bytes_6_T_1[6:0] ? phv_data_38 : _GEN_142; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_144 = 7'h27 == _match_key_bytes_6_T_1[6:0] ? phv_data_39 : _GEN_143; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_145 = 7'h28 == _match_key_bytes_6_T_1[6:0] ? phv_data_40 : _GEN_144; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_146 = 7'h29 == _match_key_bytes_6_T_1[6:0] ? phv_data_41 : _GEN_145; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_147 = 7'h2a == _match_key_bytes_6_T_1[6:0] ? phv_data_42 : _GEN_146; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_148 = 7'h2b == _match_key_bytes_6_T_1[6:0] ? phv_data_43 : _GEN_147; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_149 = 7'h2c == _match_key_bytes_6_T_1[6:0] ? phv_data_44 : _GEN_148; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_150 = 7'h2d == _match_key_bytes_6_T_1[6:0] ? phv_data_45 : _GEN_149; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_151 = 7'h2e == _match_key_bytes_6_T_1[6:0] ? phv_data_46 : _GEN_150; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_152 = 7'h2f == _match_key_bytes_6_T_1[6:0] ? phv_data_47 : _GEN_151; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_153 = 7'h30 == _match_key_bytes_6_T_1[6:0] ? phv_data_48 : _GEN_152; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_154 = 7'h31 == _match_key_bytes_6_T_1[6:0] ? phv_data_49 : _GEN_153; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_155 = 7'h32 == _match_key_bytes_6_T_1[6:0] ? phv_data_50 : _GEN_154; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_156 = 7'h33 == _match_key_bytes_6_T_1[6:0] ? phv_data_51 : _GEN_155; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_157 = 7'h34 == _match_key_bytes_6_T_1[6:0] ? phv_data_52 : _GEN_156; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_158 = 7'h35 == _match_key_bytes_6_T_1[6:0] ? phv_data_53 : _GEN_157; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_159 = 7'h36 == _match_key_bytes_6_T_1[6:0] ? phv_data_54 : _GEN_158; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_160 = 7'h37 == _match_key_bytes_6_T_1[6:0] ? phv_data_55 : _GEN_159; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_161 = 7'h38 == _match_key_bytes_6_T_1[6:0] ? phv_data_56 : _GEN_160; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_162 = 7'h39 == _match_key_bytes_6_T_1[6:0] ? phv_data_57 : _GEN_161; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_163 = 7'h3a == _match_key_bytes_6_T_1[6:0] ? phv_data_58 : _GEN_162; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_164 = 7'h3b == _match_key_bytes_6_T_1[6:0] ? phv_data_59 : _GEN_163; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_165 = 7'h3c == _match_key_bytes_6_T_1[6:0] ? phv_data_60 : _GEN_164; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_166 = 7'h3d == _match_key_bytes_6_T_1[6:0] ? phv_data_61 : _GEN_165; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_167 = 7'h3e == _match_key_bytes_6_T_1[6:0] ? phv_data_62 : _GEN_166; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_168 = 7'h3f == _match_key_bytes_6_T_1[6:0] ? phv_data_63 : _GEN_167; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_169 = 7'h40 == _match_key_bytes_6_T_1[6:0] ? phv_data_64 : _GEN_168; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_170 = 7'h41 == _match_key_bytes_6_T_1[6:0] ? phv_data_65 : _GEN_169; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_171 = 7'h42 == _match_key_bytes_6_T_1[6:0] ? phv_data_66 : _GEN_170; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_172 = 7'h43 == _match_key_bytes_6_T_1[6:0] ? phv_data_67 : _GEN_171; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_173 = 7'h44 == _match_key_bytes_6_T_1[6:0] ? phv_data_68 : _GEN_172; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_174 = 7'h45 == _match_key_bytes_6_T_1[6:0] ? phv_data_69 : _GEN_173; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_175 = 7'h46 == _match_key_bytes_6_T_1[6:0] ? phv_data_70 : _GEN_174; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_176 = 7'h47 == _match_key_bytes_6_T_1[6:0] ? phv_data_71 : _GEN_175; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_177 = 7'h48 == _match_key_bytes_6_T_1[6:0] ? phv_data_72 : _GEN_176; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_178 = 7'h49 == _match_key_bytes_6_T_1[6:0] ? phv_data_73 : _GEN_177; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_179 = 7'h4a == _match_key_bytes_6_T_1[6:0] ? phv_data_74 : _GEN_178; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_180 = 7'h4b == _match_key_bytes_6_T_1[6:0] ? phv_data_75 : _GEN_179; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_181 = 7'h4c == _match_key_bytes_6_T_1[6:0] ? phv_data_76 : _GEN_180; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_182 = 7'h4d == _match_key_bytes_6_T_1[6:0] ? phv_data_77 : _GEN_181; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_183 = 7'h4e == _match_key_bytes_6_T_1[6:0] ? phv_data_78 : _GEN_182; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_184 = 7'h4f == _match_key_bytes_6_T_1[6:0] ? phv_data_79 : _GEN_183; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_185 = 7'h50 == _match_key_bytes_6_T_1[6:0] ? phv_data_80 : _GEN_184; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_186 = 7'h51 == _match_key_bytes_6_T_1[6:0] ? phv_data_81 : _GEN_185; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_187 = 7'h52 == _match_key_bytes_6_T_1[6:0] ? phv_data_82 : _GEN_186; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_188 = 7'h53 == _match_key_bytes_6_T_1[6:0] ? phv_data_83 : _GEN_187; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_189 = 7'h54 == _match_key_bytes_6_T_1[6:0] ? phv_data_84 : _GEN_188; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_190 = 7'h55 == _match_key_bytes_6_T_1[6:0] ? phv_data_85 : _GEN_189; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_191 = 7'h56 == _match_key_bytes_6_T_1[6:0] ? phv_data_86 : _GEN_190; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_192 = 7'h57 == _match_key_bytes_6_T_1[6:0] ? phv_data_87 : _GEN_191; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_193 = 7'h58 == _match_key_bytes_6_T_1[6:0] ? phv_data_88 : _GEN_192; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_194 = 7'h59 == _match_key_bytes_6_T_1[6:0] ? phv_data_89 : _GEN_193; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_195 = 7'h5a == _match_key_bytes_6_T_1[6:0] ? phv_data_90 : _GEN_194; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_196 = 7'h5b == _match_key_bytes_6_T_1[6:0] ? phv_data_91 : _GEN_195; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_197 = 7'h5c == _match_key_bytes_6_T_1[6:0] ? phv_data_92 : _GEN_196; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_198 = 7'h5d == _match_key_bytes_6_T_1[6:0] ? phv_data_93 : _GEN_197; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_199 = 7'h5e == _match_key_bytes_6_T_1[6:0] ? phv_data_94 : _GEN_198; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_200 = 7'h5f == _match_key_bytes_6_T_1[6:0] ? phv_data_95 : _GEN_199; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_6 = 4'h1 < _GEN_6 ? _GEN_200 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_5_T_1 = key_offset + 8'h2; // @[matcher.scala 72:98]
  wire [7:0] _GEN_203 = 7'h1 == _match_key_bytes_5_T_1[6:0] ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_204 = 7'h2 == _match_key_bytes_5_T_1[6:0] ? phv_data_2 : _GEN_203; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_205 = 7'h3 == _match_key_bytes_5_T_1[6:0] ? phv_data_3 : _GEN_204; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_206 = 7'h4 == _match_key_bytes_5_T_1[6:0] ? phv_data_4 : _GEN_205; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_207 = 7'h5 == _match_key_bytes_5_T_1[6:0] ? phv_data_5 : _GEN_206; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_208 = 7'h6 == _match_key_bytes_5_T_1[6:0] ? phv_data_6 : _GEN_207; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_209 = 7'h7 == _match_key_bytes_5_T_1[6:0] ? phv_data_7 : _GEN_208; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_210 = 7'h8 == _match_key_bytes_5_T_1[6:0] ? phv_data_8 : _GEN_209; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_211 = 7'h9 == _match_key_bytes_5_T_1[6:0] ? phv_data_9 : _GEN_210; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_212 = 7'ha == _match_key_bytes_5_T_1[6:0] ? phv_data_10 : _GEN_211; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_213 = 7'hb == _match_key_bytes_5_T_1[6:0] ? phv_data_11 : _GEN_212; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_214 = 7'hc == _match_key_bytes_5_T_1[6:0] ? phv_data_12 : _GEN_213; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_215 = 7'hd == _match_key_bytes_5_T_1[6:0] ? phv_data_13 : _GEN_214; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_216 = 7'he == _match_key_bytes_5_T_1[6:0] ? phv_data_14 : _GEN_215; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_217 = 7'hf == _match_key_bytes_5_T_1[6:0] ? phv_data_15 : _GEN_216; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_218 = 7'h10 == _match_key_bytes_5_T_1[6:0] ? phv_data_16 : _GEN_217; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_219 = 7'h11 == _match_key_bytes_5_T_1[6:0] ? phv_data_17 : _GEN_218; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_220 = 7'h12 == _match_key_bytes_5_T_1[6:0] ? phv_data_18 : _GEN_219; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_221 = 7'h13 == _match_key_bytes_5_T_1[6:0] ? phv_data_19 : _GEN_220; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_222 = 7'h14 == _match_key_bytes_5_T_1[6:0] ? phv_data_20 : _GEN_221; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_223 = 7'h15 == _match_key_bytes_5_T_1[6:0] ? phv_data_21 : _GEN_222; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_224 = 7'h16 == _match_key_bytes_5_T_1[6:0] ? phv_data_22 : _GEN_223; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_225 = 7'h17 == _match_key_bytes_5_T_1[6:0] ? phv_data_23 : _GEN_224; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_226 = 7'h18 == _match_key_bytes_5_T_1[6:0] ? phv_data_24 : _GEN_225; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_227 = 7'h19 == _match_key_bytes_5_T_1[6:0] ? phv_data_25 : _GEN_226; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_228 = 7'h1a == _match_key_bytes_5_T_1[6:0] ? phv_data_26 : _GEN_227; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_229 = 7'h1b == _match_key_bytes_5_T_1[6:0] ? phv_data_27 : _GEN_228; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_230 = 7'h1c == _match_key_bytes_5_T_1[6:0] ? phv_data_28 : _GEN_229; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_231 = 7'h1d == _match_key_bytes_5_T_1[6:0] ? phv_data_29 : _GEN_230; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_232 = 7'h1e == _match_key_bytes_5_T_1[6:0] ? phv_data_30 : _GEN_231; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_233 = 7'h1f == _match_key_bytes_5_T_1[6:0] ? phv_data_31 : _GEN_232; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_234 = 7'h20 == _match_key_bytes_5_T_1[6:0] ? phv_data_32 : _GEN_233; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_235 = 7'h21 == _match_key_bytes_5_T_1[6:0] ? phv_data_33 : _GEN_234; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_236 = 7'h22 == _match_key_bytes_5_T_1[6:0] ? phv_data_34 : _GEN_235; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_237 = 7'h23 == _match_key_bytes_5_T_1[6:0] ? phv_data_35 : _GEN_236; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_238 = 7'h24 == _match_key_bytes_5_T_1[6:0] ? phv_data_36 : _GEN_237; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_239 = 7'h25 == _match_key_bytes_5_T_1[6:0] ? phv_data_37 : _GEN_238; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_240 = 7'h26 == _match_key_bytes_5_T_1[6:0] ? phv_data_38 : _GEN_239; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_241 = 7'h27 == _match_key_bytes_5_T_1[6:0] ? phv_data_39 : _GEN_240; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_242 = 7'h28 == _match_key_bytes_5_T_1[6:0] ? phv_data_40 : _GEN_241; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_243 = 7'h29 == _match_key_bytes_5_T_1[6:0] ? phv_data_41 : _GEN_242; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_244 = 7'h2a == _match_key_bytes_5_T_1[6:0] ? phv_data_42 : _GEN_243; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_245 = 7'h2b == _match_key_bytes_5_T_1[6:0] ? phv_data_43 : _GEN_244; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_246 = 7'h2c == _match_key_bytes_5_T_1[6:0] ? phv_data_44 : _GEN_245; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_247 = 7'h2d == _match_key_bytes_5_T_1[6:0] ? phv_data_45 : _GEN_246; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_248 = 7'h2e == _match_key_bytes_5_T_1[6:0] ? phv_data_46 : _GEN_247; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_249 = 7'h2f == _match_key_bytes_5_T_1[6:0] ? phv_data_47 : _GEN_248; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_250 = 7'h30 == _match_key_bytes_5_T_1[6:0] ? phv_data_48 : _GEN_249; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_251 = 7'h31 == _match_key_bytes_5_T_1[6:0] ? phv_data_49 : _GEN_250; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_252 = 7'h32 == _match_key_bytes_5_T_1[6:0] ? phv_data_50 : _GEN_251; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_253 = 7'h33 == _match_key_bytes_5_T_1[6:0] ? phv_data_51 : _GEN_252; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_254 = 7'h34 == _match_key_bytes_5_T_1[6:0] ? phv_data_52 : _GEN_253; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_255 = 7'h35 == _match_key_bytes_5_T_1[6:0] ? phv_data_53 : _GEN_254; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_256 = 7'h36 == _match_key_bytes_5_T_1[6:0] ? phv_data_54 : _GEN_255; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_257 = 7'h37 == _match_key_bytes_5_T_1[6:0] ? phv_data_55 : _GEN_256; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_258 = 7'h38 == _match_key_bytes_5_T_1[6:0] ? phv_data_56 : _GEN_257; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_259 = 7'h39 == _match_key_bytes_5_T_1[6:0] ? phv_data_57 : _GEN_258; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_260 = 7'h3a == _match_key_bytes_5_T_1[6:0] ? phv_data_58 : _GEN_259; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_261 = 7'h3b == _match_key_bytes_5_T_1[6:0] ? phv_data_59 : _GEN_260; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_262 = 7'h3c == _match_key_bytes_5_T_1[6:0] ? phv_data_60 : _GEN_261; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_263 = 7'h3d == _match_key_bytes_5_T_1[6:0] ? phv_data_61 : _GEN_262; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_264 = 7'h3e == _match_key_bytes_5_T_1[6:0] ? phv_data_62 : _GEN_263; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_265 = 7'h3f == _match_key_bytes_5_T_1[6:0] ? phv_data_63 : _GEN_264; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_266 = 7'h40 == _match_key_bytes_5_T_1[6:0] ? phv_data_64 : _GEN_265; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_267 = 7'h41 == _match_key_bytes_5_T_1[6:0] ? phv_data_65 : _GEN_266; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_268 = 7'h42 == _match_key_bytes_5_T_1[6:0] ? phv_data_66 : _GEN_267; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_269 = 7'h43 == _match_key_bytes_5_T_1[6:0] ? phv_data_67 : _GEN_268; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_270 = 7'h44 == _match_key_bytes_5_T_1[6:0] ? phv_data_68 : _GEN_269; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_271 = 7'h45 == _match_key_bytes_5_T_1[6:0] ? phv_data_69 : _GEN_270; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_272 = 7'h46 == _match_key_bytes_5_T_1[6:0] ? phv_data_70 : _GEN_271; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_273 = 7'h47 == _match_key_bytes_5_T_1[6:0] ? phv_data_71 : _GEN_272; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_274 = 7'h48 == _match_key_bytes_5_T_1[6:0] ? phv_data_72 : _GEN_273; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_275 = 7'h49 == _match_key_bytes_5_T_1[6:0] ? phv_data_73 : _GEN_274; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_276 = 7'h4a == _match_key_bytes_5_T_1[6:0] ? phv_data_74 : _GEN_275; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_277 = 7'h4b == _match_key_bytes_5_T_1[6:0] ? phv_data_75 : _GEN_276; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_278 = 7'h4c == _match_key_bytes_5_T_1[6:0] ? phv_data_76 : _GEN_277; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_279 = 7'h4d == _match_key_bytes_5_T_1[6:0] ? phv_data_77 : _GEN_278; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_280 = 7'h4e == _match_key_bytes_5_T_1[6:0] ? phv_data_78 : _GEN_279; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_281 = 7'h4f == _match_key_bytes_5_T_1[6:0] ? phv_data_79 : _GEN_280; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_282 = 7'h50 == _match_key_bytes_5_T_1[6:0] ? phv_data_80 : _GEN_281; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_283 = 7'h51 == _match_key_bytes_5_T_1[6:0] ? phv_data_81 : _GEN_282; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_284 = 7'h52 == _match_key_bytes_5_T_1[6:0] ? phv_data_82 : _GEN_283; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_285 = 7'h53 == _match_key_bytes_5_T_1[6:0] ? phv_data_83 : _GEN_284; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_286 = 7'h54 == _match_key_bytes_5_T_1[6:0] ? phv_data_84 : _GEN_285; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_287 = 7'h55 == _match_key_bytes_5_T_1[6:0] ? phv_data_85 : _GEN_286; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_288 = 7'h56 == _match_key_bytes_5_T_1[6:0] ? phv_data_86 : _GEN_287; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_289 = 7'h57 == _match_key_bytes_5_T_1[6:0] ? phv_data_87 : _GEN_288; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_290 = 7'h58 == _match_key_bytes_5_T_1[6:0] ? phv_data_88 : _GEN_289; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_291 = 7'h59 == _match_key_bytes_5_T_1[6:0] ? phv_data_89 : _GEN_290; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_292 = 7'h5a == _match_key_bytes_5_T_1[6:0] ? phv_data_90 : _GEN_291; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_293 = 7'h5b == _match_key_bytes_5_T_1[6:0] ? phv_data_91 : _GEN_292; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_294 = 7'h5c == _match_key_bytes_5_T_1[6:0] ? phv_data_92 : _GEN_293; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_295 = 7'h5d == _match_key_bytes_5_T_1[6:0] ? phv_data_93 : _GEN_294; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_296 = 7'h5e == _match_key_bytes_5_T_1[6:0] ? phv_data_94 : _GEN_295; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_297 = 7'h5f == _match_key_bytes_5_T_1[6:0] ? phv_data_95 : _GEN_296; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_5 = 4'h2 < _GEN_6 ? _GEN_297 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_4_T_1 = key_offset + 8'h3; // @[matcher.scala 72:98]
  wire [7:0] _GEN_300 = 7'h1 == _match_key_bytes_4_T_1[6:0] ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_301 = 7'h2 == _match_key_bytes_4_T_1[6:0] ? phv_data_2 : _GEN_300; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_302 = 7'h3 == _match_key_bytes_4_T_1[6:0] ? phv_data_3 : _GEN_301; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_303 = 7'h4 == _match_key_bytes_4_T_1[6:0] ? phv_data_4 : _GEN_302; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_304 = 7'h5 == _match_key_bytes_4_T_1[6:0] ? phv_data_5 : _GEN_303; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_305 = 7'h6 == _match_key_bytes_4_T_1[6:0] ? phv_data_6 : _GEN_304; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_306 = 7'h7 == _match_key_bytes_4_T_1[6:0] ? phv_data_7 : _GEN_305; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_307 = 7'h8 == _match_key_bytes_4_T_1[6:0] ? phv_data_8 : _GEN_306; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_308 = 7'h9 == _match_key_bytes_4_T_1[6:0] ? phv_data_9 : _GEN_307; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_309 = 7'ha == _match_key_bytes_4_T_1[6:0] ? phv_data_10 : _GEN_308; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_310 = 7'hb == _match_key_bytes_4_T_1[6:0] ? phv_data_11 : _GEN_309; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_311 = 7'hc == _match_key_bytes_4_T_1[6:0] ? phv_data_12 : _GEN_310; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_312 = 7'hd == _match_key_bytes_4_T_1[6:0] ? phv_data_13 : _GEN_311; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_313 = 7'he == _match_key_bytes_4_T_1[6:0] ? phv_data_14 : _GEN_312; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_314 = 7'hf == _match_key_bytes_4_T_1[6:0] ? phv_data_15 : _GEN_313; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_315 = 7'h10 == _match_key_bytes_4_T_1[6:0] ? phv_data_16 : _GEN_314; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_316 = 7'h11 == _match_key_bytes_4_T_1[6:0] ? phv_data_17 : _GEN_315; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_317 = 7'h12 == _match_key_bytes_4_T_1[6:0] ? phv_data_18 : _GEN_316; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_318 = 7'h13 == _match_key_bytes_4_T_1[6:0] ? phv_data_19 : _GEN_317; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_319 = 7'h14 == _match_key_bytes_4_T_1[6:0] ? phv_data_20 : _GEN_318; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_320 = 7'h15 == _match_key_bytes_4_T_1[6:0] ? phv_data_21 : _GEN_319; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_321 = 7'h16 == _match_key_bytes_4_T_1[6:0] ? phv_data_22 : _GEN_320; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_322 = 7'h17 == _match_key_bytes_4_T_1[6:0] ? phv_data_23 : _GEN_321; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_323 = 7'h18 == _match_key_bytes_4_T_1[6:0] ? phv_data_24 : _GEN_322; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_324 = 7'h19 == _match_key_bytes_4_T_1[6:0] ? phv_data_25 : _GEN_323; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_325 = 7'h1a == _match_key_bytes_4_T_1[6:0] ? phv_data_26 : _GEN_324; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_326 = 7'h1b == _match_key_bytes_4_T_1[6:0] ? phv_data_27 : _GEN_325; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_327 = 7'h1c == _match_key_bytes_4_T_1[6:0] ? phv_data_28 : _GEN_326; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_328 = 7'h1d == _match_key_bytes_4_T_1[6:0] ? phv_data_29 : _GEN_327; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_329 = 7'h1e == _match_key_bytes_4_T_1[6:0] ? phv_data_30 : _GEN_328; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_330 = 7'h1f == _match_key_bytes_4_T_1[6:0] ? phv_data_31 : _GEN_329; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_331 = 7'h20 == _match_key_bytes_4_T_1[6:0] ? phv_data_32 : _GEN_330; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_332 = 7'h21 == _match_key_bytes_4_T_1[6:0] ? phv_data_33 : _GEN_331; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_333 = 7'h22 == _match_key_bytes_4_T_1[6:0] ? phv_data_34 : _GEN_332; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_334 = 7'h23 == _match_key_bytes_4_T_1[6:0] ? phv_data_35 : _GEN_333; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_335 = 7'h24 == _match_key_bytes_4_T_1[6:0] ? phv_data_36 : _GEN_334; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_336 = 7'h25 == _match_key_bytes_4_T_1[6:0] ? phv_data_37 : _GEN_335; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_337 = 7'h26 == _match_key_bytes_4_T_1[6:0] ? phv_data_38 : _GEN_336; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_338 = 7'h27 == _match_key_bytes_4_T_1[6:0] ? phv_data_39 : _GEN_337; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_339 = 7'h28 == _match_key_bytes_4_T_1[6:0] ? phv_data_40 : _GEN_338; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_340 = 7'h29 == _match_key_bytes_4_T_1[6:0] ? phv_data_41 : _GEN_339; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_341 = 7'h2a == _match_key_bytes_4_T_1[6:0] ? phv_data_42 : _GEN_340; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_342 = 7'h2b == _match_key_bytes_4_T_1[6:0] ? phv_data_43 : _GEN_341; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_343 = 7'h2c == _match_key_bytes_4_T_1[6:0] ? phv_data_44 : _GEN_342; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_344 = 7'h2d == _match_key_bytes_4_T_1[6:0] ? phv_data_45 : _GEN_343; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_345 = 7'h2e == _match_key_bytes_4_T_1[6:0] ? phv_data_46 : _GEN_344; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_346 = 7'h2f == _match_key_bytes_4_T_1[6:0] ? phv_data_47 : _GEN_345; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_347 = 7'h30 == _match_key_bytes_4_T_1[6:0] ? phv_data_48 : _GEN_346; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_348 = 7'h31 == _match_key_bytes_4_T_1[6:0] ? phv_data_49 : _GEN_347; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_349 = 7'h32 == _match_key_bytes_4_T_1[6:0] ? phv_data_50 : _GEN_348; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_350 = 7'h33 == _match_key_bytes_4_T_1[6:0] ? phv_data_51 : _GEN_349; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_351 = 7'h34 == _match_key_bytes_4_T_1[6:0] ? phv_data_52 : _GEN_350; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_352 = 7'h35 == _match_key_bytes_4_T_1[6:0] ? phv_data_53 : _GEN_351; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_353 = 7'h36 == _match_key_bytes_4_T_1[6:0] ? phv_data_54 : _GEN_352; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_354 = 7'h37 == _match_key_bytes_4_T_1[6:0] ? phv_data_55 : _GEN_353; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_355 = 7'h38 == _match_key_bytes_4_T_1[6:0] ? phv_data_56 : _GEN_354; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_356 = 7'h39 == _match_key_bytes_4_T_1[6:0] ? phv_data_57 : _GEN_355; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_357 = 7'h3a == _match_key_bytes_4_T_1[6:0] ? phv_data_58 : _GEN_356; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_358 = 7'h3b == _match_key_bytes_4_T_1[6:0] ? phv_data_59 : _GEN_357; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_359 = 7'h3c == _match_key_bytes_4_T_1[6:0] ? phv_data_60 : _GEN_358; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_360 = 7'h3d == _match_key_bytes_4_T_1[6:0] ? phv_data_61 : _GEN_359; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_361 = 7'h3e == _match_key_bytes_4_T_1[6:0] ? phv_data_62 : _GEN_360; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_362 = 7'h3f == _match_key_bytes_4_T_1[6:0] ? phv_data_63 : _GEN_361; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_363 = 7'h40 == _match_key_bytes_4_T_1[6:0] ? phv_data_64 : _GEN_362; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_364 = 7'h41 == _match_key_bytes_4_T_1[6:0] ? phv_data_65 : _GEN_363; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_365 = 7'h42 == _match_key_bytes_4_T_1[6:0] ? phv_data_66 : _GEN_364; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_366 = 7'h43 == _match_key_bytes_4_T_1[6:0] ? phv_data_67 : _GEN_365; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_367 = 7'h44 == _match_key_bytes_4_T_1[6:0] ? phv_data_68 : _GEN_366; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_368 = 7'h45 == _match_key_bytes_4_T_1[6:0] ? phv_data_69 : _GEN_367; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_369 = 7'h46 == _match_key_bytes_4_T_1[6:0] ? phv_data_70 : _GEN_368; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_370 = 7'h47 == _match_key_bytes_4_T_1[6:0] ? phv_data_71 : _GEN_369; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_371 = 7'h48 == _match_key_bytes_4_T_1[6:0] ? phv_data_72 : _GEN_370; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_372 = 7'h49 == _match_key_bytes_4_T_1[6:0] ? phv_data_73 : _GEN_371; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_373 = 7'h4a == _match_key_bytes_4_T_1[6:0] ? phv_data_74 : _GEN_372; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_374 = 7'h4b == _match_key_bytes_4_T_1[6:0] ? phv_data_75 : _GEN_373; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_375 = 7'h4c == _match_key_bytes_4_T_1[6:0] ? phv_data_76 : _GEN_374; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_376 = 7'h4d == _match_key_bytes_4_T_1[6:0] ? phv_data_77 : _GEN_375; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_377 = 7'h4e == _match_key_bytes_4_T_1[6:0] ? phv_data_78 : _GEN_376; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_378 = 7'h4f == _match_key_bytes_4_T_1[6:0] ? phv_data_79 : _GEN_377; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_379 = 7'h50 == _match_key_bytes_4_T_1[6:0] ? phv_data_80 : _GEN_378; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_380 = 7'h51 == _match_key_bytes_4_T_1[6:0] ? phv_data_81 : _GEN_379; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_381 = 7'h52 == _match_key_bytes_4_T_1[6:0] ? phv_data_82 : _GEN_380; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_382 = 7'h53 == _match_key_bytes_4_T_1[6:0] ? phv_data_83 : _GEN_381; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_383 = 7'h54 == _match_key_bytes_4_T_1[6:0] ? phv_data_84 : _GEN_382; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_384 = 7'h55 == _match_key_bytes_4_T_1[6:0] ? phv_data_85 : _GEN_383; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_385 = 7'h56 == _match_key_bytes_4_T_1[6:0] ? phv_data_86 : _GEN_384; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_386 = 7'h57 == _match_key_bytes_4_T_1[6:0] ? phv_data_87 : _GEN_385; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_387 = 7'h58 == _match_key_bytes_4_T_1[6:0] ? phv_data_88 : _GEN_386; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_388 = 7'h59 == _match_key_bytes_4_T_1[6:0] ? phv_data_89 : _GEN_387; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_389 = 7'h5a == _match_key_bytes_4_T_1[6:0] ? phv_data_90 : _GEN_388; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_390 = 7'h5b == _match_key_bytes_4_T_1[6:0] ? phv_data_91 : _GEN_389; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_391 = 7'h5c == _match_key_bytes_4_T_1[6:0] ? phv_data_92 : _GEN_390; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_392 = 7'h5d == _match_key_bytes_4_T_1[6:0] ? phv_data_93 : _GEN_391; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_393 = 7'h5e == _match_key_bytes_4_T_1[6:0] ? phv_data_94 : _GEN_392; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_394 = 7'h5f == _match_key_bytes_4_T_1[6:0] ? phv_data_95 : _GEN_393; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_4 = 4'h3 < _GEN_6 ? _GEN_394 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_3_T_1 = key_offset + 8'h4; // @[matcher.scala 72:98]
  wire [7:0] _GEN_397 = 7'h1 == _match_key_bytes_3_T_1[6:0] ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_398 = 7'h2 == _match_key_bytes_3_T_1[6:0] ? phv_data_2 : _GEN_397; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_399 = 7'h3 == _match_key_bytes_3_T_1[6:0] ? phv_data_3 : _GEN_398; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_400 = 7'h4 == _match_key_bytes_3_T_1[6:0] ? phv_data_4 : _GEN_399; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_401 = 7'h5 == _match_key_bytes_3_T_1[6:0] ? phv_data_5 : _GEN_400; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_402 = 7'h6 == _match_key_bytes_3_T_1[6:0] ? phv_data_6 : _GEN_401; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_403 = 7'h7 == _match_key_bytes_3_T_1[6:0] ? phv_data_7 : _GEN_402; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_404 = 7'h8 == _match_key_bytes_3_T_1[6:0] ? phv_data_8 : _GEN_403; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_405 = 7'h9 == _match_key_bytes_3_T_1[6:0] ? phv_data_9 : _GEN_404; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_406 = 7'ha == _match_key_bytes_3_T_1[6:0] ? phv_data_10 : _GEN_405; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_407 = 7'hb == _match_key_bytes_3_T_1[6:0] ? phv_data_11 : _GEN_406; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_408 = 7'hc == _match_key_bytes_3_T_1[6:0] ? phv_data_12 : _GEN_407; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_409 = 7'hd == _match_key_bytes_3_T_1[6:0] ? phv_data_13 : _GEN_408; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_410 = 7'he == _match_key_bytes_3_T_1[6:0] ? phv_data_14 : _GEN_409; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_411 = 7'hf == _match_key_bytes_3_T_1[6:0] ? phv_data_15 : _GEN_410; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_412 = 7'h10 == _match_key_bytes_3_T_1[6:0] ? phv_data_16 : _GEN_411; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_413 = 7'h11 == _match_key_bytes_3_T_1[6:0] ? phv_data_17 : _GEN_412; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_414 = 7'h12 == _match_key_bytes_3_T_1[6:0] ? phv_data_18 : _GEN_413; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_415 = 7'h13 == _match_key_bytes_3_T_1[6:0] ? phv_data_19 : _GEN_414; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_416 = 7'h14 == _match_key_bytes_3_T_1[6:0] ? phv_data_20 : _GEN_415; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_417 = 7'h15 == _match_key_bytes_3_T_1[6:0] ? phv_data_21 : _GEN_416; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_418 = 7'h16 == _match_key_bytes_3_T_1[6:0] ? phv_data_22 : _GEN_417; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_419 = 7'h17 == _match_key_bytes_3_T_1[6:0] ? phv_data_23 : _GEN_418; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_420 = 7'h18 == _match_key_bytes_3_T_1[6:0] ? phv_data_24 : _GEN_419; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_421 = 7'h19 == _match_key_bytes_3_T_1[6:0] ? phv_data_25 : _GEN_420; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_422 = 7'h1a == _match_key_bytes_3_T_1[6:0] ? phv_data_26 : _GEN_421; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_423 = 7'h1b == _match_key_bytes_3_T_1[6:0] ? phv_data_27 : _GEN_422; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_424 = 7'h1c == _match_key_bytes_3_T_1[6:0] ? phv_data_28 : _GEN_423; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_425 = 7'h1d == _match_key_bytes_3_T_1[6:0] ? phv_data_29 : _GEN_424; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_426 = 7'h1e == _match_key_bytes_3_T_1[6:0] ? phv_data_30 : _GEN_425; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_427 = 7'h1f == _match_key_bytes_3_T_1[6:0] ? phv_data_31 : _GEN_426; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_428 = 7'h20 == _match_key_bytes_3_T_1[6:0] ? phv_data_32 : _GEN_427; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_429 = 7'h21 == _match_key_bytes_3_T_1[6:0] ? phv_data_33 : _GEN_428; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_430 = 7'h22 == _match_key_bytes_3_T_1[6:0] ? phv_data_34 : _GEN_429; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_431 = 7'h23 == _match_key_bytes_3_T_1[6:0] ? phv_data_35 : _GEN_430; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_432 = 7'h24 == _match_key_bytes_3_T_1[6:0] ? phv_data_36 : _GEN_431; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_433 = 7'h25 == _match_key_bytes_3_T_1[6:0] ? phv_data_37 : _GEN_432; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_434 = 7'h26 == _match_key_bytes_3_T_1[6:0] ? phv_data_38 : _GEN_433; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_435 = 7'h27 == _match_key_bytes_3_T_1[6:0] ? phv_data_39 : _GEN_434; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_436 = 7'h28 == _match_key_bytes_3_T_1[6:0] ? phv_data_40 : _GEN_435; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_437 = 7'h29 == _match_key_bytes_3_T_1[6:0] ? phv_data_41 : _GEN_436; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_438 = 7'h2a == _match_key_bytes_3_T_1[6:0] ? phv_data_42 : _GEN_437; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_439 = 7'h2b == _match_key_bytes_3_T_1[6:0] ? phv_data_43 : _GEN_438; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_440 = 7'h2c == _match_key_bytes_3_T_1[6:0] ? phv_data_44 : _GEN_439; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_441 = 7'h2d == _match_key_bytes_3_T_1[6:0] ? phv_data_45 : _GEN_440; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_442 = 7'h2e == _match_key_bytes_3_T_1[6:0] ? phv_data_46 : _GEN_441; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_443 = 7'h2f == _match_key_bytes_3_T_1[6:0] ? phv_data_47 : _GEN_442; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_444 = 7'h30 == _match_key_bytes_3_T_1[6:0] ? phv_data_48 : _GEN_443; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_445 = 7'h31 == _match_key_bytes_3_T_1[6:0] ? phv_data_49 : _GEN_444; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_446 = 7'h32 == _match_key_bytes_3_T_1[6:0] ? phv_data_50 : _GEN_445; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_447 = 7'h33 == _match_key_bytes_3_T_1[6:0] ? phv_data_51 : _GEN_446; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_448 = 7'h34 == _match_key_bytes_3_T_1[6:0] ? phv_data_52 : _GEN_447; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_449 = 7'h35 == _match_key_bytes_3_T_1[6:0] ? phv_data_53 : _GEN_448; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_450 = 7'h36 == _match_key_bytes_3_T_1[6:0] ? phv_data_54 : _GEN_449; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_451 = 7'h37 == _match_key_bytes_3_T_1[6:0] ? phv_data_55 : _GEN_450; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_452 = 7'h38 == _match_key_bytes_3_T_1[6:0] ? phv_data_56 : _GEN_451; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_453 = 7'h39 == _match_key_bytes_3_T_1[6:0] ? phv_data_57 : _GEN_452; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_454 = 7'h3a == _match_key_bytes_3_T_1[6:0] ? phv_data_58 : _GEN_453; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_455 = 7'h3b == _match_key_bytes_3_T_1[6:0] ? phv_data_59 : _GEN_454; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_456 = 7'h3c == _match_key_bytes_3_T_1[6:0] ? phv_data_60 : _GEN_455; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_457 = 7'h3d == _match_key_bytes_3_T_1[6:0] ? phv_data_61 : _GEN_456; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_458 = 7'h3e == _match_key_bytes_3_T_1[6:0] ? phv_data_62 : _GEN_457; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_459 = 7'h3f == _match_key_bytes_3_T_1[6:0] ? phv_data_63 : _GEN_458; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_460 = 7'h40 == _match_key_bytes_3_T_1[6:0] ? phv_data_64 : _GEN_459; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_461 = 7'h41 == _match_key_bytes_3_T_1[6:0] ? phv_data_65 : _GEN_460; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_462 = 7'h42 == _match_key_bytes_3_T_1[6:0] ? phv_data_66 : _GEN_461; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_463 = 7'h43 == _match_key_bytes_3_T_1[6:0] ? phv_data_67 : _GEN_462; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_464 = 7'h44 == _match_key_bytes_3_T_1[6:0] ? phv_data_68 : _GEN_463; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_465 = 7'h45 == _match_key_bytes_3_T_1[6:0] ? phv_data_69 : _GEN_464; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_466 = 7'h46 == _match_key_bytes_3_T_1[6:0] ? phv_data_70 : _GEN_465; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_467 = 7'h47 == _match_key_bytes_3_T_1[6:0] ? phv_data_71 : _GEN_466; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_468 = 7'h48 == _match_key_bytes_3_T_1[6:0] ? phv_data_72 : _GEN_467; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_469 = 7'h49 == _match_key_bytes_3_T_1[6:0] ? phv_data_73 : _GEN_468; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_470 = 7'h4a == _match_key_bytes_3_T_1[6:0] ? phv_data_74 : _GEN_469; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_471 = 7'h4b == _match_key_bytes_3_T_1[6:0] ? phv_data_75 : _GEN_470; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_472 = 7'h4c == _match_key_bytes_3_T_1[6:0] ? phv_data_76 : _GEN_471; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_473 = 7'h4d == _match_key_bytes_3_T_1[6:0] ? phv_data_77 : _GEN_472; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_474 = 7'h4e == _match_key_bytes_3_T_1[6:0] ? phv_data_78 : _GEN_473; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_475 = 7'h4f == _match_key_bytes_3_T_1[6:0] ? phv_data_79 : _GEN_474; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_476 = 7'h50 == _match_key_bytes_3_T_1[6:0] ? phv_data_80 : _GEN_475; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_477 = 7'h51 == _match_key_bytes_3_T_1[6:0] ? phv_data_81 : _GEN_476; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_478 = 7'h52 == _match_key_bytes_3_T_1[6:0] ? phv_data_82 : _GEN_477; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_479 = 7'h53 == _match_key_bytes_3_T_1[6:0] ? phv_data_83 : _GEN_478; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_480 = 7'h54 == _match_key_bytes_3_T_1[6:0] ? phv_data_84 : _GEN_479; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_481 = 7'h55 == _match_key_bytes_3_T_1[6:0] ? phv_data_85 : _GEN_480; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_482 = 7'h56 == _match_key_bytes_3_T_1[6:0] ? phv_data_86 : _GEN_481; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_483 = 7'h57 == _match_key_bytes_3_T_1[6:0] ? phv_data_87 : _GEN_482; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_484 = 7'h58 == _match_key_bytes_3_T_1[6:0] ? phv_data_88 : _GEN_483; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_485 = 7'h59 == _match_key_bytes_3_T_1[6:0] ? phv_data_89 : _GEN_484; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_486 = 7'h5a == _match_key_bytes_3_T_1[6:0] ? phv_data_90 : _GEN_485; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_487 = 7'h5b == _match_key_bytes_3_T_1[6:0] ? phv_data_91 : _GEN_486; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_488 = 7'h5c == _match_key_bytes_3_T_1[6:0] ? phv_data_92 : _GEN_487; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_489 = 7'h5d == _match_key_bytes_3_T_1[6:0] ? phv_data_93 : _GEN_488; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_490 = 7'h5e == _match_key_bytes_3_T_1[6:0] ? phv_data_94 : _GEN_489; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_491 = 7'h5f == _match_key_bytes_3_T_1[6:0] ? phv_data_95 : _GEN_490; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_3 = 4'h4 < _GEN_6 ? _GEN_491 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_2_T_1 = key_offset + 8'h5; // @[matcher.scala 72:98]
  wire [7:0] _GEN_494 = 7'h1 == _match_key_bytes_2_T_1[6:0] ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_495 = 7'h2 == _match_key_bytes_2_T_1[6:0] ? phv_data_2 : _GEN_494; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_496 = 7'h3 == _match_key_bytes_2_T_1[6:0] ? phv_data_3 : _GEN_495; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_497 = 7'h4 == _match_key_bytes_2_T_1[6:0] ? phv_data_4 : _GEN_496; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_498 = 7'h5 == _match_key_bytes_2_T_1[6:0] ? phv_data_5 : _GEN_497; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_499 = 7'h6 == _match_key_bytes_2_T_1[6:0] ? phv_data_6 : _GEN_498; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_500 = 7'h7 == _match_key_bytes_2_T_1[6:0] ? phv_data_7 : _GEN_499; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_501 = 7'h8 == _match_key_bytes_2_T_1[6:0] ? phv_data_8 : _GEN_500; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_502 = 7'h9 == _match_key_bytes_2_T_1[6:0] ? phv_data_9 : _GEN_501; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_503 = 7'ha == _match_key_bytes_2_T_1[6:0] ? phv_data_10 : _GEN_502; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_504 = 7'hb == _match_key_bytes_2_T_1[6:0] ? phv_data_11 : _GEN_503; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_505 = 7'hc == _match_key_bytes_2_T_1[6:0] ? phv_data_12 : _GEN_504; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_506 = 7'hd == _match_key_bytes_2_T_1[6:0] ? phv_data_13 : _GEN_505; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_507 = 7'he == _match_key_bytes_2_T_1[6:0] ? phv_data_14 : _GEN_506; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_508 = 7'hf == _match_key_bytes_2_T_1[6:0] ? phv_data_15 : _GEN_507; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_509 = 7'h10 == _match_key_bytes_2_T_1[6:0] ? phv_data_16 : _GEN_508; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_510 = 7'h11 == _match_key_bytes_2_T_1[6:0] ? phv_data_17 : _GEN_509; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_511 = 7'h12 == _match_key_bytes_2_T_1[6:0] ? phv_data_18 : _GEN_510; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_512 = 7'h13 == _match_key_bytes_2_T_1[6:0] ? phv_data_19 : _GEN_511; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_513 = 7'h14 == _match_key_bytes_2_T_1[6:0] ? phv_data_20 : _GEN_512; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_514 = 7'h15 == _match_key_bytes_2_T_1[6:0] ? phv_data_21 : _GEN_513; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_515 = 7'h16 == _match_key_bytes_2_T_1[6:0] ? phv_data_22 : _GEN_514; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_516 = 7'h17 == _match_key_bytes_2_T_1[6:0] ? phv_data_23 : _GEN_515; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_517 = 7'h18 == _match_key_bytes_2_T_1[6:0] ? phv_data_24 : _GEN_516; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_518 = 7'h19 == _match_key_bytes_2_T_1[6:0] ? phv_data_25 : _GEN_517; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_519 = 7'h1a == _match_key_bytes_2_T_1[6:0] ? phv_data_26 : _GEN_518; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_520 = 7'h1b == _match_key_bytes_2_T_1[6:0] ? phv_data_27 : _GEN_519; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_521 = 7'h1c == _match_key_bytes_2_T_1[6:0] ? phv_data_28 : _GEN_520; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_522 = 7'h1d == _match_key_bytes_2_T_1[6:0] ? phv_data_29 : _GEN_521; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_523 = 7'h1e == _match_key_bytes_2_T_1[6:0] ? phv_data_30 : _GEN_522; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_524 = 7'h1f == _match_key_bytes_2_T_1[6:0] ? phv_data_31 : _GEN_523; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_525 = 7'h20 == _match_key_bytes_2_T_1[6:0] ? phv_data_32 : _GEN_524; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_526 = 7'h21 == _match_key_bytes_2_T_1[6:0] ? phv_data_33 : _GEN_525; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_527 = 7'h22 == _match_key_bytes_2_T_1[6:0] ? phv_data_34 : _GEN_526; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_528 = 7'h23 == _match_key_bytes_2_T_1[6:0] ? phv_data_35 : _GEN_527; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_529 = 7'h24 == _match_key_bytes_2_T_1[6:0] ? phv_data_36 : _GEN_528; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_530 = 7'h25 == _match_key_bytes_2_T_1[6:0] ? phv_data_37 : _GEN_529; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_531 = 7'h26 == _match_key_bytes_2_T_1[6:0] ? phv_data_38 : _GEN_530; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_532 = 7'h27 == _match_key_bytes_2_T_1[6:0] ? phv_data_39 : _GEN_531; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_533 = 7'h28 == _match_key_bytes_2_T_1[6:0] ? phv_data_40 : _GEN_532; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_534 = 7'h29 == _match_key_bytes_2_T_1[6:0] ? phv_data_41 : _GEN_533; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_535 = 7'h2a == _match_key_bytes_2_T_1[6:0] ? phv_data_42 : _GEN_534; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_536 = 7'h2b == _match_key_bytes_2_T_1[6:0] ? phv_data_43 : _GEN_535; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_537 = 7'h2c == _match_key_bytes_2_T_1[6:0] ? phv_data_44 : _GEN_536; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_538 = 7'h2d == _match_key_bytes_2_T_1[6:0] ? phv_data_45 : _GEN_537; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_539 = 7'h2e == _match_key_bytes_2_T_1[6:0] ? phv_data_46 : _GEN_538; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_540 = 7'h2f == _match_key_bytes_2_T_1[6:0] ? phv_data_47 : _GEN_539; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_541 = 7'h30 == _match_key_bytes_2_T_1[6:0] ? phv_data_48 : _GEN_540; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_542 = 7'h31 == _match_key_bytes_2_T_1[6:0] ? phv_data_49 : _GEN_541; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_543 = 7'h32 == _match_key_bytes_2_T_1[6:0] ? phv_data_50 : _GEN_542; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_544 = 7'h33 == _match_key_bytes_2_T_1[6:0] ? phv_data_51 : _GEN_543; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_545 = 7'h34 == _match_key_bytes_2_T_1[6:0] ? phv_data_52 : _GEN_544; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_546 = 7'h35 == _match_key_bytes_2_T_1[6:0] ? phv_data_53 : _GEN_545; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_547 = 7'h36 == _match_key_bytes_2_T_1[6:0] ? phv_data_54 : _GEN_546; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_548 = 7'h37 == _match_key_bytes_2_T_1[6:0] ? phv_data_55 : _GEN_547; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_549 = 7'h38 == _match_key_bytes_2_T_1[6:0] ? phv_data_56 : _GEN_548; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_550 = 7'h39 == _match_key_bytes_2_T_1[6:0] ? phv_data_57 : _GEN_549; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_551 = 7'h3a == _match_key_bytes_2_T_1[6:0] ? phv_data_58 : _GEN_550; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_552 = 7'h3b == _match_key_bytes_2_T_1[6:0] ? phv_data_59 : _GEN_551; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_553 = 7'h3c == _match_key_bytes_2_T_1[6:0] ? phv_data_60 : _GEN_552; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_554 = 7'h3d == _match_key_bytes_2_T_1[6:0] ? phv_data_61 : _GEN_553; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_555 = 7'h3e == _match_key_bytes_2_T_1[6:0] ? phv_data_62 : _GEN_554; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_556 = 7'h3f == _match_key_bytes_2_T_1[6:0] ? phv_data_63 : _GEN_555; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_557 = 7'h40 == _match_key_bytes_2_T_1[6:0] ? phv_data_64 : _GEN_556; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_558 = 7'h41 == _match_key_bytes_2_T_1[6:0] ? phv_data_65 : _GEN_557; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_559 = 7'h42 == _match_key_bytes_2_T_1[6:0] ? phv_data_66 : _GEN_558; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_560 = 7'h43 == _match_key_bytes_2_T_1[6:0] ? phv_data_67 : _GEN_559; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_561 = 7'h44 == _match_key_bytes_2_T_1[6:0] ? phv_data_68 : _GEN_560; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_562 = 7'h45 == _match_key_bytes_2_T_1[6:0] ? phv_data_69 : _GEN_561; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_563 = 7'h46 == _match_key_bytes_2_T_1[6:0] ? phv_data_70 : _GEN_562; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_564 = 7'h47 == _match_key_bytes_2_T_1[6:0] ? phv_data_71 : _GEN_563; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_565 = 7'h48 == _match_key_bytes_2_T_1[6:0] ? phv_data_72 : _GEN_564; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_566 = 7'h49 == _match_key_bytes_2_T_1[6:0] ? phv_data_73 : _GEN_565; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_567 = 7'h4a == _match_key_bytes_2_T_1[6:0] ? phv_data_74 : _GEN_566; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_568 = 7'h4b == _match_key_bytes_2_T_1[6:0] ? phv_data_75 : _GEN_567; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_569 = 7'h4c == _match_key_bytes_2_T_1[6:0] ? phv_data_76 : _GEN_568; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_570 = 7'h4d == _match_key_bytes_2_T_1[6:0] ? phv_data_77 : _GEN_569; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_571 = 7'h4e == _match_key_bytes_2_T_1[6:0] ? phv_data_78 : _GEN_570; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_572 = 7'h4f == _match_key_bytes_2_T_1[6:0] ? phv_data_79 : _GEN_571; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_573 = 7'h50 == _match_key_bytes_2_T_1[6:0] ? phv_data_80 : _GEN_572; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_574 = 7'h51 == _match_key_bytes_2_T_1[6:0] ? phv_data_81 : _GEN_573; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_575 = 7'h52 == _match_key_bytes_2_T_1[6:0] ? phv_data_82 : _GEN_574; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_576 = 7'h53 == _match_key_bytes_2_T_1[6:0] ? phv_data_83 : _GEN_575; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_577 = 7'h54 == _match_key_bytes_2_T_1[6:0] ? phv_data_84 : _GEN_576; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_578 = 7'h55 == _match_key_bytes_2_T_1[6:0] ? phv_data_85 : _GEN_577; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_579 = 7'h56 == _match_key_bytes_2_T_1[6:0] ? phv_data_86 : _GEN_578; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_580 = 7'h57 == _match_key_bytes_2_T_1[6:0] ? phv_data_87 : _GEN_579; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_581 = 7'h58 == _match_key_bytes_2_T_1[6:0] ? phv_data_88 : _GEN_580; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_582 = 7'h59 == _match_key_bytes_2_T_1[6:0] ? phv_data_89 : _GEN_581; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_583 = 7'h5a == _match_key_bytes_2_T_1[6:0] ? phv_data_90 : _GEN_582; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_584 = 7'h5b == _match_key_bytes_2_T_1[6:0] ? phv_data_91 : _GEN_583; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_585 = 7'h5c == _match_key_bytes_2_T_1[6:0] ? phv_data_92 : _GEN_584; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_586 = 7'h5d == _match_key_bytes_2_T_1[6:0] ? phv_data_93 : _GEN_585; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_587 = 7'h5e == _match_key_bytes_2_T_1[6:0] ? phv_data_94 : _GEN_586; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_588 = 7'h5f == _match_key_bytes_2_T_1[6:0] ? phv_data_95 : _GEN_587; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_2 = 4'h5 < _GEN_6 ? _GEN_588 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_1_T_1 = key_offset + 8'h6; // @[matcher.scala 72:98]
  wire [7:0] _GEN_591 = 7'h1 == _match_key_bytes_1_T_1[6:0] ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_592 = 7'h2 == _match_key_bytes_1_T_1[6:0] ? phv_data_2 : _GEN_591; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_593 = 7'h3 == _match_key_bytes_1_T_1[6:0] ? phv_data_3 : _GEN_592; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_594 = 7'h4 == _match_key_bytes_1_T_1[6:0] ? phv_data_4 : _GEN_593; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_595 = 7'h5 == _match_key_bytes_1_T_1[6:0] ? phv_data_5 : _GEN_594; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_596 = 7'h6 == _match_key_bytes_1_T_1[6:0] ? phv_data_6 : _GEN_595; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_597 = 7'h7 == _match_key_bytes_1_T_1[6:0] ? phv_data_7 : _GEN_596; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_598 = 7'h8 == _match_key_bytes_1_T_1[6:0] ? phv_data_8 : _GEN_597; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_599 = 7'h9 == _match_key_bytes_1_T_1[6:0] ? phv_data_9 : _GEN_598; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_600 = 7'ha == _match_key_bytes_1_T_1[6:0] ? phv_data_10 : _GEN_599; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_601 = 7'hb == _match_key_bytes_1_T_1[6:0] ? phv_data_11 : _GEN_600; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_602 = 7'hc == _match_key_bytes_1_T_1[6:0] ? phv_data_12 : _GEN_601; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_603 = 7'hd == _match_key_bytes_1_T_1[6:0] ? phv_data_13 : _GEN_602; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_604 = 7'he == _match_key_bytes_1_T_1[6:0] ? phv_data_14 : _GEN_603; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_605 = 7'hf == _match_key_bytes_1_T_1[6:0] ? phv_data_15 : _GEN_604; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_606 = 7'h10 == _match_key_bytes_1_T_1[6:0] ? phv_data_16 : _GEN_605; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_607 = 7'h11 == _match_key_bytes_1_T_1[6:0] ? phv_data_17 : _GEN_606; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_608 = 7'h12 == _match_key_bytes_1_T_1[6:0] ? phv_data_18 : _GEN_607; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_609 = 7'h13 == _match_key_bytes_1_T_1[6:0] ? phv_data_19 : _GEN_608; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_610 = 7'h14 == _match_key_bytes_1_T_1[6:0] ? phv_data_20 : _GEN_609; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_611 = 7'h15 == _match_key_bytes_1_T_1[6:0] ? phv_data_21 : _GEN_610; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_612 = 7'h16 == _match_key_bytes_1_T_1[6:0] ? phv_data_22 : _GEN_611; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_613 = 7'h17 == _match_key_bytes_1_T_1[6:0] ? phv_data_23 : _GEN_612; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_614 = 7'h18 == _match_key_bytes_1_T_1[6:0] ? phv_data_24 : _GEN_613; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_615 = 7'h19 == _match_key_bytes_1_T_1[6:0] ? phv_data_25 : _GEN_614; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_616 = 7'h1a == _match_key_bytes_1_T_1[6:0] ? phv_data_26 : _GEN_615; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_617 = 7'h1b == _match_key_bytes_1_T_1[6:0] ? phv_data_27 : _GEN_616; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_618 = 7'h1c == _match_key_bytes_1_T_1[6:0] ? phv_data_28 : _GEN_617; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_619 = 7'h1d == _match_key_bytes_1_T_1[6:0] ? phv_data_29 : _GEN_618; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_620 = 7'h1e == _match_key_bytes_1_T_1[6:0] ? phv_data_30 : _GEN_619; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_621 = 7'h1f == _match_key_bytes_1_T_1[6:0] ? phv_data_31 : _GEN_620; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_622 = 7'h20 == _match_key_bytes_1_T_1[6:0] ? phv_data_32 : _GEN_621; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_623 = 7'h21 == _match_key_bytes_1_T_1[6:0] ? phv_data_33 : _GEN_622; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_624 = 7'h22 == _match_key_bytes_1_T_1[6:0] ? phv_data_34 : _GEN_623; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_625 = 7'h23 == _match_key_bytes_1_T_1[6:0] ? phv_data_35 : _GEN_624; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_626 = 7'h24 == _match_key_bytes_1_T_1[6:0] ? phv_data_36 : _GEN_625; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_627 = 7'h25 == _match_key_bytes_1_T_1[6:0] ? phv_data_37 : _GEN_626; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_628 = 7'h26 == _match_key_bytes_1_T_1[6:0] ? phv_data_38 : _GEN_627; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_629 = 7'h27 == _match_key_bytes_1_T_1[6:0] ? phv_data_39 : _GEN_628; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_630 = 7'h28 == _match_key_bytes_1_T_1[6:0] ? phv_data_40 : _GEN_629; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_631 = 7'h29 == _match_key_bytes_1_T_1[6:0] ? phv_data_41 : _GEN_630; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_632 = 7'h2a == _match_key_bytes_1_T_1[6:0] ? phv_data_42 : _GEN_631; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_633 = 7'h2b == _match_key_bytes_1_T_1[6:0] ? phv_data_43 : _GEN_632; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_634 = 7'h2c == _match_key_bytes_1_T_1[6:0] ? phv_data_44 : _GEN_633; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_635 = 7'h2d == _match_key_bytes_1_T_1[6:0] ? phv_data_45 : _GEN_634; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_636 = 7'h2e == _match_key_bytes_1_T_1[6:0] ? phv_data_46 : _GEN_635; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_637 = 7'h2f == _match_key_bytes_1_T_1[6:0] ? phv_data_47 : _GEN_636; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_638 = 7'h30 == _match_key_bytes_1_T_1[6:0] ? phv_data_48 : _GEN_637; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_639 = 7'h31 == _match_key_bytes_1_T_1[6:0] ? phv_data_49 : _GEN_638; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_640 = 7'h32 == _match_key_bytes_1_T_1[6:0] ? phv_data_50 : _GEN_639; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_641 = 7'h33 == _match_key_bytes_1_T_1[6:0] ? phv_data_51 : _GEN_640; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_642 = 7'h34 == _match_key_bytes_1_T_1[6:0] ? phv_data_52 : _GEN_641; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_643 = 7'h35 == _match_key_bytes_1_T_1[6:0] ? phv_data_53 : _GEN_642; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_644 = 7'h36 == _match_key_bytes_1_T_1[6:0] ? phv_data_54 : _GEN_643; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_645 = 7'h37 == _match_key_bytes_1_T_1[6:0] ? phv_data_55 : _GEN_644; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_646 = 7'h38 == _match_key_bytes_1_T_1[6:0] ? phv_data_56 : _GEN_645; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_647 = 7'h39 == _match_key_bytes_1_T_1[6:0] ? phv_data_57 : _GEN_646; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_648 = 7'h3a == _match_key_bytes_1_T_1[6:0] ? phv_data_58 : _GEN_647; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_649 = 7'h3b == _match_key_bytes_1_T_1[6:0] ? phv_data_59 : _GEN_648; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_650 = 7'h3c == _match_key_bytes_1_T_1[6:0] ? phv_data_60 : _GEN_649; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_651 = 7'h3d == _match_key_bytes_1_T_1[6:0] ? phv_data_61 : _GEN_650; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_652 = 7'h3e == _match_key_bytes_1_T_1[6:0] ? phv_data_62 : _GEN_651; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_653 = 7'h3f == _match_key_bytes_1_T_1[6:0] ? phv_data_63 : _GEN_652; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_654 = 7'h40 == _match_key_bytes_1_T_1[6:0] ? phv_data_64 : _GEN_653; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_655 = 7'h41 == _match_key_bytes_1_T_1[6:0] ? phv_data_65 : _GEN_654; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_656 = 7'h42 == _match_key_bytes_1_T_1[6:0] ? phv_data_66 : _GEN_655; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_657 = 7'h43 == _match_key_bytes_1_T_1[6:0] ? phv_data_67 : _GEN_656; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_658 = 7'h44 == _match_key_bytes_1_T_1[6:0] ? phv_data_68 : _GEN_657; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_659 = 7'h45 == _match_key_bytes_1_T_1[6:0] ? phv_data_69 : _GEN_658; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_660 = 7'h46 == _match_key_bytes_1_T_1[6:0] ? phv_data_70 : _GEN_659; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_661 = 7'h47 == _match_key_bytes_1_T_1[6:0] ? phv_data_71 : _GEN_660; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_662 = 7'h48 == _match_key_bytes_1_T_1[6:0] ? phv_data_72 : _GEN_661; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_663 = 7'h49 == _match_key_bytes_1_T_1[6:0] ? phv_data_73 : _GEN_662; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_664 = 7'h4a == _match_key_bytes_1_T_1[6:0] ? phv_data_74 : _GEN_663; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_665 = 7'h4b == _match_key_bytes_1_T_1[6:0] ? phv_data_75 : _GEN_664; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_666 = 7'h4c == _match_key_bytes_1_T_1[6:0] ? phv_data_76 : _GEN_665; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_667 = 7'h4d == _match_key_bytes_1_T_1[6:0] ? phv_data_77 : _GEN_666; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_668 = 7'h4e == _match_key_bytes_1_T_1[6:0] ? phv_data_78 : _GEN_667; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_669 = 7'h4f == _match_key_bytes_1_T_1[6:0] ? phv_data_79 : _GEN_668; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_670 = 7'h50 == _match_key_bytes_1_T_1[6:0] ? phv_data_80 : _GEN_669; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_671 = 7'h51 == _match_key_bytes_1_T_1[6:0] ? phv_data_81 : _GEN_670; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_672 = 7'h52 == _match_key_bytes_1_T_1[6:0] ? phv_data_82 : _GEN_671; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_673 = 7'h53 == _match_key_bytes_1_T_1[6:0] ? phv_data_83 : _GEN_672; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_674 = 7'h54 == _match_key_bytes_1_T_1[6:0] ? phv_data_84 : _GEN_673; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_675 = 7'h55 == _match_key_bytes_1_T_1[6:0] ? phv_data_85 : _GEN_674; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_676 = 7'h56 == _match_key_bytes_1_T_1[6:0] ? phv_data_86 : _GEN_675; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_677 = 7'h57 == _match_key_bytes_1_T_1[6:0] ? phv_data_87 : _GEN_676; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_678 = 7'h58 == _match_key_bytes_1_T_1[6:0] ? phv_data_88 : _GEN_677; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_679 = 7'h59 == _match_key_bytes_1_T_1[6:0] ? phv_data_89 : _GEN_678; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_680 = 7'h5a == _match_key_bytes_1_T_1[6:0] ? phv_data_90 : _GEN_679; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_681 = 7'h5b == _match_key_bytes_1_T_1[6:0] ? phv_data_91 : _GEN_680; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_682 = 7'h5c == _match_key_bytes_1_T_1[6:0] ? phv_data_92 : _GEN_681; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_683 = 7'h5d == _match_key_bytes_1_T_1[6:0] ? phv_data_93 : _GEN_682; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_684 = 7'h5e == _match_key_bytes_1_T_1[6:0] ? phv_data_94 : _GEN_683; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_685 = 7'h5f == _match_key_bytes_1_T_1[6:0] ? phv_data_95 : _GEN_684; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_1 = 4'h6 < _GEN_6 ? _GEN_685 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [7:0] _match_key_bytes_0_T_1 = key_offset + 8'h7; // @[matcher.scala 72:98]
  wire [7:0] _GEN_688 = 7'h1 == _match_key_bytes_0_T_1[6:0] ? phv_data_1 : phv_data_0; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_689 = 7'h2 == _match_key_bytes_0_T_1[6:0] ? phv_data_2 : _GEN_688; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_690 = 7'h3 == _match_key_bytes_0_T_1[6:0] ? phv_data_3 : _GEN_689; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_691 = 7'h4 == _match_key_bytes_0_T_1[6:0] ? phv_data_4 : _GEN_690; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_692 = 7'h5 == _match_key_bytes_0_T_1[6:0] ? phv_data_5 : _GEN_691; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_693 = 7'h6 == _match_key_bytes_0_T_1[6:0] ? phv_data_6 : _GEN_692; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_694 = 7'h7 == _match_key_bytes_0_T_1[6:0] ? phv_data_7 : _GEN_693; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_695 = 7'h8 == _match_key_bytes_0_T_1[6:0] ? phv_data_8 : _GEN_694; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_696 = 7'h9 == _match_key_bytes_0_T_1[6:0] ? phv_data_9 : _GEN_695; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_697 = 7'ha == _match_key_bytes_0_T_1[6:0] ? phv_data_10 : _GEN_696; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_698 = 7'hb == _match_key_bytes_0_T_1[6:0] ? phv_data_11 : _GEN_697; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_699 = 7'hc == _match_key_bytes_0_T_1[6:0] ? phv_data_12 : _GEN_698; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_700 = 7'hd == _match_key_bytes_0_T_1[6:0] ? phv_data_13 : _GEN_699; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_701 = 7'he == _match_key_bytes_0_T_1[6:0] ? phv_data_14 : _GEN_700; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_702 = 7'hf == _match_key_bytes_0_T_1[6:0] ? phv_data_15 : _GEN_701; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_703 = 7'h10 == _match_key_bytes_0_T_1[6:0] ? phv_data_16 : _GEN_702; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_704 = 7'h11 == _match_key_bytes_0_T_1[6:0] ? phv_data_17 : _GEN_703; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_705 = 7'h12 == _match_key_bytes_0_T_1[6:0] ? phv_data_18 : _GEN_704; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_706 = 7'h13 == _match_key_bytes_0_T_1[6:0] ? phv_data_19 : _GEN_705; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_707 = 7'h14 == _match_key_bytes_0_T_1[6:0] ? phv_data_20 : _GEN_706; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_708 = 7'h15 == _match_key_bytes_0_T_1[6:0] ? phv_data_21 : _GEN_707; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_709 = 7'h16 == _match_key_bytes_0_T_1[6:0] ? phv_data_22 : _GEN_708; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_710 = 7'h17 == _match_key_bytes_0_T_1[6:0] ? phv_data_23 : _GEN_709; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_711 = 7'h18 == _match_key_bytes_0_T_1[6:0] ? phv_data_24 : _GEN_710; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_712 = 7'h19 == _match_key_bytes_0_T_1[6:0] ? phv_data_25 : _GEN_711; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_713 = 7'h1a == _match_key_bytes_0_T_1[6:0] ? phv_data_26 : _GEN_712; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_714 = 7'h1b == _match_key_bytes_0_T_1[6:0] ? phv_data_27 : _GEN_713; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_715 = 7'h1c == _match_key_bytes_0_T_1[6:0] ? phv_data_28 : _GEN_714; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_716 = 7'h1d == _match_key_bytes_0_T_1[6:0] ? phv_data_29 : _GEN_715; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_717 = 7'h1e == _match_key_bytes_0_T_1[6:0] ? phv_data_30 : _GEN_716; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_718 = 7'h1f == _match_key_bytes_0_T_1[6:0] ? phv_data_31 : _GEN_717; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_719 = 7'h20 == _match_key_bytes_0_T_1[6:0] ? phv_data_32 : _GEN_718; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_720 = 7'h21 == _match_key_bytes_0_T_1[6:0] ? phv_data_33 : _GEN_719; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_721 = 7'h22 == _match_key_bytes_0_T_1[6:0] ? phv_data_34 : _GEN_720; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_722 = 7'h23 == _match_key_bytes_0_T_1[6:0] ? phv_data_35 : _GEN_721; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_723 = 7'h24 == _match_key_bytes_0_T_1[6:0] ? phv_data_36 : _GEN_722; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_724 = 7'h25 == _match_key_bytes_0_T_1[6:0] ? phv_data_37 : _GEN_723; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_725 = 7'h26 == _match_key_bytes_0_T_1[6:0] ? phv_data_38 : _GEN_724; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_726 = 7'h27 == _match_key_bytes_0_T_1[6:0] ? phv_data_39 : _GEN_725; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_727 = 7'h28 == _match_key_bytes_0_T_1[6:0] ? phv_data_40 : _GEN_726; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_728 = 7'h29 == _match_key_bytes_0_T_1[6:0] ? phv_data_41 : _GEN_727; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_729 = 7'h2a == _match_key_bytes_0_T_1[6:0] ? phv_data_42 : _GEN_728; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_730 = 7'h2b == _match_key_bytes_0_T_1[6:0] ? phv_data_43 : _GEN_729; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_731 = 7'h2c == _match_key_bytes_0_T_1[6:0] ? phv_data_44 : _GEN_730; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_732 = 7'h2d == _match_key_bytes_0_T_1[6:0] ? phv_data_45 : _GEN_731; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_733 = 7'h2e == _match_key_bytes_0_T_1[6:0] ? phv_data_46 : _GEN_732; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_734 = 7'h2f == _match_key_bytes_0_T_1[6:0] ? phv_data_47 : _GEN_733; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_735 = 7'h30 == _match_key_bytes_0_T_1[6:0] ? phv_data_48 : _GEN_734; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_736 = 7'h31 == _match_key_bytes_0_T_1[6:0] ? phv_data_49 : _GEN_735; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_737 = 7'h32 == _match_key_bytes_0_T_1[6:0] ? phv_data_50 : _GEN_736; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_738 = 7'h33 == _match_key_bytes_0_T_1[6:0] ? phv_data_51 : _GEN_737; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_739 = 7'h34 == _match_key_bytes_0_T_1[6:0] ? phv_data_52 : _GEN_738; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_740 = 7'h35 == _match_key_bytes_0_T_1[6:0] ? phv_data_53 : _GEN_739; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_741 = 7'h36 == _match_key_bytes_0_T_1[6:0] ? phv_data_54 : _GEN_740; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_742 = 7'h37 == _match_key_bytes_0_T_1[6:0] ? phv_data_55 : _GEN_741; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_743 = 7'h38 == _match_key_bytes_0_T_1[6:0] ? phv_data_56 : _GEN_742; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_744 = 7'h39 == _match_key_bytes_0_T_1[6:0] ? phv_data_57 : _GEN_743; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_745 = 7'h3a == _match_key_bytes_0_T_1[6:0] ? phv_data_58 : _GEN_744; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_746 = 7'h3b == _match_key_bytes_0_T_1[6:0] ? phv_data_59 : _GEN_745; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_747 = 7'h3c == _match_key_bytes_0_T_1[6:0] ? phv_data_60 : _GEN_746; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_748 = 7'h3d == _match_key_bytes_0_T_1[6:0] ? phv_data_61 : _GEN_747; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_749 = 7'h3e == _match_key_bytes_0_T_1[6:0] ? phv_data_62 : _GEN_748; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_750 = 7'h3f == _match_key_bytes_0_T_1[6:0] ? phv_data_63 : _GEN_749; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_751 = 7'h40 == _match_key_bytes_0_T_1[6:0] ? phv_data_64 : _GEN_750; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_752 = 7'h41 == _match_key_bytes_0_T_1[6:0] ? phv_data_65 : _GEN_751; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_753 = 7'h42 == _match_key_bytes_0_T_1[6:0] ? phv_data_66 : _GEN_752; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_754 = 7'h43 == _match_key_bytes_0_T_1[6:0] ? phv_data_67 : _GEN_753; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_755 = 7'h44 == _match_key_bytes_0_T_1[6:0] ? phv_data_68 : _GEN_754; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_756 = 7'h45 == _match_key_bytes_0_T_1[6:0] ? phv_data_69 : _GEN_755; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_757 = 7'h46 == _match_key_bytes_0_T_1[6:0] ? phv_data_70 : _GEN_756; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_758 = 7'h47 == _match_key_bytes_0_T_1[6:0] ? phv_data_71 : _GEN_757; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_759 = 7'h48 == _match_key_bytes_0_T_1[6:0] ? phv_data_72 : _GEN_758; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_760 = 7'h49 == _match_key_bytes_0_T_1[6:0] ? phv_data_73 : _GEN_759; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_761 = 7'h4a == _match_key_bytes_0_T_1[6:0] ? phv_data_74 : _GEN_760; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_762 = 7'h4b == _match_key_bytes_0_T_1[6:0] ? phv_data_75 : _GEN_761; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_763 = 7'h4c == _match_key_bytes_0_T_1[6:0] ? phv_data_76 : _GEN_762; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_764 = 7'h4d == _match_key_bytes_0_T_1[6:0] ? phv_data_77 : _GEN_763; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_765 = 7'h4e == _match_key_bytes_0_T_1[6:0] ? phv_data_78 : _GEN_764; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_766 = 7'h4f == _match_key_bytes_0_T_1[6:0] ? phv_data_79 : _GEN_765; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_767 = 7'h50 == _match_key_bytes_0_T_1[6:0] ? phv_data_80 : _GEN_766; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_768 = 7'h51 == _match_key_bytes_0_T_1[6:0] ? phv_data_81 : _GEN_767; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_769 = 7'h52 == _match_key_bytes_0_T_1[6:0] ? phv_data_82 : _GEN_768; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_770 = 7'h53 == _match_key_bytes_0_T_1[6:0] ? phv_data_83 : _GEN_769; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_771 = 7'h54 == _match_key_bytes_0_T_1[6:0] ? phv_data_84 : _GEN_770; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_772 = 7'h55 == _match_key_bytes_0_T_1[6:0] ? phv_data_85 : _GEN_771; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_773 = 7'h56 == _match_key_bytes_0_T_1[6:0] ? phv_data_86 : _GEN_772; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_774 = 7'h57 == _match_key_bytes_0_T_1[6:0] ? phv_data_87 : _GEN_773; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_775 = 7'h58 == _match_key_bytes_0_T_1[6:0] ? phv_data_88 : _GEN_774; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_776 = 7'h59 == _match_key_bytes_0_T_1[6:0] ? phv_data_89 : _GEN_775; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_777 = 7'h5a == _match_key_bytes_0_T_1[6:0] ? phv_data_90 : _GEN_776; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_778 = 7'h5b == _match_key_bytes_0_T_1[6:0] ? phv_data_91 : _GEN_777; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_779 = 7'h5c == _match_key_bytes_0_T_1[6:0] ? phv_data_92 : _GEN_778; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_780 = 7'h5d == _match_key_bytes_0_T_1[6:0] ? phv_data_93 : _GEN_779; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_781 = 7'h5e == _match_key_bytes_0_T_1[6:0] ? phv_data_94 : _GEN_780; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] _GEN_782 = 7'h5f == _match_key_bytes_0_T_1[6:0] ? phv_data_95 : _GEN_781; // @[matcher.scala 72:75 matcher.scala 72:75]
  wire [7:0] match_key_bytes_0 = 4'h7 < _GEN_6 ? _GEN_782 : 8'h0; // @[matcher.scala 71:84 matcher.scala 72:75 matcher.scala 74:75]
  wire [63:0] match_key = {match_key_bytes_0,match_key_bytes_1,match_key_bytes_2,match_key_bytes_3,match_key_bytes_4,
    match_key_bytes_5,match_key_bytes_6,match_key_bytes_7}; // @[Cat.scala 30:58]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[matcher.scala 60:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[matcher.scala 60:25]
  assign io_match_key = phv_is_valid_processor ? match_key : 64'h0; // @[matcher.scala 65:39 matcher.scala 79:26 matcher.scala 81:26]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[matcher.scala 59:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[matcher.scala 59:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[matcher.scala 59:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[matcher.scala 59:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[matcher.scala 59:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[matcher.scala 59:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[matcher.scala 59:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[matcher.scala 59:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[matcher.scala 59:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[matcher.scala 59:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[matcher.scala 59:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[matcher.scala 59:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[matcher.scala 59:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[matcher.scala 59:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[matcher.scala 59:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[matcher.scala 59:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[matcher.scala 59:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[matcher.scala 59:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[matcher.scala 59:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[matcher.scala 59:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[matcher.scala 59:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[matcher.scala 59:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[matcher.scala 59:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[matcher.scala 59:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[matcher.scala 59:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[matcher.scala 59:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[matcher.scala 59:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[matcher.scala 59:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[matcher.scala 59:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[matcher.scala 59:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[matcher.scala 59:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[matcher.scala 59:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[matcher.scala 59:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[matcher.scala 59:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[matcher.scala 59:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[matcher.scala 59:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[matcher.scala 59:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[matcher.scala 59:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[matcher.scala 59:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[matcher.scala 59:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[matcher.scala 59:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[matcher.scala 59:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[matcher.scala 59:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[matcher.scala 59:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[matcher.scala 59:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[matcher.scala 59:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[matcher.scala 59:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[matcher.scala 59:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[matcher.scala 59:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[matcher.scala 59:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[matcher.scala 59:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[matcher.scala 59:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[matcher.scala 59:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[matcher.scala 59:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[matcher.scala 59:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[matcher.scala 59:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[matcher.scala 59:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[matcher.scala 59:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[matcher.scala 59:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[matcher.scala 59:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[matcher.scala 59:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[matcher.scala 59:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[matcher.scala 59:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[matcher.scala 59:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[matcher.scala 59:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[matcher.scala 59:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[matcher.scala 59:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[matcher.scala 59:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[matcher.scala 59:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[matcher.scala 59:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[matcher.scala 59:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[matcher.scala 59:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[matcher.scala 59:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[matcher.scala 59:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[matcher.scala 59:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[matcher.scala 59:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[matcher.scala 59:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[matcher.scala 59:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[matcher.scala 59:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[matcher.scala 59:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[matcher.scala 59:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[matcher.scala 59:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[matcher.scala 59:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[matcher.scala 59:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[matcher.scala 59:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[matcher.scala 59:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[matcher.scala 59:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[matcher.scala 59:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[matcher.scala 59:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[matcher.scala 59:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[matcher.scala 59:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[matcher.scala 59:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[matcher.scala 59:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[matcher.scala 59:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[matcher.scala 59:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[matcher.scala 59:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[matcher.scala 59:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[matcher.scala 59:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[matcher.scala 59:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[matcher.scala 59:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[matcher.scala 59:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[matcher.scala 59:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[matcher.scala 59:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[matcher.scala 59:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[matcher.scala 59:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[matcher.scala 59:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[matcher.scala 59:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[matcher.scala 59:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[matcher.scala 59:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[matcher.scala 59:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[matcher.scala 59:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[matcher.scala 59:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[matcher.scala 59:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[matcher.scala 59:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[matcher.scala 59:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[matcher.scala 59:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[matcher.scala 59:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[matcher.scala 59:13]
    key_offset <= io_key_offset; // @[matcher.scala 63:20]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  phv_next_config_id = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  key_offset = _RAND_118[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HashSumLevel(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input  [63:0] io_key_in,
  output [63:0] io_key_out,
  input  [15:0] io_sum_in,
  output [15:0] io_sum_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [31:0] _RAND_119;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[hash.scala 37:22]
  reg [7:0] phv_data_1; // @[hash.scala 37:22]
  reg [7:0] phv_data_2; // @[hash.scala 37:22]
  reg [7:0] phv_data_3; // @[hash.scala 37:22]
  reg [7:0] phv_data_4; // @[hash.scala 37:22]
  reg [7:0] phv_data_5; // @[hash.scala 37:22]
  reg [7:0] phv_data_6; // @[hash.scala 37:22]
  reg [7:0] phv_data_7; // @[hash.scala 37:22]
  reg [7:0] phv_data_8; // @[hash.scala 37:22]
  reg [7:0] phv_data_9; // @[hash.scala 37:22]
  reg [7:0] phv_data_10; // @[hash.scala 37:22]
  reg [7:0] phv_data_11; // @[hash.scala 37:22]
  reg [7:0] phv_data_12; // @[hash.scala 37:22]
  reg [7:0] phv_data_13; // @[hash.scala 37:22]
  reg [7:0] phv_data_14; // @[hash.scala 37:22]
  reg [7:0] phv_data_15; // @[hash.scala 37:22]
  reg [7:0] phv_data_16; // @[hash.scala 37:22]
  reg [7:0] phv_data_17; // @[hash.scala 37:22]
  reg [7:0] phv_data_18; // @[hash.scala 37:22]
  reg [7:0] phv_data_19; // @[hash.scala 37:22]
  reg [7:0] phv_data_20; // @[hash.scala 37:22]
  reg [7:0] phv_data_21; // @[hash.scala 37:22]
  reg [7:0] phv_data_22; // @[hash.scala 37:22]
  reg [7:0] phv_data_23; // @[hash.scala 37:22]
  reg [7:0] phv_data_24; // @[hash.scala 37:22]
  reg [7:0] phv_data_25; // @[hash.scala 37:22]
  reg [7:0] phv_data_26; // @[hash.scala 37:22]
  reg [7:0] phv_data_27; // @[hash.scala 37:22]
  reg [7:0] phv_data_28; // @[hash.scala 37:22]
  reg [7:0] phv_data_29; // @[hash.scala 37:22]
  reg [7:0] phv_data_30; // @[hash.scala 37:22]
  reg [7:0] phv_data_31; // @[hash.scala 37:22]
  reg [7:0] phv_data_32; // @[hash.scala 37:22]
  reg [7:0] phv_data_33; // @[hash.scala 37:22]
  reg [7:0] phv_data_34; // @[hash.scala 37:22]
  reg [7:0] phv_data_35; // @[hash.scala 37:22]
  reg [7:0] phv_data_36; // @[hash.scala 37:22]
  reg [7:0] phv_data_37; // @[hash.scala 37:22]
  reg [7:0] phv_data_38; // @[hash.scala 37:22]
  reg [7:0] phv_data_39; // @[hash.scala 37:22]
  reg [7:0] phv_data_40; // @[hash.scala 37:22]
  reg [7:0] phv_data_41; // @[hash.scala 37:22]
  reg [7:0] phv_data_42; // @[hash.scala 37:22]
  reg [7:0] phv_data_43; // @[hash.scala 37:22]
  reg [7:0] phv_data_44; // @[hash.scala 37:22]
  reg [7:0] phv_data_45; // @[hash.scala 37:22]
  reg [7:0] phv_data_46; // @[hash.scala 37:22]
  reg [7:0] phv_data_47; // @[hash.scala 37:22]
  reg [7:0] phv_data_48; // @[hash.scala 37:22]
  reg [7:0] phv_data_49; // @[hash.scala 37:22]
  reg [7:0] phv_data_50; // @[hash.scala 37:22]
  reg [7:0] phv_data_51; // @[hash.scala 37:22]
  reg [7:0] phv_data_52; // @[hash.scala 37:22]
  reg [7:0] phv_data_53; // @[hash.scala 37:22]
  reg [7:0] phv_data_54; // @[hash.scala 37:22]
  reg [7:0] phv_data_55; // @[hash.scala 37:22]
  reg [7:0] phv_data_56; // @[hash.scala 37:22]
  reg [7:0] phv_data_57; // @[hash.scala 37:22]
  reg [7:0] phv_data_58; // @[hash.scala 37:22]
  reg [7:0] phv_data_59; // @[hash.scala 37:22]
  reg [7:0] phv_data_60; // @[hash.scala 37:22]
  reg [7:0] phv_data_61; // @[hash.scala 37:22]
  reg [7:0] phv_data_62; // @[hash.scala 37:22]
  reg [7:0] phv_data_63; // @[hash.scala 37:22]
  reg [7:0] phv_data_64; // @[hash.scala 37:22]
  reg [7:0] phv_data_65; // @[hash.scala 37:22]
  reg [7:0] phv_data_66; // @[hash.scala 37:22]
  reg [7:0] phv_data_67; // @[hash.scala 37:22]
  reg [7:0] phv_data_68; // @[hash.scala 37:22]
  reg [7:0] phv_data_69; // @[hash.scala 37:22]
  reg [7:0] phv_data_70; // @[hash.scala 37:22]
  reg [7:0] phv_data_71; // @[hash.scala 37:22]
  reg [7:0] phv_data_72; // @[hash.scala 37:22]
  reg [7:0] phv_data_73; // @[hash.scala 37:22]
  reg [7:0] phv_data_74; // @[hash.scala 37:22]
  reg [7:0] phv_data_75; // @[hash.scala 37:22]
  reg [7:0] phv_data_76; // @[hash.scala 37:22]
  reg [7:0] phv_data_77; // @[hash.scala 37:22]
  reg [7:0] phv_data_78; // @[hash.scala 37:22]
  reg [7:0] phv_data_79; // @[hash.scala 37:22]
  reg [7:0] phv_data_80; // @[hash.scala 37:22]
  reg [7:0] phv_data_81; // @[hash.scala 37:22]
  reg [7:0] phv_data_82; // @[hash.scala 37:22]
  reg [7:0] phv_data_83; // @[hash.scala 37:22]
  reg [7:0] phv_data_84; // @[hash.scala 37:22]
  reg [7:0] phv_data_85; // @[hash.scala 37:22]
  reg [7:0] phv_data_86; // @[hash.scala 37:22]
  reg [7:0] phv_data_87; // @[hash.scala 37:22]
  reg [7:0] phv_data_88; // @[hash.scala 37:22]
  reg [7:0] phv_data_89; // @[hash.scala 37:22]
  reg [7:0] phv_data_90; // @[hash.scala 37:22]
  reg [7:0] phv_data_91; // @[hash.scala 37:22]
  reg [7:0] phv_data_92; // @[hash.scala 37:22]
  reg [7:0] phv_data_93; // @[hash.scala 37:22]
  reg [7:0] phv_data_94; // @[hash.scala 37:22]
  reg [7:0] phv_data_95; // @[hash.scala 37:22]
  reg [15:0] phv_header_0; // @[hash.scala 37:22]
  reg [15:0] phv_header_1; // @[hash.scala 37:22]
  reg [15:0] phv_header_2; // @[hash.scala 37:22]
  reg [15:0] phv_header_3; // @[hash.scala 37:22]
  reg [15:0] phv_header_4; // @[hash.scala 37:22]
  reg [15:0] phv_header_5; // @[hash.scala 37:22]
  reg [15:0] phv_header_6; // @[hash.scala 37:22]
  reg [15:0] phv_header_7; // @[hash.scala 37:22]
  reg [15:0] phv_header_8; // @[hash.scala 37:22]
  reg [15:0] phv_header_9; // @[hash.scala 37:22]
  reg [15:0] phv_header_10; // @[hash.scala 37:22]
  reg [15:0] phv_header_11; // @[hash.scala 37:22]
  reg [15:0] phv_header_12; // @[hash.scala 37:22]
  reg [15:0] phv_header_13; // @[hash.scala 37:22]
  reg [15:0] phv_header_14; // @[hash.scala 37:22]
  reg [15:0] phv_header_15; // @[hash.scala 37:22]
  reg [7:0] phv_parse_current_state; // @[hash.scala 37:22]
  reg [7:0] phv_parse_current_offset; // @[hash.scala 37:22]
  reg [15:0] phv_parse_transition_field; // @[hash.scala 37:22]
  reg [1:0] phv_next_processor_id; // @[hash.scala 37:22]
  reg  phv_next_config_id; // @[hash.scala 37:22]
  reg  phv_is_valid_processor; // @[hash.scala 37:22]
  reg [63:0] key; // @[hash.scala 41:22]
  reg [15:0] sum; // @[hash.scala 45:22]
  wire [15:0] _io_sum_out_T_2 = sum + key[31:16]; // @[hash.scala 49:31]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[hash.scala 39:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[hash.scala 39:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[hash.scala 39:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[hash.scala 39:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[hash.scala 39:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[hash.scala 39:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[hash.scala 39:25]
  assign io_key_out = key; // @[hash.scala 43:20]
  assign io_sum_out = phv_is_valid_processor ? _io_sum_out_T_2 : sum; // @[hash.scala 48:39 hash.scala 49:24 hash.scala 51:24]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[hash.scala 38:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[hash.scala 38:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[hash.scala 38:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[hash.scala 38:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[hash.scala 38:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[hash.scala 38:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[hash.scala 38:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[hash.scala 38:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[hash.scala 38:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[hash.scala 38:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[hash.scala 38:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[hash.scala 38:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[hash.scala 38:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[hash.scala 38:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[hash.scala 38:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[hash.scala 38:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[hash.scala 38:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[hash.scala 38:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[hash.scala 38:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[hash.scala 38:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[hash.scala 38:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[hash.scala 38:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[hash.scala 38:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[hash.scala 38:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[hash.scala 38:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[hash.scala 38:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[hash.scala 38:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[hash.scala 38:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[hash.scala 38:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[hash.scala 38:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[hash.scala 38:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[hash.scala 38:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[hash.scala 38:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[hash.scala 38:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[hash.scala 38:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[hash.scala 38:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[hash.scala 38:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[hash.scala 38:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[hash.scala 38:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[hash.scala 38:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[hash.scala 38:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[hash.scala 38:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[hash.scala 38:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[hash.scala 38:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[hash.scala 38:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[hash.scala 38:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[hash.scala 38:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[hash.scala 38:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[hash.scala 38:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[hash.scala 38:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[hash.scala 38:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[hash.scala 38:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[hash.scala 38:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[hash.scala 38:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[hash.scala 38:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[hash.scala 38:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[hash.scala 38:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[hash.scala 38:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[hash.scala 38:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[hash.scala 38:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[hash.scala 38:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[hash.scala 38:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[hash.scala 38:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[hash.scala 38:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[hash.scala 38:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[hash.scala 38:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[hash.scala 38:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[hash.scala 38:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[hash.scala 38:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[hash.scala 38:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[hash.scala 38:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[hash.scala 38:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[hash.scala 38:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[hash.scala 38:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[hash.scala 38:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[hash.scala 38:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[hash.scala 38:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[hash.scala 38:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[hash.scala 38:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[hash.scala 38:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[hash.scala 38:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[hash.scala 38:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[hash.scala 38:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[hash.scala 38:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[hash.scala 38:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[hash.scala 38:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[hash.scala 38:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[hash.scala 38:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[hash.scala 38:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[hash.scala 38:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[hash.scala 38:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[hash.scala 38:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[hash.scala 38:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[hash.scala 38:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[hash.scala 38:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[hash.scala 38:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[hash.scala 38:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[hash.scala 38:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[hash.scala 38:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[hash.scala 38:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[hash.scala 38:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[hash.scala 38:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[hash.scala 38:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[hash.scala 38:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[hash.scala 38:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[hash.scala 38:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[hash.scala 38:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[hash.scala 38:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[hash.scala 38:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[hash.scala 38:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[hash.scala 38:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[hash.scala 38:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[hash.scala 38:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[hash.scala 38:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[hash.scala 38:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[hash.scala 38:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[hash.scala 38:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[hash.scala 38:13]
    key <= io_key_in; // @[hash.scala 42:13]
    sum <= io_sum_in; // @[hash.scala 46:13]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  phv_next_config_id = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_117[0:0];
  _RAND_118 = {2{`RANDOM}};
  key = _RAND_118[63:0];
  _RAND_119 = {1{`RANDOM}};
  sum = _RAND_119[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HashSumLevel_1(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input  [63:0] io_key_in,
  output [63:0] io_key_out,
  input  [15:0] io_sum_in,
  output [15:0] io_sum_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [31:0] _RAND_119;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[hash.scala 37:22]
  reg [7:0] phv_data_1; // @[hash.scala 37:22]
  reg [7:0] phv_data_2; // @[hash.scala 37:22]
  reg [7:0] phv_data_3; // @[hash.scala 37:22]
  reg [7:0] phv_data_4; // @[hash.scala 37:22]
  reg [7:0] phv_data_5; // @[hash.scala 37:22]
  reg [7:0] phv_data_6; // @[hash.scala 37:22]
  reg [7:0] phv_data_7; // @[hash.scala 37:22]
  reg [7:0] phv_data_8; // @[hash.scala 37:22]
  reg [7:0] phv_data_9; // @[hash.scala 37:22]
  reg [7:0] phv_data_10; // @[hash.scala 37:22]
  reg [7:0] phv_data_11; // @[hash.scala 37:22]
  reg [7:0] phv_data_12; // @[hash.scala 37:22]
  reg [7:0] phv_data_13; // @[hash.scala 37:22]
  reg [7:0] phv_data_14; // @[hash.scala 37:22]
  reg [7:0] phv_data_15; // @[hash.scala 37:22]
  reg [7:0] phv_data_16; // @[hash.scala 37:22]
  reg [7:0] phv_data_17; // @[hash.scala 37:22]
  reg [7:0] phv_data_18; // @[hash.scala 37:22]
  reg [7:0] phv_data_19; // @[hash.scala 37:22]
  reg [7:0] phv_data_20; // @[hash.scala 37:22]
  reg [7:0] phv_data_21; // @[hash.scala 37:22]
  reg [7:0] phv_data_22; // @[hash.scala 37:22]
  reg [7:0] phv_data_23; // @[hash.scala 37:22]
  reg [7:0] phv_data_24; // @[hash.scala 37:22]
  reg [7:0] phv_data_25; // @[hash.scala 37:22]
  reg [7:0] phv_data_26; // @[hash.scala 37:22]
  reg [7:0] phv_data_27; // @[hash.scala 37:22]
  reg [7:0] phv_data_28; // @[hash.scala 37:22]
  reg [7:0] phv_data_29; // @[hash.scala 37:22]
  reg [7:0] phv_data_30; // @[hash.scala 37:22]
  reg [7:0] phv_data_31; // @[hash.scala 37:22]
  reg [7:0] phv_data_32; // @[hash.scala 37:22]
  reg [7:0] phv_data_33; // @[hash.scala 37:22]
  reg [7:0] phv_data_34; // @[hash.scala 37:22]
  reg [7:0] phv_data_35; // @[hash.scala 37:22]
  reg [7:0] phv_data_36; // @[hash.scala 37:22]
  reg [7:0] phv_data_37; // @[hash.scala 37:22]
  reg [7:0] phv_data_38; // @[hash.scala 37:22]
  reg [7:0] phv_data_39; // @[hash.scala 37:22]
  reg [7:0] phv_data_40; // @[hash.scala 37:22]
  reg [7:0] phv_data_41; // @[hash.scala 37:22]
  reg [7:0] phv_data_42; // @[hash.scala 37:22]
  reg [7:0] phv_data_43; // @[hash.scala 37:22]
  reg [7:0] phv_data_44; // @[hash.scala 37:22]
  reg [7:0] phv_data_45; // @[hash.scala 37:22]
  reg [7:0] phv_data_46; // @[hash.scala 37:22]
  reg [7:0] phv_data_47; // @[hash.scala 37:22]
  reg [7:0] phv_data_48; // @[hash.scala 37:22]
  reg [7:0] phv_data_49; // @[hash.scala 37:22]
  reg [7:0] phv_data_50; // @[hash.scala 37:22]
  reg [7:0] phv_data_51; // @[hash.scala 37:22]
  reg [7:0] phv_data_52; // @[hash.scala 37:22]
  reg [7:0] phv_data_53; // @[hash.scala 37:22]
  reg [7:0] phv_data_54; // @[hash.scala 37:22]
  reg [7:0] phv_data_55; // @[hash.scala 37:22]
  reg [7:0] phv_data_56; // @[hash.scala 37:22]
  reg [7:0] phv_data_57; // @[hash.scala 37:22]
  reg [7:0] phv_data_58; // @[hash.scala 37:22]
  reg [7:0] phv_data_59; // @[hash.scala 37:22]
  reg [7:0] phv_data_60; // @[hash.scala 37:22]
  reg [7:0] phv_data_61; // @[hash.scala 37:22]
  reg [7:0] phv_data_62; // @[hash.scala 37:22]
  reg [7:0] phv_data_63; // @[hash.scala 37:22]
  reg [7:0] phv_data_64; // @[hash.scala 37:22]
  reg [7:0] phv_data_65; // @[hash.scala 37:22]
  reg [7:0] phv_data_66; // @[hash.scala 37:22]
  reg [7:0] phv_data_67; // @[hash.scala 37:22]
  reg [7:0] phv_data_68; // @[hash.scala 37:22]
  reg [7:0] phv_data_69; // @[hash.scala 37:22]
  reg [7:0] phv_data_70; // @[hash.scala 37:22]
  reg [7:0] phv_data_71; // @[hash.scala 37:22]
  reg [7:0] phv_data_72; // @[hash.scala 37:22]
  reg [7:0] phv_data_73; // @[hash.scala 37:22]
  reg [7:0] phv_data_74; // @[hash.scala 37:22]
  reg [7:0] phv_data_75; // @[hash.scala 37:22]
  reg [7:0] phv_data_76; // @[hash.scala 37:22]
  reg [7:0] phv_data_77; // @[hash.scala 37:22]
  reg [7:0] phv_data_78; // @[hash.scala 37:22]
  reg [7:0] phv_data_79; // @[hash.scala 37:22]
  reg [7:0] phv_data_80; // @[hash.scala 37:22]
  reg [7:0] phv_data_81; // @[hash.scala 37:22]
  reg [7:0] phv_data_82; // @[hash.scala 37:22]
  reg [7:0] phv_data_83; // @[hash.scala 37:22]
  reg [7:0] phv_data_84; // @[hash.scala 37:22]
  reg [7:0] phv_data_85; // @[hash.scala 37:22]
  reg [7:0] phv_data_86; // @[hash.scala 37:22]
  reg [7:0] phv_data_87; // @[hash.scala 37:22]
  reg [7:0] phv_data_88; // @[hash.scala 37:22]
  reg [7:0] phv_data_89; // @[hash.scala 37:22]
  reg [7:0] phv_data_90; // @[hash.scala 37:22]
  reg [7:0] phv_data_91; // @[hash.scala 37:22]
  reg [7:0] phv_data_92; // @[hash.scala 37:22]
  reg [7:0] phv_data_93; // @[hash.scala 37:22]
  reg [7:0] phv_data_94; // @[hash.scala 37:22]
  reg [7:0] phv_data_95; // @[hash.scala 37:22]
  reg [15:0] phv_header_0; // @[hash.scala 37:22]
  reg [15:0] phv_header_1; // @[hash.scala 37:22]
  reg [15:0] phv_header_2; // @[hash.scala 37:22]
  reg [15:0] phv_header_3; // @[hash.scala 37:22]
  reg [15:0] phv_header_4; // @[hash.scala 37:22]
  reg [15:0] phv_header_5; // @[hash.scala 37:22]
  reg [15:0] phv_header_6; // @[hash.scala 37:22]
  reg [15:0] phv_header_7; // @[hash.scala 37:22]
  reg [15:0] phv_header_8; // @[hash.scala 37:22]
  reg [15:0] phv_header_9; // @[hash.scala 37:22]
  reg [15:0] phv_header_10; // @[hash.scala 37:22]
  reg [15:0] phv_header_11; // @[hash.scala 37:22]
  reg [15:0] phv_header_12; // @[hash.scala 37:22]
  reg [15:0] phv_header_13; // @[hash.scala 37:22]
  reg [15:0] phv_header_14; // @[hash.scala 37:22]
  reg [15:0] phv_header_15; // @[hash.scala 37:22]
  reg [7:0] phv_parse_current_state; // @[hash.scala 37:22]
  reg [7:0] phv_parse_current_offset; // @[hash.scala 37:22]
  reg [15:0] phv_parse_transition_field; // @[hash.scala 37:22]
  reg [1:0] phv_next_processor_id; // @[hash.scala 37:22]
  reg  phv_next_config_id; // @[hash.scala 37:22]
  reg  phv_is_valid_processor; // @[hash.scala 37:22]
  reg [63:0] key; // @[hash.scala 41:22]
  reg [15:0] sum; // @[hash.scala 45:22]
  wire [15:0] _io_sum_out_T_2 = sum + key[47:32]; // @[hash.scala 49:31]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[hash.scala 39:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[hash.scala 39:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[hash.scala 39:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[hash.scala 39:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[hash.scala 39:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[hash.scala 39:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[hash.scala 39:25]
  assign io_key_out = key; // @[hash.scala 43:20]
  assign io_sum_out = phv_is_valid_processor ? _io_sum_out_T_2 : sum; // @[hash.scala 48:39 hash.scala 49:24 hash.scala 51:24]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[hash.scala 38:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[hash.scala 38:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[hash.scala 38:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[hash.scala 38:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[hash.scala 38:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[hash.scala 38:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[hash.scala 38:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[hash.scala 38:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[hash.scala 38:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[hash.scala 38:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[hash.scala 38:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[hash.scala 38:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[hash.scala 38:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[hash.scala 38:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[hash.scala 38:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[hash.scala 38:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[hash.scala 38:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[hash.scala 38:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[hash.scala 38:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[hash.scala 38:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[hash.scala 38:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[hash.scala 38:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[hash.scala 38:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[hash.scala 38:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[hash.scala 38:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[hash.scala 38:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[hash.scala 38:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[hash.scala 38:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[hash.scala 38:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[hash.scala 38:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[hash.scala 38:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[hash.scala 38:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[hash.scala 38:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[hash.scala 38:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[hash.scala 38:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[hash.scala 38:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[hash.scala 38:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[hash.scala 38:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[hash.scala 38:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[hash.scala 38:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[hash.scala 38:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[hash.scala 38:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[hash.scala 38:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[hash.scala 38:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[hash.scala 38:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[hash.scala 38:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[hash.scala 38:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[hash.scala 38:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[hash.scala 38:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[hash.scala 38:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[hash.scala 38:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[hash.scala 38:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[hash.scala 38:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[hash.scala 38:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[hash.scala 38:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[hash.scala 38:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[hash.scala 38:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[hash.scala 38:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[hash.scala 38:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[hash.scala 38:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[hash.scala 38:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[hash.scala 38:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[hash.scala 38:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[hash.scala 38:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[hash.scala 38:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[hash.scala 38:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[hash.scala 38:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[hash.scala 38:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[hash.scala 38:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[hash.scala 38:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[hash.scala 38:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[hash.scala 38:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[hash.scala 38:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[hash.scala 38:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[hash.scala 38:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[hash.scala 38:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[hash.scala 38:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[hash.scala 38:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[hash.scala 38:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[hash.scala 38:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[hash.scala 38:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[hash.scala 38:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[hash.scala 38:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[hash.scala 38:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[hash.scala 38:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[hash.scala 38:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[hash.scala 38:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[hash.scala 38:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[hash.scala 38:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[hash.scala 38:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[hash.scala 38:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[hash.scala 38:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[hash.scala 38:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[hash.scala 38:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[hash.scala 38:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[hash.scala 38:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[hash.scala 38:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[hash.scala 38:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[hash.scala 38:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[hash.scala 38:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[hash.scala 38:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[hash.scala 38:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[hash.scala 38:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[hash.scala 38:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[hash.scala 38:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[hash.scala 38:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[hash.scala 38:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[hash.scala 38:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[hash.scala 38:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[hash.scala 38:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[hash.scala 38:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[hash.scala 38:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[hash.scala 38:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[hash.scala 38:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[hash.scala 38:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[hash.scala 38:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[hash.scala 38:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[hash.scala 38:13]
    key <= io_key_in; // @[hash.scala 42:13]
    sum <= io_sum_in; // @[hash.scala 46:13]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  phv_next_config_id = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_117[0:0];
  _RAND_118 = {2{`RANDOM}};
  key = _RAND_118[63:0];
  _RAND_119 = {1{`RANDOM}};
  sum = _RAND_119[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HashSumLevel_2(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input  [63:0] io_key_in,
  output [63:0] io_key_out,
  input  [15:0] io_sum_in,
  output [15:0] io_sum_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [31:0] _RAND_119;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[hash.scala 37:22]
  reg [7:0] phv_data_1; // @[hash.scala 37:22]
  reg [7:0] phv_data_2; // @[hash.scala 37:22]
  reg [7:0] phv_data_3; // @[hash.scala 37:22]
  reg [7:0] phv_data_4; // @[hash.scala 37:22]
  reg [7:0] phv_data_5; // @[hash.scala 37:22]
  reg [7:0] phv_data_6; // @[hash.scala 37:22]
  reg [7:0] phv_data_7; // @[hash.scala 37:22]
  reg [7:0] phv_data_8; // @[hash.scala 37:22]
  reg [7:0] phv_data_9; // @[hash.scala 37:22]
  reg [7:0] phv_data_10; // @[hash.scala 37:22]
  reg [7:0] phv_data_11; // @[hash.scala 37:22]
  reg [7:0] phv_data_12; // @[hash.scala 37:22]
  reg [7:0] phv_data_13; // @[hash.scala 37:22]
  reg [7:0] phv_data_14; // @[hash.scala 37:22]
  reg [7:0] phv_data_15; // @[hash.scala 37:22]
  reg [7:0] phv_data_16; // @[hash.scala 37:22]
  reg [7:0] phv_data_17; // @[hash.scala 37:22]
  reg [7:0] phv_data_18; // @[hash.scala 37:22]
  reg [7:0] phv_data_19; // @[hash.scala 37:22]
  reg [7:0] phv_data_20; // @[hash.scala 37:22]
  reg [7:0] phv_data_21; // @[hash.scala 37:22]
  reg [7:0] phv_data_22; // @[hash.scala 37:22]
  reg [7:0] phv_data_23; // @[hash.scala 37:22]
  reg [7:0] phv_data_24; // @[hash.scala 37:22]
  reg [7:0] phv_data_25; // @[hash.scala 37:22]
  reg [7:0] phv_data_26; // @[hash.scala 37:22]
  reg [7:0] phv_data_27; // @[hash.scala 37:22]
  reg [7:0] phv_data_28; // @[hash.scala 37:22]
  reg [7:0] phv_data_29; // @[hash.scala 37:22]
  reg [7:0] phv_data_30; // @[hash.scala 37:22]
  reg [7:0] phv_data_31; // @[hash.scala 37:22]
  reg [7:0] phv_data_32; // @[hash.scala 37:22]
  reg [7:0] phv_data_33; // @[hash.scala 37:22]
  reg [7:0] phv_data_34; // @[hash.scala 37:22]
  reg [7:0] phv_data_35; // @[hash.scala 37:22]
  reg [7:0] phv_data_36; // @[hash.scala 37:22]
  reg [7:0] phv_data_37; // @[hash.scala 37:22]
  reg [7:0] phv_data_38; // @[hash.scala 37:22]
  reg [7:0] phv_data_39; // @[hash.scala 37:22]
  reg [7:0] phv_data_40; // @[hash.scala 37:22]
  reg [7:0] phv_data_41; // @[hash.scala 37:22]
  reg [7:0] phv_data_42; // @[hash.scala 37:22]
  reg [7:0] phv_data_43; // @[hash.scala 37:22]
  reg [7:0] phv_data_44; // @[hash.scala 37:22]
  reg [7:0] phv_data_45; // @[hash.scala 37:22]
  reg [7:0] phv_data_46; // @[hash.scala 37:22]
  reg [7:0] phv_data_47; // @[hash.scala 37:22]
  reg [7:0] phv_data_48; // @[hash.scala 37:22]
  reg [7:0] phv_data_49; // @[hash.scala 37:22]
  reg [7:0] phv_data_50; // @[hash.scala 37:22]
  reg [7:0] phv_data_51; // @[hash.scala 37:22]
  reg [7:0] phv_data_52; // @[hash.scala 37:22]
  reg [7:0] phv_data_53; // @[hash.scala 37:22]
  reg [7:0] phv_data_54; // @[hash.scala 37:22]
  reg [7:0] phv_data_55; // @[hash.scala 37:22]
  reg [7:0] phv_data_56; // @[hash.scala 37:22]
  reg [7:0] phv_data_57; // @[hash.scala 37:22]
  reg [7:0] phv_data_58; // @[hash.scala 37:22]
  reg [7:0] phv_data_59; // @[hash.scala 37:22]
  reg [7:0] phv_data_60; // @[hash.scala 37:22]
  reg [7:0] phv_data_61; // @[hash.scala 37:22]
  reg [7:0] phv_data_62; // @[hash.scala 37:22]
  reg [7:0] phv_data_63; // @[hash.scala 37:22]
  reg [7:0] phv_data_64; // @[hash.scala 37:22]
  reg [7:0] phv_data_65; // @[hash.scala 37:22]
  reg [7:0] phv_data_66; // @[hash.scala 37:22]
  reg [7:0] phv_data_67; // @[hash.scala 37:22]
  reg [7:0] phv_data_68; // @[hash.scala 37:22]
  reg [7:0] phv_data_69; // @[hash.scala 37:22]
  reg [7:0] phv_data_70; // @[hash.scala 37:22]
  reg [7:0] phv_data_71; // @[hash.scala 37:22]
  reg [7:0] phv_data_72; // @[hash.scala 37:22]
  reg [7:0] phv_data_73; // @[hash.scala 37:22]
  reg [7:0] phv_data_74; // @[hash.scala 37:22]
  reg [7:0] phv_data_75; // @[hash.scala 37:22]
  reg [7:0] phv_data_76; // @[hash.scala 37:22]
  reg [7:0] phv_data_77; // @[hash.scala 37:22]
  reg [7:0] phv_data_78; // @[hash.scala 37:22]
  reg [7:0] phv_data_79; // @[hash.scala 37:22]
  reg [7:0] phv_data_80; // @[hash.scala 37:22]
  reg [7:0] phv_data_81; // @[hash.scala 37:22]
  reg [7:0] phv_data_82; // @[hash.scala 37:22]
  reg [7:0] phv_data_83; // @[hash.scala 37:22]
  reg [7:0] phv_data_84; // @[hash.scala 37:22]
  reg [7:0] phv_data_85; // @[hash.scala 37:22]
  reg [7:0] phv_data_86; // @[hash.scala 37:22]
  reg [7:0] phv_data_87; // @[hash.scala 37:22]
  reg [7:0] phv_data_88; // @[hash.scala 37:22]
  reg [7:0] phv_data_89; // @[hash.scala 37:22]
  reg [7:0] phv_data_90; // @[hash.scala 37:22]
  reg [7:0] phv_data_91; // @[hash.scala 37:22]
  reg [7:0] phv_data_92; // @[hash.scala 37:22]
  reg [7:0] phv_data_93; // @[hash.scala 37:22]
  reg [7:0] phv_data_94; // @[hash.scala 37:22]
  reg [7:0] phv_data_95; // @[hash.scala 37:22]
  reg [15:0] phv_header_0; // @[hash.scala 37:22]
  reg [15:0] phv_header_1; // @[hash.scala 37:22]
  reg [15:0] phv_header_2; // @[hash.scala 37:22]
  reg [15:0] phv_header_3; // @[hash.scala 37:22]
  reg [15:0] phv_header_4; // @[hash.scala 37:22]
  reg [15:0] phv_header_5; // @[hash.scala 37:22]
  reg [15:0] phv_header_6; // @[hash.scala 37:22]
  reg [15:0] phv_header_7; // @[hash.scala 37:22]
  reg [15:0] phv_header_8; // @[hash.scala 37:22]
  reg [15:0] phv_header_9; // @[hash.scala 37:22]
  reg [15:0] phv_header_10; // @[hash.scala 37:22]
  reg [15:0] phv_header_11; // @[hash.scala 37:22]
  reg [15:0] phv_header_12; // @[hash.scala 37:22]
  reg [15:0] phv_header_13; // @[hash.scala 37:22]
  reg [15:0] phv_header_14; // @[hash.scala 37:22]
  reg [15:0] phv_header_15; // @[hash.scala 37:22]
  reg [7:0] phv_parse_current_state; // @[hash.scala 37:22]
  reg [7:0] phv_parse_current_offset; // @[hash.scala 37:22]
  reg [15:0] phv_parse_transition_field; // @[hash.scala 37:22]
  reg [1:0] phv_next_processor_id; // @[hash.scala 37:22]
  reg  phv_next_config_id; // @[hash.scala 37:22]
  reg  phv_is_valid_processor; // @[hash.scala 37:22]
  reg [63:0] key; // @[hash.scala 41:22]
  reg [15:0] sum; // @[hash.scala 45:22]
  wire [15:0] _io_sum_out_T_2 = sum + key[63:48]; // @[hash.scala 49:31]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[hash.scala 39:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[hash.scala 39:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[hash.scala 39:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[hash.scala 39:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[hash.scala 39:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[hash.scala 39:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[hash.scala 39:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[hash.scala 39:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[hash.scala 39:25]
  assign io_key_out = key; // @[hash.scala 43:20]
  assign io_sum_out = phv_is_valid_processor ? _io_sum_out_T_2 : sum; // @[hash.scala 48:39 hash.scala 49:24 hash.scala 51:24]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[hash.scala 38:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[hash.scala 38:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[hash.scala 38:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[hash.scala 38:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[hash.scala 38:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[hash.scala 38:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[hash.scala 38:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[hash.scala 38:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[hash.scala 38:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[hash.scala 38:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[hash.scala 38:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[hash.scala 38:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[hash.scala 38:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[hash.scala 38:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[hash.scala 38:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[hash.scala 38:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[hash.scala 38:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[hash.scala 38:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[hash.scala 38:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[hash.scala 38:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[hash.scala 38:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[hash.scala 38:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[hash.scala 38:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[hash.scala 38:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[hash.scala 38:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[hash.scala 38:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[hash.scala 38:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[hash.scala 38:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[hash.scala 38:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[hash.scala 38:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[hash.scala 38:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[hash.scala 38:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[hash.scala 38:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[hash.scala 38:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[hash.scala 38:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[hash.scala 38:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[hash.scala 38:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[hash.scala 38:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[hash.scala 38:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[hash.scala 38:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[hash.scala 38:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[hash.scala 38:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[hash.scala 38:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[hash.scala 38:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[hash.scala 38:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[hash.scala 38:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[hash.scala 38:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[hash.scala 38:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[hash.scala 38:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[hash.scala 38:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[hash.scala 38:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[hash.scala 38:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[hash.scala 38:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[hash.scala 38:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[hash.scala 38:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[hash.scala 38:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[hash.scala 38:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[hash.scala 38:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[hash.scala 38:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[hash.scala 38:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[hash.scala 38:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[hash.scala 38:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[hash.scala 38:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[hash.scala 38:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[hash.scala 38:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[hash.scala 38:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[hash.scala 38:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[hash.scala 38:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[hash.scala 38:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[hash.scala 38:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[hash.scala 38:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[hash.scala 38:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[hash.scala 38:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[hash.scala 38:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[hash.scala 38:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[hash.scala 38:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[hash.scala 38:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[hash.scala 38:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[hash.scala 38:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[hash.scala 38:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[hash.scala 38:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[hash.scala 38:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[hash.scala 38:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[hash.scala 38:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[hash.scala 38:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[hash.scala 38:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[hash.scala 38:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[hash.scala 38:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[hash.scala 38:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[hash.scala 38:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[hash.scala 38:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[hash.scala 38:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[hash.scala 38:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[hash.scala 38:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[hash.scala 38:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[hash.scala 38:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[hash.scala 38:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[hash.scala 38:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[hash.scala 38:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[hash.scala 38:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[hash.scala 38:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[hash.scala 38:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[hash.scala 38:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[hash.scala 38:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[hash.scala 38:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[hash.scala 38:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[hash.scala 38:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[hash.scala 38:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[hash.scala 38:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[hash.scala 38:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[hash.scala 38:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[hash.scala 38:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[hash.scala 38:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[hash.scala 38:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[hash.scala 38:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[hash.scala 38:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[hash.scala 38:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[hash.scala 38:13]
    key <= io_key_in; // @[hash.scala 42:13]
    sum <= io_sum_in; // @[hash.scala 46:13]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  phv_next_config_id = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_117[0:0];
  _RAND_118 = {2{`RANDOM}};
  key = _RAND_118[63:0];
  _RAND_119 = {1{`RANDOM}};
  sum = _RAND_119[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HashReshapeLevel(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input  [2:0]  io_hash_depth_0,
  input  [2:0]  io_hash_depth_1,
  input  [63:0] io_key_in,
  output [63:0] io_key_out,
  input  [15:0] io_sum_in,
  output [15:0] io_sum_out,
  output [15:0] io_val_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[hash.scala 68:22]
  reg [7:0] phv_data_1; // @[hash.scala 68:22]
  reg [7:0] phv_data_2; // @[hash.scala 68:22]
  reg [7:0] phv_data_3; // @[hash.scala 68:22]
  reg [7:0] phv_data_4; // @[hash.scala 68:22]
  reg [7:0] phv_data_5; // @[hash.scala 68:22]
  reg [7:0] phv_data_6; // @[hash.scala 68:22]
  reg [7:0] phv_data_7; // @[hash.scala 68:22]
  reg [7:0] phv_data_8; // @[hash.scala 68:22]
  reg [7:0] phv_data_9; // @[hash.scala 68:22]
  reg [7:0] phv_data_10; // @[hash.scala 68:22]
  reg [7:0] phv_data_11; // @[hash.scala 68:22]
  reg [7:0] phv_data_12; // @[hash.scala 68:22]
  reg [7:0] phv_data_13; // @[hash.scala 68:22]
  reg [7:0] phv_data_14; // @[hash.scala 68:22]
  reg [7:0] phv_data_15; // @[hash.scala 68:22]
  reg [7:0] phv_data_16; // @[hash.scala 68:22]
  reg [7:0] phv_data_17; // @[hash.scala 68:22]
  reg [7:0] phv_data_18; // @[hash.scala 68:22]
  reg [7:0] phv_data_19; // @[hash.scala 68:22]
  reg [7:0] phv_data_20; // @[hash.scala 68:22]
  reg [7:0] phv_data_21; // @[hash.scala 68:22]
  reg [7:0] phv_data_22; // @[hash.scala 68:22]
  reg [7:0] phv_data_23; // @[hash.scala 68:22]
  reg [7:0] phv_data_24; // @[hash.scala 68:22]
  reg [7:0] phv_data_25; // @[hash.scala 68:22]
  reg [7:0] phv_data_26; // @[hash.scala 68:22]
  reg [7:0] phv_data_27; // @[hash.scala 68:22]
  reg [7:0] phv_data_28; // @[hash.scala 68:22]
  reg [7:0] phv_data_29; // @[hash.scala 68:22]
  reg [7:0] phv_data_30; // @[hash.scala 68:22]
  reg [7:0] phv_data_31; // @[hash.scala 68:22]
  reg [7:0] phv_data_32; // @[hash.scala 68:22]
  reg [7:0] phv_data_33; // @[hash.scala 68:22]
  reg [7:0] phv_data_34; // @[hash.scala 68:22]
  reg [7:0] phv_data_35; // @[hash.scala 68:22]
  reg [7:0] phv_data_36; // @[hash.scala 68:22]
  reg [7:0] phv_data_37; // @[hash.scala 68:22]
  reg [7:0] phv_data_38; // @[hash.scala 68:22]
  reg [7:0] phv_data_39; // @[hash.scala 68:22]
  reg [7:0] phv_data_40; // @[hash.scala 68:22]
  reg [7:0] phv_data_41; // @[hash.scala 68:22]
  reg [7:0] phv_data_42; // @[hash.scala 68:22]
  reg [7:0] phv_data_43; // @[hash.scala 68:22]
  reg [7:0] phv_data_44; // @[hash.scala 68:22]
  reg [7:0] phv_data_45; // @[hash.scala 68:22]
  reg [7:0] phv_data_46; // @[hash.scala 68:22]
  reg [7:0] phv_data_47; // @[hash.scala 68:22]
  reg [7:0] phv_data_48; // @[hash.scala 68:22]
  reg [7:0] phv_data_49; // @[hash.scala 68:22]
  reg [7:0] phv_data_50; // @[hash.scala 68:22]
  reg [7:0] phv_data_51; // @[hash.scala 68:22]
  reg [7:0] phv_data_52; // @[hash.scala 68:22]
  reg [7:0] phv_data_53; // @[hash.scala 68:22]
  reg [7:0] phv_data_54; // @[hash.scala 68:22]
  reg [7:0] phv_data_55; // @[hash.scala 68:22]
  reg [7:0] phv_data_56; // @[hash.scala 68:22]
  reg [7:0] phv_data_57; // @[hash.scala 68:22]
  reg [7:0] phv_data_58; // @[hash.scala 68:22]
  reg [7:0] phv_data_59; // @[hash.scala 68:22]
  reg [7:0] phv_data_60; // @[hash.scala 68:22]
  reg [7:0] phv_data_61; // @[hash.scala 68:22]
  reg [7:0] phv_data_62; // @[hash.scala 68:22]
  reg [7:0] phv_data_63; // @[hash.scala 68:22]
  reg [7:0] phv_data_64; // @[hash.scala 68:22]
  reg [7:0] phv_data_65; // @[hash.scala 68:22]
  reg [7:0] phv_data_66; // @[hash.scala 68:22]
  reg [7:0] phv_data_67; // @[hash.scala 68:22]
  reg [7:0] phv_data_68; // @[hash.scala 68:22]
  reg [7:0] phv_data_69; // @[hash.scala 68:22]
  reg [7:0] phv_data_70; // @[hash.scala 68:22]
  reg [7:0] phv_data_71; // @[hash.scala 68:22]
  reg [7:0] phv_data_72; // @[hash.scala 68:22]
  reg [7:0] phv_data_73; // @[hash.scala 68:22]
  reg [7:0] phv_data_74; // @[hash.scala 68:22]
  reg [7:0] phv_data_75; // @[hash.scala 68:22]
  reg [7:0] phv_data_76; // @[hash.scala 68:22]
  reg [7:0] phv_data_77; // @[hash.scala 68:22]
  reg [7:0] phv_data_78; // @[hash.scala 68:22]
  reg [7:0] phv_data_79; // @[hash.scala 68:22]
  reg [7:0] phv_data_80; // @[hash.scala 68:22]
  reg [7:0] phv_data_81; // @[hash.scala 68:22]
  reg [7:0] phv_data_82; // @[hash.scala 68:22]
  reg [7:0] phv_data_83; // @[hash.scala 68:22]
  reg [7:0] phv_data_84; // @[hash.scala 68:22]
  reg [7:0] phv_data_85; // @[hash.scala 68:22]
  reg [7:0] phv_data_86; // @[hash.scala 68:22]
  reg [7:0] phv_data_87; // @[hash.scala 68:22]
  reg [7:0] phv_data_88; // @[hash.scala 68:22]
  reg [7:0] phv_data_89; // @[hash.scala 68:22]
  reg [7:0] phv_data_90; // @[hash.scala 68:22]
  reg [7:0] phv_data_91; // @[hash.scala 68:22]
  reg [7:0] phv_data_92; // @[hash.scala 68:22]
  reg [7:0] phv_data_93; // @[hash.scala 68:22]
  reg [7:0] phv_data_94; // @[hash.scala 68:22]
  reg [7:0] phv_data_95; // @[hash.scala 68:22]
  reg [15:0] phv_header_0; // @[hash.scala 68:22]
  reg [15:0] phv_header_1; // @[hash.scala 68:22]
  reg [15:0] phv_header_2; // @[hash.scala 68:22]
  reg [15:0] phv_header_3; // @[hash.scala 68:22]
  reg [15:0] phv_header_4; // @[hash.scala 68:22]
  reg [15:0] phv_header_5; // @[hash.scala 68:22]
  reg [15:0] phv_header_6; // @[hash.scala 68:22]
  reg [15:0] phv_header_7; // @[hash.scala 68:22]
  reg [15:0] phv_header_8; // @[hash.scala 68:22]
  reg [15:0] phv_header_9; // @[hash.scala 68:22]
  reg [15:0] phv_header_10; // @[hash.scala 68:22]
  reg [15:0] phv_header_11; // @[hash.scala 68:22]
  reg [15:0] phv_header_12; // @[hash.scala 68:22]
  reg [15:0] phv_header_13; // @[hash.scala 68:22]
  reg [15:0] phv_header_14; // @[hash.scala 68:22]
  reg [15:0] phv_header_15; // @[hash.scala 68:22]
  reg [7:0] phv_parse_current_state; // @[hash.scala 68:22]
  reg [7:0] phv_parse_current_offset; // @[hash.scala 68:22]
  reg [15:0] phv_parse_transition_field; // @[hash.scala 68:22]
  reg [1:0] phv_next_processor_id; // @[hash.scala 68:22]
  reg  phv_next_config_id; // @[hash.scala 68:22]
  reg  phv_is_valid_processor; // @[hash.scala 68:22]
  reg [63:0] key; // @[hash.scala 72:22]
  reg [15:0] sum; // @[hash.scala 76:22]
  reg [2:0] hash_depth; // @[hash.scala 80:29]
  wire [16:0] _io_val_out_T_1 = {{1'd0}, sum}; // @[hash.scala 90:44]
  wire [15:0] _GEN_2 = hash_depth[0] ? _io_val_out_T_1[15:0] : 16'h0; // @[hash.scala 89:42 hash.scala 90:32 hash.scala 92:32]
  wire [15:0] _GEN_3 = hash_depth == 3'h0 ? sum : _GEN_2; // @[hash.scala 86:71 hash.scala 87:28]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[hash.scala 70:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[hash.scala 70:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[hash.scala 70:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[hash.scala 70:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[hash.scala 70:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[hash.scala 70:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[hash.scala 70:25]
  assign io_key_out = key; // @[hash.scala 74:20]
  assign io_sum_out = sum; // @[hash.scala 78:20]
  assign io_val_out = phv_is_valid_processor ? _GEN_3 : 16'h0; // @[hash.scala 85:39 hash.scala 96:24]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[hash.scala 69:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[hash.scala 69:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[hash.scala 69:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[hash.scala 69:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[hash.scala 69:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[hash.scala 69:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[hash.scala 69:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[hash.scala 69:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[hash.scala 69:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[hash.scala 69:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[hash.scala 69:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[hash.scala 69:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[hash.scala 69:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[hash.scala 69:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[hash.scala 69:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[hash.scala 69:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[hash.scala 69:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[hash.scala 69:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[hash.scala 69:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[hash.scala 69:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[hash.scala 69:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[hash.scala 69:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[hash.scala 69:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[hash.scala 69:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[hash.scala 69:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[hash.scala 69:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[hash.scala 69:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[hash.scala 69:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[hash.scala 69:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[hash.scala 69:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[hash.scala 69:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[hash.scala 69:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[hash.scala 69:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[hash.scala 69:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[hash.scala 69:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[hash.scala 69:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[hash.scala 69:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[hash.scala 69:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[hash.scala 69:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[hash.scala 69:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[hash.scala 69:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[hash.scala 69:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[hash.scala 69:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[hash.scala 69:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[hash.scala 69:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[hash.scala 69:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[hash.scala 69:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[hash.scala 69:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[hash.scala 69:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[hash.scala 69:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[hash.scala 69:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[hash.scala 69:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[hash.scala 69:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[hash.scala 69:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[hash.scala 69:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[hash.scala 69:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[hash.scala 69:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[hash.scala 69:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[hash.scala 69:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[hash.scala 69:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[hash.scala 69:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[hash.scala 69:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[hash.scala 69:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[hash.scala 69:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[hash.scala 69:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[hash.scala 69:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[hash.scala 69:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[hash.scala 69:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[hash.scala 69:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[hash.scala 69:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[hash.scala 69:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[hash.scala 69:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[hash.scala 69:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[hash.scala 69:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[hash.scala 69:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[hash.scala 69:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[hash.scala 69:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[hash.scala 69:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[hash.scala 69:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[hash.scala 69:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[hash.scala 69:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[hash.scala 69:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[hash.scala 69:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[hash.scala 69:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[hash.scala 69:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[hash.scala 69:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[hash.scala 69:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[hash.scala 69:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[hash.scala 69:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[hash.scala 69:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[hash.scala 69:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[hash.scala 69:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[hash.scala 69:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[hash.scala 69:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[hash.scala 69:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[hash.scala 69:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[hash.scala 69:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[hash.scala 69:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[hash.scala 69:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[hash.scala 69:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[hash.scala 69:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[hash.scala 69:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[hash.scala 69:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[hash.scala 69:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[hash.scala 69:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[hash.scala 69:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[hash.scala 69:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[hash.scala 69:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[hash.scala 69:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[hash.scala 69:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[hash.scala 69:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[hash.scala 69:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[hash.scala 69:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[hash.scala 69:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[hash.scala 69:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[hash.scala 69:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[hash.scala 69:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[hash.scala 69:13]
    key <= io_key_in; // @[hash.scala 73:13]
    sum <= io_sum_in; // @[hash.scala 77:13]
    if (io_pipe_phv_in_next_config_id) begin // @[hash.scala 81:20]
      hash_depth <= io_hash_depth_1; // @[hash.scala 81:20]
    end else begin
      hash_depth <= io_hash_depth_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  phv_next_config_id = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_117[0:0];
  _RAND_118 = {2{`RANDOM}};
  key = _RAND_118[63:0];
  _RAND_119 = {1{`RANDOM}};
  sum = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  hash_depth = _RAND_120[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HashReshapeLevel_1(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input  [2:0]  io_hash_depth_0,
  input  [2:0]  io_hash_depth_1,
  input  [63:0] io_key_in,
  output [63:0] io_key_out,
  input  [15:0] io_sum_in,
  output [15:0] io_sum_out,
  input  [15:0] io_val_in,
  output [15:0] io_val_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[hash.scala 68:22]
  reg [7:0] phv_data_1; // @[hash.scala 68:22]
  reg [7:0] phv_data_2; // @[hash.scala 68:22]
  reg [7:0] phv_data_3; // @[hash.scala 68:22]
  reg [7:0] phv_data_4; // @[hash.scala 68:22]
  reg [7:0] phv_data_5; // @[hash.scala 68:22]
  reg [7:0] phv_data_6; // @[hash.scala 68:22]
  reg [7:0] phv_data_7; // @[hash.scala 68:22]
  reg [7:0] phv_data_8; // @[hash.scala 68:22]
  reg [7:0] phv_data_9; // @[hash.scala 68:22]
  reg [7:0] phv_data_10; // @[hash.scala 68:22]
  reg [7:0] phv_data_11; // @[hash.scala 68:22]
  reg [7:0] phv_data_12; // @[hash.scala 68:22]
  reg [7:0] phv_data_13; // @[hash.scala 68:22]
  reg [7:0] phv_data_14; // @[hash.scala 68:22]
  reg [7:0] phv_data_15; // @[hash.scala 68:22]
  reg [7:0] phv_data_16; // @[hash.scala 68:22]
  reg [7:0] phv_data_17; // @[hash.scala 68:22]
  reg [7:0] phv_data_18; // @[hash.scala 68:22]
  reg [7:0] phv_data_19; // @[hash.scala 68:22]
  reg [7:0] phv_data_20; // @[hash.scala 68:22]
  reg [7:0] phv_data_21; // @[hash.scala 68:22]
  reg [7:0] phv_data_22; // @[hash.scala 68:22]
  reg [7:0] phv_data_23; // @[hash.scala 68:22]
  reg [7:0] phv_data_24; // @[hash.scala 68:22]
  reg [7:0] phv_data_25; // @[hash.scala 68:22]
  reg [7:0] phv_data_26; // @[hash.scala 68:22]
  reg [7:0] phv_data_27; // @[hash.scala 68:22]
  reg [7:0] phv_data_28; // @[hash.scala 68:22]
  reg [7:0] phv_data_29; // @[hash.scala 68:22]
  reg [7:0] phv_data_30; // @[hash.scala 68:22]
  reg [7:0] phv_data_31; // @[hash.scala 68:22]
  reg [7:0] phv_data_32; // @[hash.scala 68:22]
  reg [7:0] phv_data_33; // @[hash.scala 68:22]
  reg [7:0] phv_data_34; // @[hash.scala 68:22]
  reg [7:0] phv_data_35; // @[hash.scala 68:22]
  reg [7:0] phv_data_36; // @[hash.scala 68:22]
  reg [7:0] phv_data_37; // @[hash.scala 68:22]
  reg [7:0] phv_data_38; // @[hash.scala 68:22]
  reg [7:0] phv_data_39; // @[hash.scala 68:22]
  reg [7:0] phv_data_40; // @[hash.scala 68:22]
  reg [7:0] phv_data_41; // @[hash.scala 68:22]
  reg [7:0] phv_data_42; // @[hash.scala 68:22]
  reg [7:0] phv_data_43; // @[hash.scala 68:22]
  reg [7:0] phv_data_44; // @[hash.scala 68:22]
  reg [7:0] phv_data_45; // @[hash.scala 68:22]
  reg [7:0] phv_data_46; // @[hash.scala 68:22]
  reg [7:0] phv_data_47; // @[hash.scala 68:22]
  reg [7:0] phv_data_48; // @[hash.scala 68:22]
  reg [7:0] phv_data_49; // @[hash.scala 68:22]
  reg [7:0] phv_data_50; // @[hash.scala 68:22]
  reg [7:0] phv_data_51; // @[hash.scala 68:22]
  reg [7:0] phv_data_52; // @[hash.scala 68:22]
  reg [7:0] phv_data_53; // @[hash.scala 68:22]
  reg [7:0] phv_data_54; // @[hash.scala 68:22]
  reg [7:0] phv_data_55; // @[hash.scala 68:22]
  reg [7:0] phv_data_56; // @[hash.scala 68:22]
  reg [7:0] phv_data_57; // @[hash.scala 68:22]
  reg [7:0] phv_data_58; // @[hash.scala 68:22]
  reg [7:0] phv_data_59; // @[hash.scala 68:22]
  reg [7:0] phv_data_60; // @[hash.scala 68:22]
  reg [7:0] phv_data_61; // @[hash.scala 68:22]
  reg [7:0] phv_data_62; // @[hash.scala 68:22]
  reg [7:0] phv_data_63; // @[hash.scala 68:22]
  reg [7:0] phv_data_64; // @[hash.scala 68:22]
  reg [7:0] phv_data_65; // @[hash.scala 68:22]
  reg [7:0] phv_data_66; // @[hash.scala 68:22]
  reg [7:0] phv_data_67; // @[hash.scala 68:22]
  reg [7:0] phv_data_68; // @[hash.scala 68:22]
  reg [7:0] phv_data_69; // @[hash.scala 68:22]
  reg [7:0] phv_data_70; // @[hash.scala 68:22]
  reg [7:0] phv_data_71; // @[hash.scala 68:22]
  reg [7:0] phv_data_72; // @[hash.scala 68:22]
  reg [7:0] phv_data_73; // @[hash.scala 68:22]
  reg [7:0] phv_data_74; // @[hash.scala 68:22]
  reg [7:0] phv_data_75; // @[hash.scala 68:22]
  reg [7:0] phv_data_76; // @[hash.scala 68:22]
  reg [7:0] phv_data_77; // @[hash.scala 68:22]
  reg [7:0] phv_data_78; // @[hash.scala 68:22]
  reg [7:0] phv_data_79; // @[hash.scala 68:22]
  reg [7:0] phv_data_80; // @[hash.scala 68:22]
  reg [7:0] phv_data_81; // @[hash.scala 68:22]
  reg [7:0] phv_data_82; // @[hash.scala 68:22]
  reg [7:0] phv_data_83; // @[hash.scala 68:22]
  reg [7:0] phv_data_84; // @[hash.scala 68:22]
  reg [7:0] phv_data_85; // @[hash.scala 68:22]
  reg [7:0] phv_data_86; // @[hash.scala 68:22]
  reg [7:0] phv_data_87; // @[hash.scala 68:22]
  reg [7:0] phv_data_88; // @[hash.scala 68:22]
  reg [7:0] phv_data_89; // @[hash.scala 68:22]
  reg [7:0] phv_data_90; // @[hash.scala 68:22]
  reg [7:0] phv_data_91; // @[hash.scala 68:22]
  reg [7:0] phv_data_92; // @[hash.scala 68:22]
  reg [7:0] phv_data_93; // @[hash.scala 68:22]
  reg [7:0] phv_data_94; // @[hash.scala 68:22]
  reg [7:0] phv_data_95; // @[hash.scala 68:22]
  reg [15:0] phv_header_0; // @[hash.scala 68:22]
  reg [15:0] phv_header_1; // @[hash.scala 68:22]
  reg [15:0] phv_header_2; // @[hash.scala 68:22]
  reg [15:0] phv_header_3; // @[hash.scala 68:22]
  reg [15:0] phv_header_4; // @[hash.scala 68:22]
  reg [15:0] phv_header_5; // @[hash.scala 68:22]
  reg [15:0] phv_header_6; // @[hash.scala 68:22]
  reg [15:0] phv_header_7; // @[hash.scala 68:22]
  reg [15:0] phv_header_8; // @[hash.scala 68:22]
  reg [15:0] phv_header_9; // @[hash.scala 68:22]
  reg [15:0] phv_header_10; // @[hash.scala 68:22]
  reg [15:0] phv_header_11; // @[hash.scala 68:22]
  reg [15:0] phv_header_12; // @[hash.scala 68:22]
  reg [15:0] phv_header_13; // @[hash.scala 68:22]
  reg [15:0] phv_header_14; // @[hash.scala 68:22]
  reg [15:0] phv_header_15; // @[hash.scala 68:22]
  reg [7:0] phv_parse_current_state; // @[hash.scala 68:22]
  reg [7:0] phv_parse_current_offset; // @[hash.scala 68:22]
  reg [15:0] phv_parse_transition_field; // @[hash.scala 68:22]
  reg [1:0] phv_next_processor_id; // @[hash.scala 68:22]
  reg  phv_next_config_id; // @[hash.scala 68:22]
  reg  phv_is_valid_processor; // @[hash.scala 68:22]
  reg [63:0] key; // @[hash.scala 72:22]
  reg [15:0] sum; // @[hash.scala 76:22]
  reg [2:0] hash_depth; // @[hash.scala 80:29]
  reg [15:0] hash_val; // @[hash.scala 82:27]
  wire [15:0] _GEN_5 = {{1'd0}, sum[14:0]}; // @[hash.scala 90:44]
  wire [15:0] _io_val_out_T_2 = hash_val + _GEN_5; // @[hash.scala 90:44]
  wire [15:0] _GEN_2 = hash_depth[1] ? _io_val_out_T_2 : hash_val; // @[hash.scala 89:42 hash.scala 90:32 hash.scala 92:32]
  wire [15:0] _GEN_3 = hash_depth == 3'h0 ? sum : _GEN_2; // @[hash.scala 86:71 hash.scala 87:28]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[hash.scala 70:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[hash.scala 70:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[hash.scala 70:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[hash.scala 70:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[hash.scala 70:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[hash.scala 70:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[hash.scala 70:25]
  assign io_key_out = key; // @[hash.scala 74:20]
  assign io_sum_out = sum; // @[hash.scala 78:20]
  assign io_val_out = phv_is_valid_processor ? _GEN_3 : hash_val; // @[hash.scala 85:39 hash.scala 96:24]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[hash.scala 69:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[hash.scala 69:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[hash.scala 69:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[hash.scala 69:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[hash.scala 69:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[hash.scala 69:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[hash.scala 69:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[hash.scala 69:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[hash.scala 69:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[hash.scala 69:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[hash.scala 69:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[hash.scala 69:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[hash.scala 69:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[hash.scala 69:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[hash.scala 69:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[hash.scala 69:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[hash.scala 69:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[hash.scala 69:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[hash.scala 69:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[hash.scala 69:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[hash.scala 69:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[hash.scala 69:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[hash.scala 69:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[hash.scala 69:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[hash.scala 69:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[hash.scala 69:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[hash.scala 69:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[hash.scala 69:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[hash.scala 69:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[hash.scala 69:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[hash.scala 69:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[hash.scala 69:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[hash.scala 69:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[hash.scala 69:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[hash.scala 69:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[hash.scala 69:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[hash.scala 69:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[hash.scala 69:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[hash.scala 69:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[hash.scala 69:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[hash.scala 69:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[hash.scala 69:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[hash.scala 69:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[hash.scala 69:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[hash.scala 69:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[hash.scala 69:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[hash.scala 69:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[hash.scala 69:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[hash.scala 69:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[hash.scala 69:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[hash.scala 69:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[hash.scala 69:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[hash.scala 69:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[hash.scala 69:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[hash.scala 69:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[hash.scala 69:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[hash.scala 69:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[hash.scala 69:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[hash.scala 69:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[hash.scala 69:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[hash.scala 69:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[hash.scala 69:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[hash.scala 69:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[hash.scala 69:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[hash.scala 69:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[hash.scala 69:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[hash.scala 69:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[hash.scala 69:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[hash.scala 69:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[hash.scala 69:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[hash.scala 69:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[hash.scala 69:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[hash.scala 69:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[hash.scala 69:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[hash.scala 69:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[hash.scala 69:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[hash.scala 69:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[hash.scala 69:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[hash.scala 69:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[hash.scala 69:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[hash.scala 69:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[hash.scala 69:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[hash.scala 69:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[hash.scala 69:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[hash.scala 69:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[hash.scala 69:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[hash.scala 69:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[hash.scala 69:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[hash.scala 69:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[hash.scala 69:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[hash.scala 69:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[hash.scala 69:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[hash.scala 69:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[hash.scala 69:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[hash.scala 69:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[hash.scala 69:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[hash.scala 69:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[hash.scala 69:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[hash.scala 69:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[hash.scala 69:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[hash.scala 69:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[hash.scala 69:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[hash.scala 69:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[hash.scala 69:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[hash.scala 69:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[hash.scala 69:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[hash.scala 69:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[hash.scala 69:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[hash.scala 69:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[hash.scala 69:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[hash.scala 69:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[hash.scala 69:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[hash.scala 69:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[hash.scala 69:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[hash.scala 69:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[hash.scala 69:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[hash.scala 69:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[hash.scala 69:13]
    key <= io_key_in; // @[hash.scala 73:13]
    sum <= io_sum_in; // @[hash.scala 77:13]
    if (io_pipe_phv_in_next_config_id) begin // @[hash.scala 81:20]
      hash_depth <= io_hash_depth_1; // @[hash.scala 81:20]
    end else begin
      hash_depth <= io_hash_depth_0;
    end
    hash_val <= io_val_in; // @[hash.scala 83:18]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  phv_next_config_id = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_117[0:0];
  _RAND_118 = {2{`RANDOM}};
  key = _RAND_118[63:0];
  _RAND_119 = {1{`RANDOM}};
  sum = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  hash_depth = _RAND_120[2:0];
  _RAND_121 = {1{`RANDOM}};
  hash_val = _RAND_121[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HashReshapeLevel_2(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input  [2:0]  io_hash_depth_0,
  input  [2:0]  io_hash_depth_1,
  input  [63:0] io_key_in,
  output [63:0] io_key_out,
  input  [15:0] io_sum_in,
  output [15:0] io_sum_out,
  input  [15:0] io_val_in,
  output [15:0] io_val_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[hash.scala 68:22]
  reg [7:0] phv_data_1; // @[hash.scala 68:22]
  reg [7:0] phv_data_2; // @[hash.scala 68:22]
  reg [7:0] phv_data_3; // @[hash.scala 68:22]
  reg [7:0] phv_data_4; // @[hash.scala 68:22]
  reg [7:0] phv_data_5; // @[hash.scala 68:22]
  reg [7:0] phv_data_6; // @[hash.scala 68:22]
  reg [7:0] phv_data_7; // @[hash.scala 68:22]
  reg [7:0] phv_data_8; // @[hash.scala 68:22]
  reg [7:0] phv_data_9; // @[hash.scala 68:22]
  reg [7:0] phv_data_10; // @[hash.scala 68:22]
  reg [7:0] phv_data_11; // @[hash.scala 68:22]
  reg [7:0] phv_data_12; // @[hash.scala 68:22]
  reg [7:0] phv_data_13; // @[hash.scala 68:22]
  reg [7:0] phv_data_14; // @[hash.scala 68:22]
  reg [7:0] phv_data_15; // @[hash.scala 68:22]
  reg [7:0] phv_data_16; // @[hash.scala 68:22]
  reg [7:0] phv_data_17; // @[hash.scala 68:22]
  reg [7:0] phv_data_18; // @[hash.scala 68:22]
  reg [7:0] phv_data_19; // @[hash.scala 68:22]
  reg [7:0] phv_data_20; // @[hash.scala 68:22]
  reg [7:0] phv_data_21; // @[hash.scala 68:22]
  reg [7:0] phv_data_22; // @[hash.scala 68:22]
  reg [7:0] phv_data_23; // @[hash.scala 68:22]
  reg [7:0] phv_data_24; // @[hash.scala 68:22]
  reg [7:0] phv_data_25; // @[hash.scala 68:22]
  reg [7:0] phv_data_26; // @[hash.scala 68:22]
  reg [7:0] phv_data_27; // @[hash.scala 68:22]
  reg [7:0] phv_data_28; // @[hash.scala 68:22]
  reg [7:0] phv_data_29; // @[hash.scala 68:22]
  reg [7:0] phv_data_30; // @[hash.scala 68:22]
  reg [7:0] phv_data_31; // @[hash.scala 68:22]
  reg [7:0] phv_data_32; // @[hash.scala 68:22]
  reg [7:0] phv_data_33; // @[hash.scala 68:22]
  reg [7:0] phv_data_34; // @[hash.scala 68:22]
  reg [7:0] phv_data_35; // @[hash.scala 68:22]
  reg [7:0] phv_data_36; // @[hash.scala 68:22]
  reg [7:0] phv_data_37; // @[hash.scala 68:22]
  reg [7:0] phv_data_38; // @[hash.scala 68:22]
  reg [7:0] phv_data_39; // @[hash.scala 68:22]
  reg [7:0] phv_data_40; // @[hash.scala 68:22]
  reg [7:0] phv_data_41; // @[hash.scala 68:22]
  reg [7:0] phv_data_42; // @[hash.scala 68:22]
  reg [7:0] phv_data_43; // @[hash.scala 68:22]
  reg [7:0] phv_data_44; // @[hash.scala 68:22]
  reg [7:0] phv_data_45; // @[hash.scala 68:22]
  reg [7:0] phv_data_46; // @[hash.scala 68:22]
  reg [7:0] phv_data_47; // @[hash.scala 68:22]
  reg [7:0] phv_data_48; // @[hash.scala 68:22]
  reg [7:0] phv_data_49; // @[hash.scala 68:22]
  reg [7:0] phv_data_50; // @[hash.scala 68:22]
  reg [7:0] phv_data_51; // @[hash.scala 68:22]
  reg [7:0] phv_data_52; // @[hash.scala 68:22]
  reg [7:0] phv_data_53; // @[hash.scala 68:22]
  reg [7:0] phv_data_54; // @[hash.scala 68:22]
  reg [7:0] phv_data_55; // @[hash.scala 68:22]
  reg [7:0] phv_data_56; // @[hash.scala 68:22]
  reg [7:0] phv_data_57; // @[hash.scala 68:22]
  reg [7:0] phv_data_58; // @[hash.scala 68:22]
  reg [7:0] phv_data_59; // @[hash.scala 68:22]
  reg [7:0] phv_data_60; // @[hash.scala 68:22]
  reg [7:0] phv_data_61; // @[hash.scala 68:22]
  reg [7:0] phv_data_62; // @[hash.scala 68:22]
  reg [7:0] phv_data_63; // @[hash.scala 68:22]
  reg [7:0] phv_data_64; // @[hash.scala 68:22]
  reg [7:0] phv_data_65; // @[hash.scala 68:22]
  reg [7:0] phv_data_66; // @[hash.scala 68:22]
  reg [7:0] phv_data_67; // @[hash.scala 68:22]
  reg [7:0] phv_data_68; // @[hash.scala 68:22]
  reg [7:0] phv_data_69; // @[hash.scala 68:22]
  reg [7:0] phv_data_70; // @[hash.scala 68:22]
  reg [7:0] phv_data_71; // @[hash.scala 68:22]
  reg [7:0] phv_data_72; // @[hash.scala 68:22]
  reg [7:0] phv_data_73; // @[hash.scala 68:22]
  reg [7:0] phv_data_74; // @[hash.scala 68:22]
  reg [7:0] phv_data_75; // @[hash.scala 68:22]
  reg [7:0] phv_data_76; // @[hash.scala 68:22]
  reg [7:0] phv_data_77; // @[hash.scala 68:22]
  reg [7:0] phv_data_78; // @[hash.scala 68:22]
  reg [7:0] phv_data_79; // @[hash.scala 68:22]
  reg [7:0] phv_data_80; // @[hash.scala 68:22]
  reg [7:0] phv_data_81; // @[hash.scala 68:22]
  reg [7:0] phv_data_82; // @[hash.scala 68:22]
  reg [7:0] phv_data_83; // @[hash.scala 68:22]
  reg [7:0] phv_data_84; // @[hash.scala 68:22]
  reg [7:0] phv_data_85; // @[hash.scala 68:22]
  reg [7:0] phv_data_86; // @[hash.scala 68:22]
  reg [7:0] phv_data_87; // @[hash.scala 68:22]
  reg [7:0] phv_data_88; // @[hash.scala 68:22]
  reg [7:0] phv_data_89; // @[hash.scala 68:22]
  reg [7:0] phv_data_90; // @[hash.scala 68:22]
  reg [7:0] phv_data_91; // @[hash.scala 68:22]
  reg [7:0] phv_data_92; // @[hash.scala 68:22]
  reg [7:0] phv_data_93; // @[hash.scala 68:22]
  reg [7:0] phv_data_94; // @[hash.scala 68:22]
  reg [7:0] phv_data_95; // @[hash.scala 68:22]
  reg [15:0] phv_header_0; // @[hash.scala 68:22]
  reg [15:0] phv_header_1; // @[hash.scala 68:22]
  reg [15:0] phv_header_2; // @[hash.scala 68:22]
  reg [15:0] phv_header_3; // @[hash.scala 68:22]
  reg [15:0] phv_header_4; // @[hash.scala 68:22]
  reg [15:0] phv_header_5; // @[hash.scala 68:22]
  reg [15:0] phv_header_6; // @[hash.scala 68:22]
  reg [15:0] phv_header_7; // @[hash.scala 68:22]
  reg [15:0] phv_header_8; // @[hash.scala 68:22]
  reg [15:0] phv_header_9; // @[hash.scala 68:22]
  reg [15:0] phv_header_10; // @[hash.scala 68:22]
  reg [15:0] phv_header_11; // @[hash.scala 68:22]
  reg [15:0] phv_header_12; // @[hash.scala 68:22]
  reg [15:0] phv_header_13; // @[hash.scala 68:22]
  reg [15:0] phv_header_14; // @[hash.scala 68:22]
  reg [15:0] phv_header_15; // @[hash.scala 68:22]
  reg [7:0] phv_parse_current_state; // @[hash.scala 68:22]
  reg [7:0] phv_parse_current_offset; // @[hash.scala 68:22]
  reg [15:0] phv_parse_transition_field; // @[hash.scala 68:22]
  reg [1:0] phv_next_processor_id; // @[hash.scala 68:22]
  reg  phv_next_config_id; // @[hash.scala 68:22]
  reg  phv_is_valid_processor; // @[hash.scala 68:22]
  reg [63:0] key; // @[hash.scala 72:22]
  reg [15:0] sum; // @[hash.scala 76:22]
  reg [2:0] hash_depth; // @[hash.scala 80:29]
  reg [15:0] hash_val; // @[hash.scala 82:27]
  wire [15:0] _GEN_5 = {{2'd0}, sum[13:0]}; // @[hash.scala 90:44]
  wire [15:0] _io_val_out_T_2 = hash_val + _GEN_5; // @[hash.scala 90:44]
  wire [15:0] _GEN_2 = hash_depth[2] ? _io_val_out_T_2 : hash_val; // @[hash.scala 89:42 hash.scala 90:32 hash.scala 92:32]
  wire [15:0] _GEN_3 = hash_depth == 3'h0 ? sum : _GEN_2; // @[hash.scala 86:71 hash.scala 87:28]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[hash.scala 70:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[hash.scala 70:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[hash.scala 70:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[hash.scala 70:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[hash.scala 70:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[hash.scala 70:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[hash.scala 70:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[hash.scala 70:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[hash.scala 70:25]
  assign io_key_out = key; // @[hash.scala 74:20]
  assign io_sum_out = sum; // @[hash.scala 78:20]
  assign io_val_out = phv_is_valid_processor ? _GEN_3 : hash_val; // @[hash.scala 85:39 hash.scala 96:24]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[hash.scala 69:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[hash.scala 69:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[hash.scala 69:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[hash.scala 69:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[hash.scala 69:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[hash.scala 69:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[hash.scala 69:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[hash.scala 69:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[hash.scala 69:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[hash.scala 69:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[hash.scala 69:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[hash.scala 69:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[hash.scala 69:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[hash.scala 69:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[hash.scala 69:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[hash.scala 69:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[hash.scala 69:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[hash.scala 69:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[hash.scala 69:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[hash.scala 69:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[hash.scala 69:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[hash.scala 69:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[hash.scala 69:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[hash.scala 69:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[hash.scala 69:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[hash.scala 69:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[hash.scala 69:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[hash.scala 69:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[hash.scala 69:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[hash.scala 69:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[hash.scala 69:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[hash.scala 69:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[hash.scala 69:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[hash.scala 69:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[hash.scala 69:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[hash.scala 69:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[hash.scala 69:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[hash.scala 69:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[hash.scala 69:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[hash.scala 69:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[hash.scala 69:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[hash.scala 69:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[hash.scala 69:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[hash.scala 69:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[hash.scala 69:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[hash.scala 69:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[hash.scala 69:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[hash.scala 69:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[hash.scala 69:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[hash.scala 69:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[hash.scala 69:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[hash.scala 69:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[hash.scala 69:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[hash.scala 69:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[hash.scala 69:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[hash.scala 69:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[hash.scala 69:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[hash.scala 69:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[hash.scala 69:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[hash.scala 69:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[hash.scala 69:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[hash.scala 69:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[hash.scala 69:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[hash.scala 69:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[hash.scala 69:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[hash.scala 69:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[hash.scala 69:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[hash.scala 69:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[hash.scala 69:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[hash.scala 69:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[hash.scala 69:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[hash.scala 69:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[hash.scala 69:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[hash.scala 69:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[hash.scala 69:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[hash.scala 69:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[hash.scala 69:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[hash.scala 69:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[hash.scala 69:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[hash.scala 69:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[hash.scala 69:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[hash.scala 69:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[hash.scala 69:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[hash.scala 69:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[hash.scala 69:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[hash.scala 69:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[hash.scala 69:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[hash.scala 69:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[hash.scala 69:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[hash.scala 69:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[hash.scala 69:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[hash.scala 69:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[hash.scala 69:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[hash.scala 69:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[hash.scala 69:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[hash.scala 69:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[hash.scala 69:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[hash.scala 69:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[hash.scala 69:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[hash.scala 69:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[hash.scala 69:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[hash.scala 69:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[hash.scala 69:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[hash.scala 69:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[hash.scala 69:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[hash.scala 69:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[hash.scala 69:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[hash.scala 69:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[hash.scala 69:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[hash.scala 69:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[hash.scala 69:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[hash.scala 69:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[hash.scala 69:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[hash.scala 69:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[hash.scala 69:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[hash.scala 69:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[hash.scala 69:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[hash.scala 69:13]
    key <= io_key_in; // @[hash.scala 73:13]
    sum <= io_sum_in; // @[hash.scala 77:13]
    if (io_pipe_phv_in_next_config_id) begin // @[hash.scala 81:20]
      hash_depth <= io_hash_depth_1; // @[hash.scala 81:20]
    end else begin
      hash_depth <= io_hash_depth_0;
    end
    hash_val <= io_val_in; // @[hash.scala 83:18]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  phv_next_config_id = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_117[0:0];
  _RAND_118 = {2{`RANDOM}};
  key = _RAND_118[63:0];
  _RAND_119 = {1{`RANDOM}};
  sum = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  hash_depth = _RAND_120[2:0];
  _RAND_121 = {1{`RANDOM}};
  hash_val = _RAND_121[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Hash(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input         io_mod_hash_depth_mod,
  input         io_mod_config_id,
  input  [2:0]  io_mod_hash_depth,
  input  [63:0] io_key_in,
  output [63:0] io_key_out,
  output [7:0]  io_hash_val,
  output [2:0]  io_hash_val_cs
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  pipe1_clock; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_0; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_1; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_2; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_3; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_4; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_5; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_6; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_7; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_8; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_9; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_10; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_11; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_12; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_13; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_14; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_15; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_16; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_17; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_18; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_19; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_20; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_21; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_22; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_23; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_24; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_25; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_26; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_27; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_28; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_29; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_30; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_31; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_32; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_33; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_34; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_35; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_36; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_37; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_38; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_39; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_40; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_41; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_42; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_43; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_44; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_45; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_46; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_47; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_48; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_49; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_50; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_51; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_52; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_53; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_54; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_55; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_56; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_57; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_58; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_59; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_60; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_61; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_62; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_63; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_64; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_65; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_66; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_67; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_68; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_69; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_70; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_71; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_72; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_73; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_74; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_75; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_76; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_77; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_78; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_79; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_80; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_81; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_82; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_83; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_84; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_85; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_86; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_87; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_88; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_89; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_90; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_91; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_92; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_93; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_94; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_95; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_0; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_1; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_2; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_3; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_4; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_5; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_6; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_7; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_8; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_9; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_10; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_11; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_12; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_13; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_14; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_15; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_state; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_offset; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_parse_transition_field; // @[hash.scala 101:23]
  wire [1:0] pipe1_io_pipe_phv_in_next_processor_id; // @[hash.scala 101:23]
  wire  pipe1_io_pipe_phv_in_next_config_id; // @[hash.scala 101:23]
  wire  pipe1_io_pipe_phv_in_is_valid_processor; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_0; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_1; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_2; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_3; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_4; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_5; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_6; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_7; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_8; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_9; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_10; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_11; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_12; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_13; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_14; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_15; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_16; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_17; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_18; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_19; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_20; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_21; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_22; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_23; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_24; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_25; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_26; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_27; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_28; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_29; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_30; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_31; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_32; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_33; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_34; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_35; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_36; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_37; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_38; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_39; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_40; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_41; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_42; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_43; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_44; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_45; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_46; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_47; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_48; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_49; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_50; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_51; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_52; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_53; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_54; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_55; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_56; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_57; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_58; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_59; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_60; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_61; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_62; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_63; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_64; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_65; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_66; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_67; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_68; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_69; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_70; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_71; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_72; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_73; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_74; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_75; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_76; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_77; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_78; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_79; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_80; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_81; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_82; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_83; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_84; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_85; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_86; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_87; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_88; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_89; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_90; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_91; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_92; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_93; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_94; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_95; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_0; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_1; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_2; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_3; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_4; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_5; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_6; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_7; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_8; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_9; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_10; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_11; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_12; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_13; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_14; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_15; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_state; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_offset; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_parse_transition_field; // @[hash.scala 101:23]
  wire [1:0] pipe1_io_pipe_phv_out_next_processor_id; // @[hash.scala 101:23]
  wire  pipe1_io_pipe_phv_out_next_config_id; // @[hash.scala 101:23]
  wire  pipe1_io_pipe_phv_out_is_valid_processor; // @[hash.scala 101:23]
  wire [63:0] pipe1_io_key_in; // @[hash.scala 101:23]
  wire [63:0] pipe1_io_key_out; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_sum_in; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_sum_out; // @[hash.scala 101:23]
  wire  pipe2_clock; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_0; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_1; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_2; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_3; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_4; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_5; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_6; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_7; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_8; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_9; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_10; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_11; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_12; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_13; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_14; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_15; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_16; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_17; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_18; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_19; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_20; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_21; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_22; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_23; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_24; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_25; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_26; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_27; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_28; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_29; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_30; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_31; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_32; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_33; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_34; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_35; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_36; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_37; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_38; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_39; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_40; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_41; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_42; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_43; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_44; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_45; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_46; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_47; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_48; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_49; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_50; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_51; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_52; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_53; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_54; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_55; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_56; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_57; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_58; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_59; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_60; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_61; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_62; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_63; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_64; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_65; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_66; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_67; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_68; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_69; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_70; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_71; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_72; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_73; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_74; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_75; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_76; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_77; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_78; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_79; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_80; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_81; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_82; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_83; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_84; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_85; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_86; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_87; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_88; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_89; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_90; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_91; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_92; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_93; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_94; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_95; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_0; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_1; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_2; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_3; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_4; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_5; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_6; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_7; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_8; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_9; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_10; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_11; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_12; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_13; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_14; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_15; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_state; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_offset; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_parse_transition_field; // @[hash.scala 102:23]
  wire [1:0] pipe2_io_pipe_phv_in_next_processor_id; // @[hash.scala 102:23]
  wire  pipe2_io_pipe_phv_in_next_config_id; // @[hash.scala 102:23]
  wire  pipe2_io_pipe_phv_in_is_valid_processor; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_0; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_1; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_2; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_3; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_4; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_5; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_6; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_7; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_8; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_9; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_10; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_11; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_12; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_13; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_14; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_15; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_16; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_17; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_18; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_19; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_20; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_21; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_22; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_23; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_24; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_25; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_26; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_27; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_28; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_29; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_30; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_31; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_32; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_33; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_34; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_35; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_36; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_37; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_38; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_39; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_40; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_41; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_42; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_43; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_44; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_45; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_46; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_47; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_48; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_49; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_50; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_51; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_52; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_53; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_54; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_55; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_56; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_57; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_58; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_59; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_60; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_61; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_62; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_63; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_64; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_65; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_66; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_67; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_68; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_69; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_70; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_71; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_72; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_73; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_74; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_75; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_76; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_77; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_78; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_79; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_80; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_81; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_82; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_83; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_84; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_85; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_86; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_87; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_88; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_89; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_90; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_91; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_92; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_93; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_94; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_95; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_0; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_1; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_2; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_3; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_4; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_5; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_6; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_7; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_8; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_9; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_10; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_11; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_12; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_13; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_14; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_15; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_state; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_offset; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_parse_transition_field; // @[hash.scala 102:23]
  wire [1:0] pipe2_io_pipe_phv_out_next_processor_id; // @[hash.scala 102:23]
  wire  pipe2_io_pipe_phv_out_next_config_id; // @[hash.scala 102:23]
  wire  pipe2_io_pipe_phv_out_is_valid_processor; // @[hash.scala 102:23]
  wire [63:0] pipe2_io_key_in; // @[hash.scala 102:23]
  wire [63:0] pipe2_io_key_out; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_sum_in; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_sum_out; // @[hash.scala 102:23]
  wire  pipe3_clock; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_0; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_1; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_2; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_3; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_4; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_5; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_6; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_7; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_8; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_9; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_10; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_11; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_12; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_13; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_14; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_15; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_16; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_17; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_18; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_19; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_20; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_21; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_22; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_23; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_24; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_25; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_26; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_27; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_28; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_29; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_30; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_31; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_32; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_33; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_34; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_35; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_36; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_37; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_38; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_39; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_40; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_41; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_42; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_43; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_44; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_45; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_46; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_47; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_48; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_49; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_50; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_51; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_52; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_53; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_54; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_55; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_56; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_57; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_58; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_59; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_60; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_61; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_62; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_63; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_64; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_65; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_66; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_67; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_68; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_69; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_70; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_71; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_72; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_73; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_74; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_75; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_76; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_77; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_78; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_79; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_80; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_81; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_82; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_83; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_84; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_85; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_86; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_87; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_88; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_89; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_90; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_91; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_92; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_93; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_94; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_95; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_0; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_1; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_2; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_3; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_4; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_5; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_6; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_7; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_8; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_9; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_10; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_11; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_12; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_13; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_14; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_15; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_parse_current_state; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_parse_current_offset; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_parse_transition_field; // @[hash.scala 103:23]
  wire [1:0] pipe3_io_pipe_phv_in_next_processor_id; // @[hash.scala 103:23]
  wire  pipe3_io_pipe_phv_in_next_config_id; // @[hash.scala 103:23]
  wire  pipe3_io_pipe_phv_in_is_valid_processor; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_0; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_1; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_2; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_3; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_4; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_5; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_6; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_7; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_8; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_9; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_10; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_11; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_12; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_13; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_14; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_15; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_16; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_17; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_18; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_19; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_20; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_21; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_22; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_23; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_24; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_25; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_26; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_27; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_28; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_29; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_30; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_31; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_32; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_33; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_34; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_35; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_36; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_37; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_38; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_39; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_40; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_41; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_42; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_43; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_44; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_45; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_46; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_47; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_48; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_49; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_50; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_51; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_52; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_53; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_54; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_55; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_56; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_57; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_58; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_59; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_60; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_61; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_62; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_63; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_64; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_65; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_66; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_67; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_68; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_69; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_70; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_71; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_72; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_73; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_74; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_75; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_76; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_77; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_78; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_79; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_80; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_81; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_82; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_83; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_84; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_85; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_86; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_87; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_88; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_89; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_90; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_91; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_92; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_93; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_94; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_95; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_0; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_1; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_2; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_3; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_4; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_5; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_6; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_7; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_8; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_9; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_10; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_11; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_12; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_13; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_14; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_15; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_parse_current_state; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_parse_current_offset; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_parse_transition_field; // @[hash.scala 103:23]
  wire [1:0] pipe3_io_pipe_phv_out_next_processor_id; // @[hash.scala 103:23]
  wire  pipe3_io_pipe_phv_out_next_config_id; // @[hash.scala 103:23]
  wire  pipe3_io_pipe_phv_out_is_valid_processor; // @[hash.scala 103:23]
  wire [63:0] pipe3_io_key_in; // @[hash.scala 103:23]
  wire [63:0] pipe3_io_key_out; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_sum_in; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_sum_out; // @[hash.scala 103:23]
  wire  pipe4_clock; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_0; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_1; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_2; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_3; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_4; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_5; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_6; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_7; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_8; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_9; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_10; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_11; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_12; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_13; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_14; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_15; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_16; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_17; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_18; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_19; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_20; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_21; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_22; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_23; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_24; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_25; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_26; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_27; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_28; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_29; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_30; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_31; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_32; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_33; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_34; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_35; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_36; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_37; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_38; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_39; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_40; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_41; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_42; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_43; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_44; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_45; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_46; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_47; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_48; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_49; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_50; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_51; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_52; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_53; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_54; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_55; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_56; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_57; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_58; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_59; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_60; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_61; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_62; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_63; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_64; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_65; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_66; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_67; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_68; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_69; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_70; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_71; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_72; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_73; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_74; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_75; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_76; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_77; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_78; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_79; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_80; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_81; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_82; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_83; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_84; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_85; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_86; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_87; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_88; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_89; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_90; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_91; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_92; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_93; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_94; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_95; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_0; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_1; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_2; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_3; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_4; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_5; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_6; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_7; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_8; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_9; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_10; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_11; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_12; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_13; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_14; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_15; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_parse_current_state; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_parse_current_offset; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_parse_transition_field; // @[hash.scala 104:23]
  wire [1:0] pipe4_io_pipe_phv_in_next_processor_id; // @[hash.scala 104:23]
  wire  pipe4_io_pipe_phv_in_next_config_id; // @[hash.scala 104:23]
  wire  pipe4_io_pipe_phv_in_is_valid_processor; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_0; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_1; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_2; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_3; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_4; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_5; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_6; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_7; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_8; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_9; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_10; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_11; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_12; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_13; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_14; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_15; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_16; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_17; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_18; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_19; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_20; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_21; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_22; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_23; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_24; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_25; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_26; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_27; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_28; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_29; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_30; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_31; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_32; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_33; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_34; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_35; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_36; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_37; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_38; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_39; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_40; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_41; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_42; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_43; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_44; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_45; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_46; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_47; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_48; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_49; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_50; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_51; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_52; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_53; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_54; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_55; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_56; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_57; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_58; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_59; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_60; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_61; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_62; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_63; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_64; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_65; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_66; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_67; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_68; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_69; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_70; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_71; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_72; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_73; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_74; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_75; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_76; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_77; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_78; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_79; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_80; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_81; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_82; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_83; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_84; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_85; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_86; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_87; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_88; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_89; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_90; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_91; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_92; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_93; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_94; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_95; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_0; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_1; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_2; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_3; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_4; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_5; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_6; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_7; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_8; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_9; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_10; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_11; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_12; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_13; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_14; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_15; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_parse_current_state; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_parse_current_offset; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_parse_transition_field; // @[hash.scala 104:23]
  wire [1:0] pipe4_io_pipe_phv_out_next_processor_id; // @[hash.scala 104:23]
  wire  pipe4_io_pipe_phv_out_next_config_id; // @[hash.scala 104:23]
  wire  pipe4_io_pipe_phv_out_is_valid_processor; // @[hash.scala 104:23]
  wire [2:0] pipe4_io_hash_depth_0; // @[hash.scala 104:23]
  wire [2:0] pipe4_io_hash_depth_1; // @[hash.scala 104:23]
  wire [63:0] pipe4_io_key_in; // @[hash.scala 104:23]
  wire [63:0] pipe4_io_key_out; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_sum_in; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_sum_out; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_val_out; // @[hash.scala 104:23]
  wire  pipe5_clock; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_0; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_1; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_2; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_3; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_4; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_5; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_6; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_7; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_8; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_9; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_10; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_11; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_12; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_13; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_14; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_15; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_16; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_17; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_18; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_19; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_20; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_21; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_22; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_23; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_24; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_25; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_26; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_27; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_28; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_29; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_30; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_31; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_32; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_33; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_34; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_35; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_36; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_37; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_38; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_39; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_40; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_41; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_42; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_43; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_44; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_45; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_46; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_47; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_48; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_49; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_50; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_51; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_52; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_53; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_54; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_55; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_56; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_57; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_58; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_59; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_60; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_61; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_62; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_63; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_64; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_65; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_66; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_67; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_68; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_69; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_70; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_71; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_72; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_73; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_74; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_75; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_76; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_77; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_78; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_79; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_80; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_81; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_82; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_83; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_84; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_85; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_86; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_87; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_88; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_89; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_90; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_91; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_92; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_93; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_94; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_95; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_0; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_1; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_2; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_3; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_4; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_5; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_6; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_7; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_8; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_9; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_10; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_11; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_12; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_13; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_14; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_15; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_parse_current_state; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_parse_current_offset; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_parse_transition_field; // @[hash.scala 105:23]
  wire [1:0] pipe5_io_pipe_phv_in_next_processor_id; // @[hash.scala 105:23]
  wire  pipe5_io_pipe_phv_in_next_config_id; // @[hash.scala 105:23]
  wire  pipe5_io_pipe_phv_in_is_valid_processor; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_0; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_1; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_2; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_3; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_4; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_5; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_6; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_7; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_8; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_9; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_10; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_11; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_12; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_13; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_14; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_15; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_16; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_17; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_18; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_19; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_20; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_21; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_22; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_23; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_24; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_25; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_26; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_27; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_28; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_29; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_30; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_31; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_32; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_33; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_34; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_35; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_36; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_37; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_38; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_39; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_40; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_41; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_42; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_43; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_44; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_45; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_46; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_47; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_48; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_49; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_50; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_51; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_52; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_53; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_54; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_55; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_56; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_57; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_58; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_59; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_60; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_61; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_62; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_63; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_64; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_65; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_66; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_67; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_68; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_69; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_70; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_71; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_72; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_73; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_74; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_75; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_76; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_77; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_78; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_79; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_80; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_81; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_82; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_83; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_84; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_85; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_86; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_87; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_88; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_89; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_90; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_91; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_92; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_93; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_94; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_95; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_0; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_1; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_2; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_3; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_4; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_5; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_6; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_7; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_8; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_9; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_10; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_11; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_12; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_13; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_14; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_15; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_parse_current_state; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_parse_current_offset; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_parse_transition_field; // @[hash.scala 105:23]
  wire [1:0] pipe5_io_pipe_phv_out_next_processor_id; // @[hash.scala 105:23]
  wire  pipe5_io_pipe_phv_out_next_config_id; // @[hash.scala 105:23]
  wire  pipe5_io_pipe_phv_out_is_valid_processor; // @[hash.scala 105:23]
  wire [2:0] pipe5_io_hash_depth_0; // @[hash.scala 105:23]
  wire [2:0] pipe5_io_hash_depth_1; // @[hash.scala 105:23]
  wire [63:0] pipe5_io_key_in; // @[hash.scala 105:23]
  wire [63:0] pipe5_io_key_out; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_sum_in; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_sum_out; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_val_in; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_val_out; // @[hash.scala 105:23]
  wire  pipe6_clock; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_0; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_1; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_2; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_3; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_4; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_5; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_6; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_7; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_8; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_9; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_10; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_11; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_12; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_13; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_14; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_15; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_16; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_17; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_18; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_19; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_20; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_21; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_22; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_23; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_24; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_25; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_26; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_27; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_28; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_29; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_30; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_31; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_32; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_33; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_34; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_35; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_36; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_37; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_38; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_39; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_40; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_41; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_42; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_43; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_44; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_45; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_46; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_47; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_48; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_49; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_50; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_51; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_52; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_53; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_54; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_55; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_56; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_57; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_58; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_59; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_60; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_61; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_62; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_63; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_64; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_65; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_66; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_67; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_68; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_69; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_70; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_71; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_72; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_73; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_74; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_75; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_76; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_77; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_78; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_79; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_80; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_81; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_82; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_83; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_84; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_85; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_86; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_87; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_88; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_89; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_90; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_91; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_92; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_93; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_94; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_95; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_0; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_1; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_2; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_3; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_4; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_5; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_6; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_7; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_8; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_9; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_10; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_11; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_12; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_13; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_14; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_15; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_parse_current_state; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_parse_current_offset; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_parse_transition_field; // @[hash.scala 106:23]
  wire [1:0] pipe6_io_pipe_phv_in_next_processor_id; // @[hash.scala 106:23]
  wire  pipe6_io_pipe_phv_in_next_config_id; // @[hash.scala 106:23]
  wire  pipe6_io_pipe_phv_in_is_valid_processor; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_0; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_1; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_2; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_3; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_4; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_5; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_6; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_7; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_8; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_9; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_10; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_11; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_12; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_13; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_14; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_15; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_16; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_17; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_18; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_19; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_20; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_21; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_22; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_23; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_24; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_25; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_26; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_27; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_28; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_29; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_30; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_31; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_32; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_33; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_34; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_35; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_36; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_37; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_38; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_39; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_40; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_41; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_42; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_43; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_44; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_45; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_46; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_47; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_48; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_49; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_50; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_51; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_52; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_53; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_54; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_55; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_56; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_57; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_58; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_59; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_60; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_61; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_62; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_63; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_64; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_65; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_66; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_67; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_68; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_69; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_70; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_71; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_72; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_73; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_74; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_75; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_76; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_77; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_78; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_79; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_80; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_81; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_82; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_83; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_84; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_85; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_86; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_87; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_88; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_89; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_90; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_91; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_92; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_93; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_94; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_95; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_0; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_1; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_2; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_3; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_4; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_5; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_6; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_7; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_8; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_9; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_10; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_11; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_12; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_13; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_14; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_15; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_parse_current_state; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_parse_current_offset; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_parse_transition_field; // @[hash.scala 106:23]
  wire [1:0] pipe6_io_pipe_phv_out_next_processor_id; // @[hash.scala 106:23]
  wire  pipe6_io_pipe_phv_out_next_config_id; // @[hash.scala 106:23]
  wire  pipe6_io_pipe_phv_out_is_valid_processor; // @[hash.scala 106:23]
  wire [2:0] pipe6_io_hash_depth_0; // @[hash.scala 106:23]
  wire [2:0] pipe6_io_hash_depth_1; // @[hash.scala 106:23]
  wire [63:0] pipe6_io_key_in; // @[hash.scala 106:23]
  wire [63:0] pipe6_io_key_out; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_sum_in; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_sum_out; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_val_in; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_val_out; // @[hash.scala 106:23]
  reg [2:0] hash_depth_0; // @[hash.scala 18:26]
  reg [2:0] hash_depth_1; // @[hash.scala 18:26]
  HashSumLevel pipe1 ( // @[hash.scala 101:23]
    .clock(pipe1_clock),
    .io_pipe_phv_in_data_0(pipe1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe1_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe1_io_key_in),
    .io_key_out(pipe1_io_key_out),
    .io_sum_in(pipe1_io_sum_in),
    .io_sum_out(pipe1_io_sum_out)
  );
  HashSumLevel_1 pipe2 ( // @[hash.scala 102:23]
    .clock(pipe2_clock),
    .io_pipe_phv_in_data_0(pipe2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe2_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe2_io_key_in),
    .io_key_out(pipe2_io_key_out),
    .io_sum_in(pipe2_io_sum_in),
    .io_sum_out(pipe2_io_sum_out)
  );
  HashSumLevel_2 pipe3 ( // @[hash.scala 103:23]
    .clock(pipe3_clock),
    .io_pipe_phv_in_data_0(pipe3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe3_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe3_io_key_in),
    .io_key_out(pipe3_io_key_out),
    .io_sum_in(pipe3_io_sum_in),
    .io_sum_out(pipe3_io_sum_out)
  );
  HashReshapeLevel pipe4 ( // @[hash.scala 104:23]
    .clock(pipe4_clock),
    .io_pipe_phv_in_data_0(pipe4_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe4_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe4_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe4_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe4_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe4_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe4_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe4_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe4_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe4_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe4_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe4_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe4_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe4_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe4_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe4_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe4_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe4_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe4_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe4_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe4_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe4_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe4_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe4_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe4_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe4_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe4_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe4_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe4_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe4_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe4_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe4_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe4_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe4_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe4_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe4_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe4_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe4_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe4_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe4_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe4_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe4_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe4_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe4_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe4_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe4_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe4_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe4_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe4_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe4_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe4_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe4_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe4_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe4_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe4_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe4_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe4_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe4_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe4_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe4_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe4_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe4_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe4_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe4_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe4_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe4_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe4_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe4_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe4_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe4_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe4_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe4_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe4_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe4_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe4_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe4_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe4_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe4_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe4_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe4_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe4_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe4_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe4_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe4_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe4_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe4_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe4_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe4_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe4_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe4_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe4_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe4_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe4_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe4_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe4_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe4_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe4_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe4_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe4_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe4_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe4_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe4_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe4_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe4_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe4_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe4_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe4_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe4_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe4_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe4_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe4_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe4_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe4_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe4_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe4_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe4_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe4_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe4_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe4_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe4_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe4_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe4_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe4_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe4_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe4_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe4_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe4_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe4_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe4_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe4_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe4_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe4_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe4_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe4_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe4_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe4_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe4_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe4_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe4_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe4_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe4_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe4_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe4_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe4_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe4_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe4_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe4_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe4_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe4_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe4_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe4_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe4_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe4_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe4_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe4_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe4_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe4_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe4_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe4_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe4_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe4_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe4_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe4_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe4_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe4_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe4_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe4_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe4_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe4_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe4_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe4_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe4_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe4_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe4_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe4_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe4_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe4_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe4_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe4_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe4_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe4_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe4_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe4_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe4_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe4_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe4_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe4_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe4_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe4_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe4_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe4_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe4_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe4_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe4_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe4_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe4_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe4_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe4_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe4_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe4_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe4_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe4_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe4_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe4_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe4_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe4_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe4_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe4_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe4_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe4_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe4_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe4_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe4_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe4_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe4_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe4_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe4_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe4_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe4_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe4_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe4_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe4_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe4_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe4_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe4_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe4_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe4_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe4_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe4_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe4_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe4_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe4_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe4_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe4_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe4_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe4_io_pipe_phv_out_is_valid_processor),
    .io_hash_depth_0(pipe4_io_hash_depth_0),
    .io_hash_depth_1(pipe4_io_hash_depth_1),
    .io_key_in(pipe4_io_key_in),
    .io_key_out(pipe4_io_key_out),
    .io_sum_in(pipe4_io_sum_in),
    .io_sum_out(pipe4_io_sum_out),
    .io_val_out(pipe4_io_val_out)
  );
  HashReshapeLevel_1 pipe5 ( // @[hash.scala 105:23]
    .clock(pipe5_clock),
    .io_pipe_phv_in_data_0(pipe5_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe5_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe5_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe5_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe5_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe5_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe5_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe5_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe5_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe5_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe5_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe5_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe5_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe5_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe5_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe5_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe5_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe5_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe5_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe5_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe5_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe5_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe5_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe5_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe5_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe5_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe5_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe5_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe5_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe5_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe5_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe5_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe5_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe5_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe5_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe5_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe5_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe5_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe5_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe5_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe5_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe5_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe5_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe5_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe5_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe5_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe5_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe5_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe5_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe5_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe5_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe5_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe5_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe5_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe5_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe5_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe5_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe5_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe5_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe5_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe5_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe5_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe5_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe5_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe5_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe5_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe5_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe5_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe5_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe5_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe5_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe5_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe5_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe5_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe5_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe5_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe5_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe5_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe5_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe5_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe5_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe5_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe5_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe5_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe5_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe5_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe5_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe5_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe5_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe5_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe5_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe5_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe5_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe5_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe5_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe5_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe5_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe5_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe5_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe5_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe5_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe5_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe5_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe5_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe5_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe5_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe5_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe5_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe5_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe5_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe5_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe5_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe5_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe5_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe5_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe5_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe5_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe5_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe5_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe5_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe5_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe5_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe5_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe5_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe5_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe5_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe5_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe5_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe5_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe5_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe5_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe5_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe5_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe5_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe5_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe5_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe5_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe5_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe5_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe5_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe5_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe5_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe5_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe5_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe5_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe5_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe5_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe5_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe5_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe5_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe5_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe5_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe5_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe5_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe5_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe5_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe5_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe5_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe5_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe5_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe5_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe5_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe5_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe5_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe5_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe5_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe5_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe5_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe5_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe5_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe5_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe5_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe5_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe5_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe5_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe5_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe5_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe5_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe5_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe5_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe5_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe5_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe5_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe5_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe5_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe5_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe5_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe5_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe5_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe5_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe5_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe5_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe5_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe5_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe5_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe5_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe5_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe5_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe5_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe5_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe5_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe5_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe5_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe5_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe5_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe5_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe5_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe5_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe5_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe5_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe5_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe5_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe5_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe5_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe5_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe5_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe5_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe5_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe5_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe5_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe5_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe5_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe5_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe5_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe5_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe5_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe5_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe5_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe5_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe5_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe5_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe5_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe5_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe5_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe5_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe5_io_pipe_phv_out_is_valid_processor),
    .io_hash_depth_0(pipe5_io_hash_depth_0),
    .io_hash_depth_1(pipe5_io_hash_depth_1),
    .io_key_in(pipe5_io_key_in),
    .io_key_out(pipe5_io_key_out),
    .io_sum_in(pipe5_io_sum_in),
    .io_sum_out(pipe5_io_sum_out),
    .io_val_in(pipe5_io_val_in),
    .io_val_out(pipe5_io_val_out)
  );
  HashReshapeLevel_2 pipe6 ( // @[hash.scala 106:23]
    .clock(pipe6_clock),
    .io_pipe_phv_in_data_0(pipe6_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe6_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe6_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe6_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe6_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe6_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe6_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe6_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe6_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe6_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe6_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe6_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe6_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe6_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe6_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe6_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe6_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe6_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe6_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe6_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe6_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe6_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe6_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe6_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe6_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe6_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe6_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe6_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe6_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe6_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe6_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe6_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe6_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe6_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe6_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe6_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe6_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe6_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe6_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe6_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe6_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe6_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe6_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe6_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe6_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe6_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe6_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe6_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe6_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe6_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe6_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe6_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe6_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe6_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe6_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe6_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe6_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe6_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe6_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe6_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe6_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe6_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe6_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe6_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe6_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe6_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe6_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe6_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe6_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe6_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe6_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe6_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe6_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe6_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe6_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe6_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe6_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe6_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe6_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe6_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe6_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe6_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe6_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe6_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe6_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe6_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe6_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe6_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe6_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe6_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe6_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe6_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe6_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe6_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe6_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe6_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe6_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe6_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe6_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe6_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe6_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe6_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe6_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe6_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe6_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe6_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe6_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe6_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe6_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe6_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe6_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe6_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe6_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe6_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe6_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe6_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe6_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe6_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe6_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe6_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe6_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe6_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe6_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe6_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe6_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe6_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe6_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe6_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe6_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe6_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe6_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe6_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe6_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe6_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe6_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe6_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe6_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe6_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe6_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe6_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe6_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe6_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe6_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe6_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe6_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe6_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe6_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe6_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe6_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe6_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe6_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe6_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe6_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe6_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe6_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe6_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe6_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe6_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe6_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe6_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe6_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe6_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe6_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe6_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe6_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe6_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe6_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe6_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe6_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe6_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe6_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe6_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe6_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe6_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe6_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe6_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe6_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe6_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe6_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe6_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe6_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe6_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe6_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe6_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe6_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe6_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe6_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe6_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe6_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe6_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe6_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe6_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe6_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe6_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe6_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe6_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe6_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe6_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe6_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe6_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe6_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe6_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe6_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe6_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe6_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe6_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe6_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe6_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe6_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe6_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe6_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe6_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe6_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe6_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe6_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe6_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe6_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe6_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe6_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe6_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe6_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe6_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe6_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe6_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe6_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe6_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe6_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe6_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe6_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe6_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe6_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe6_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe6_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe6_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe6_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe6_io_pipe_phv_out_is_valid_processor),
    .io_hash_depth_0(pipe6_io_hash_depth_0),
    .io_hash_depth_1(pipe6_io_hash_depth_1),
    .io_key_in(pipe6_io_key_in),
    .io_key_out(pipe6_io_key_out),
    .io_sum_in(pipe6_io_sum_in),
    .io_sum_out(pipe6_io_sum_out),
    .io_val_in(pipe6_io_val_in),
    .io_val_out(pipe6_io_val_out)
  );
  assign io_pipe_phv_out_data_0 = pipe6_io_pipe_phv_out_data_0; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_1 = pipe6_io_pipe_phv_out_data_1; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_2 = pipe6_io_pipe_phv_out_data_2; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_3 = pipe6_io_pipe_phv_out_data_3; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_4 = pipe6_io_pipe_phv_out_data_4; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_5 = pipe6_io_pipe_phv_out_data_5; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_6 = pipe6_io_pipe_phv_out_data_6; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_7 = pipe6_io_pipe_phv_out_data_7; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_8 = pipe6_io_pipe_phv_out_data_8; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_9 = pipe6_io_pipe_phv_out_data_9; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_10 = pipe6_io_pipe_phv_out_data_10; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_11 = pipe6_io_pipe_phv_out_data_11; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_12 = pipe6_io_pipe_phv_out_data_12; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_13 = pipe6_io_pipe_phv_out_data_13; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_14 = pipe6_io_pipe_phv_out_data_14; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_15 = pipe6_io_pipe_phv_out_data_15; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_16 = pipe6_io_pipe_phv_out_data_16; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_17 = pipe6_io_pipe_phv_out_data_17; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_18 = pipe6_io_pipe_phv_out_data_18; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_19 = pipe6_io_pipe_phv_out_data_19; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_20 = pipe6_io_pipe_phv_out_data_20; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_21 = pipe6_io_pipe_phv_out_data_21; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_22 = pipe6_io_pipe_phv_out_data_22; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_23 = pipe6_io_pipe_phv_out_data_23; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_24 = pipe6_io_pipe_phv_out_data_24; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_25 = pipe6_io_pipe_phv_out_data_25; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_26 = pipe6_io_pipe_phv_out_data_26; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_27 = pipe6_io_pipe_phv_out_data_27; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_28 = pipe6_io_pipe_phv_out_data_28; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_29 = pipe6_io_pipe_phv_out_data_29; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_30 = pipe6_io_pipe_phv_out_data_30; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_31 = pipe6_io_pipe_phv_out_data_31; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_32 = pipe6_io_pipe_phv_out_data_32; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_33 = pipe6_io_pipe_phv_out_data_33; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_34 = pipe6_io_pipe_phv_out_data_34; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_35 = pipe6_io_pipe_phv_out_data_35; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_36 = pipe6_io_pipe_phv_out_data_36; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_37 = pipe6_io_pipe_phv_out_data_37; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_38 = pipe6_io_pipe_phv_out_data_38; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_39 = pipe6_io_pipe_phv_out_data_39; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_40 = pipe6_io_pipe_phv_out_data_40; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_41 = pipe6_io_pipe_phv_out_data_41; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_42 = pipe6_io_pipe_phv_out_data_42; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_43 = pipe6_io_pipe_phv_out_data_43; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_44 = pipe6_io_pipe_phv_out_data_44; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_45 = pipe6_io_pipe_phv_out_data_45; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_46 = pipe6_io_pipe_phv_out_data_46; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_47 = pipe6_io_pipe_phv_out_data_47; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_48 = pipe6_io_pipe_phv_out_data_48; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_49 = pipe6_io_pipe_phv_out_data_49; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_50 = pipe6_io_pipe_phv_out_data_50; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_51 = pipe6_io_pipe_phv_out_data_51; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_52 = pipe6_io_pipe_phv_out_data_52; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_53 = pipe6_io_pipe_phv_out_data_53; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_54 = pipe6_io_pipe_phv_out_data_54; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_55 = pipe6_io_pipe_phv_out_data_55; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_56 = pipe6_io_pipe_phv_out_data_56; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_57 = pipe6_io_pipe_phv_out_data_57; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_58 = pipe6_io_pipe_phv_out_data_58; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_59 = pipe6_io_pipe_phv_out_data_59; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_60 = pipe6_io_pipe_phv_out_data_60; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_61 = pipe6_io_pipe_phv_out_data_61; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_62 = pipe6_io_pipe_phv_out_data_62; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_63 = pipe6_io_pipe_phv_out_data_63; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_64 = pipe6_io_pipe_phv_out_data_64; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_65 = pipe6_io_pipe_phv_out_data_65; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_66 = pipe6_io_pipe_phv_out_data_66; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_67 = pipe6_io_pipe_phv_out_data_67; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_68 = pipe6_io_pipe_phv_out_data_68; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_69 = pipe6_io_pipe_phv_out_data_69; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_70 = pipe6_io_pipe_phv_out_data_70; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_71 = pipe6_io_pipe_phv_out_data_71; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_72 = pipe6_io_pipe_phv_out_data_72; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_73 = pipe6_io_pipe_phv_out_data_73; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_74 = pipe6_io_pipe_phv_out_data_74; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_75 = pipe6_io_pipe_phv_out_data_75; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_76 = pipe6_io_pipe_phv_out_data_76; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_77 = pipe6_io_pipe_phv_out_data_77; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_78 = pipe6_io_pipe_phv_out_data_78; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_79 = pipe6_io_pipe_phv_out_data_79; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_80 = pipe6_io_pipe_phv_out_data_80; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_81 = pipe6_io_pipe_phv_out_data_81; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_82 = pipe6_io_pipe_phv_out_data_82; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_83 = pipe6_io_pipe_phv_out_data_83; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_84 = pipe6_io_pipe_phv_out_data_84; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_85 = pipe6_io_pipe_phv_out_data_85; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_86 = pipe6_io_pipe_phv_out_data_86; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_87 = pipe6_io_pipe_phv_out_data_87; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_88 = pipe6_io_pipe_phv_out_data_88; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_89 = pipe6_io_pipe_phv_out_data_89; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_90 = pipe6_io_pipe_phv_out_data_90; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_91 = pipe6_io_pipe_phv_out_data_91; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_92 = pipe6_io_pipe_phv_out_data_92; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_93 = pipe6_io_pipe_phv_out_data_93; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_94 = pipe6_io_pipe_phv_out_data_94; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_95 = pipe6_io_pipe_phv_out_data_95; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_0 = pipe6_io_pipe_phv_out_header_0; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_1 = pipe6_io_pipe_phv_out_header_1; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_2 = pipe6_io_pipe_phv_out_header_2; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_3 = pipe6_io_pipe_phv_out_header_3; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_4 = pipe6_io_pipe_phv_out_header_4; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_5 = pipe6_io_pipe_phv_out_header_5; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_6 = pipe6_io_pipe_phv_out_header_6; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_7 = pipe6_io_pipe_phv_out_header_7; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_8 = pipe6_io_pipe_phv_out_header_8; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_9 = pipe6_io_pipe_phv_out_header_9; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_10 = pipe6_io_pipe_phv_out_header_10; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_11 = pipe6_io_pipe_phv_out_header_11; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_12 = pipe6_io_pipe_phv_out_header_12; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_13 = pipe6_io_pipe_phv_out_header_13; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_14 = pipe6_io_pipe_phv_out_header_14; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_15 = pipe6_io_pipe_phv_out_header_15; // @[hash.scala 138:27]
  assign io_pipe_phv_out_parse_current_state = pipe6_io_pipe_phv_out_parse_current_state; // @[hash.scala 138:27]
  assign io_pipe_phv_out_parse_current_offset = pipe6_io_pipe_phv_out_parse_current_offset; // @[hash.scala 138:27]
  assign io_pipe_phv_out_parse_transition_field = pipe6_io_pipe_phv_out_parse_transition_field; // @[hash.scala 138:27]
  assign io_pipe_phv_out_next_processor_id = pipe6_io_pipe_phv_out_next_processor_id; // @[hash.scala 138:27]
  assign io_pipe_phv_out_next_config_id = pipe6_io_pipe_phv_out_next_config_id; // @[hash.scala 138:27]
  assign io_pipe_phv_out_is_valid_processor = pipe6_io_pipe_phv_out_is_valid_processor; // @[hash.scala 138:27]
  assign io_key_out = pipe6_io_key_out; // @[hash.scala 139:27]
  assign io_hash_val = pipe6_io_sum_out[7:0]; // @[hash.scala 140:46]
  assign io_hash_val_cs = pipe6_io_val_out[7:5]; // @[hash.scala 141:46]
  assign pipe1_clock = clock;
  assign pipe1_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[hash.scala 108:27]
  assign pipe1_io_key_in = io_key_in; // @[hash.scala 109:27]
  assign pipe1_io_sum_in = io_key_in[15:0]; // @[hash.scala 110:39]
  assign pipe2_clock = clock;
  assign pipe2_io_pipe_phv_in_data_0 = pipe1_io_pipe_phv_out_data_0; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_1 = pipe1_io_pipe_phv_out_data_1; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_2 = pipe1_io_pipe_phv_out_data_2; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_3 = pipe1_io_pipe_phv_out_data_3; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_4 = pipe1_io_pipe_phv_out_data_4; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_5 = pipe1_io_pipe_phv_out_data_5; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_6 = pipe1_io_pipe_phv_out_data_6; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_7 = pipe1_io_pipe_phv_out_data_7; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_8 = pipe1_io_pipe_phv_out_data_8; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_9 = pipe1_io_pipe_phv_out_data_9; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_10 = pipe1_io_pipe_phv_out_data_10; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_11 = pipe1_io_pipe_phv_out_data_11; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_12 = pipe1_io_pipe_phv_out_data_12; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_13 = pipe1_io_pipe_phv_out_data_13; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_14 = pipe1_io_pipe_phv_out_data_14; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_15 = pipe1_io_pipe_phv_out_data_15; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_16 = pipe1_io_pipe_phv_out_data_16; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_17 = pipe1_io_pipe_phv_out_data_17; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_18 = pipe1_io_pipe_phv_out_data_18; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_19 = pipe1_io_pipe_phv_out_data_19; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_20 = pipe1_io_pipe_phv_out_data_20; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_21 = pipe1_io_pipe_phv_out_data_21; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_22 = pipe1_io_pipe_phv_out_data_22; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_23 = pipe1_io_pipe_phv_out_data_23; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_24 = pipe1_io_pipe_phv_out_data_24; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_25 = pipe1_io_pipe_phv_out_data_25; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_26 = pipe1_io_pipe_phv_out_data_26; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_27 = pipe1_io_pipe_phv_out_data_27; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_28 = pipe1_io_pipe_phv_out_data_28; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_29 = pipe1_io_pipe_phv_out_data_29; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_30 = pipe1_io_pipe_phv_out_data_30; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_31 = pipe1_io_pipe_phv_out_data_31; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_32 = pipe1_io_pipe_phv_out_data_32; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_33 = pipe1_io_pipe_phv_out_data_33; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_34 = pipe1_io_pipe_phv_out_data_34; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_35 = pipe1_io_pipe_phv_out_data_35; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_36 = pipe1_io_pipe_phv_out_data_36; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_37 = pipe1_io_pipe_phv_out_data_37; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_38 = pipe1_io_pipe_phv_out_data_38; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_39 = pipe1_io_pipe_phv_out_data_39; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_40 = pipe1_io_pipe_phv_out_data_40; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_41 = pipe1_io_pipe_phv_out_data_41; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_42 = pipe1_io_pipe_phv_out_data_42; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_43 = pipe1_io_pipe_phv_out_data_43; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_44 = pipe1_io_pipe_phv_out_data_44; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_45 = pipe1_io_pipe_phv_out_data_45; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_46 = pipe1_io_pipe_phv_out_data_46; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_47 = pipe1_io_pipe_phv_out_data_47; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_48 = pipe1_io_pipe_phv_out_data_48; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_49 = pipe1_io_pipe_phv_out_data_49; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_50 = pipe1_io_pipe_phv_out_data_50; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_51 = pipe1_io_pipe_phv_out_data_51; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_52 = pipe1_io_pipe_phv_out_data_52; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_53 = pipe1_io_pipe_phv_out_data_53; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_54 = pipe1_io_pipe_phv_out_data_54; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_55 = pipe1_io_pipe_phv_out_data_55; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_56 = pipe1_io_pipe_phv_out_data_56; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_57 = pipe1_io_pipe_phv_out_data_57; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_58 = pipe1_io_pipe_phv_out_data_58; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_59 = pipe1_io_pipe_phv_out_data_59; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_60 = pipe1_io_pipe_phv_out_data_60; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_61 = pipe1_io_pipe_phv_out_data_61; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_62 = pipe1_io_pipe_phv_out_data_62; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_63 = pipe1_io_pipe_phv_out_data_63; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_64 = pipe1_io_pipe_phv_out_data_64; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_65 = pipe1_io_pipe_phv_out_data_65; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_66 = pipe1_io_pipe_phv_out_data_66; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_67 = pipe1_io_pipe_phv_out_data_67; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_68 = pipe1_io_pipe_phv_out_data_68; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_69 = pipe1_io_pipe_phv_out_data_69; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_70 = pipe1_io_pipe_phv_out_data_70; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_71 = pipe1_io_pipe_phv_out_data_71; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_72 = pipe1_io_pipe_phv_out_data_72; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_73 = pipe1_io_pipe_phv_out_data_73; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_74 = pipe1_io_pipe_phv_out_data_74; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_75 = pipe1_io_pipe_phv_out_data_75; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_76 = pipe1_io_pipe_phv_out_data_76; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_77 = pipe1_io_pipe_phv_out_data_77; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_78 = pipe1_io_pipe_phv_out_data_78; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_79 = pipe1_io_pipe_phv_out_data_79; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_80 = pipe1_io_pipe_phv_out_data_80; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_81 = pipe1_io_pipe_phv_out_data_81; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_82 = pipe1_io_pipe_phv_out_data_82; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_83 = pipe1_io_pipe_phv_out_data_83; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_84 = pipe1_io_pipe_phv_out_data_84; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_85 = pipe1_io_pipe_phv_out_data_85; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_86 = pipe1_io_pipe_phv_out_data_86; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_87 = pipe1_io_pipe_phv_out_data_87; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_88 = pipe1_io_pipe_phv_out_data_88; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_89 = pipe1_io_pipe_phv_out_data_89; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_90 = pipe1_io_pipe_phv_out_data_90; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_91 = pipe1_io_pipe_phv_out_data_91; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_92 = pipe1_io_pipe_phv_out_data_92; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_93 = pipe1_io_pipe_phv_out_data_93; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_94 = pipe1_io_pipe_phv_out_data_94; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_95 = pipe1_io_pipe_phv_out_data_95; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_0 = pipe1_io_pipe_phv_out_header_0; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_1 = pipe1_io_pipe_phv_out_header_1; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_2 = pipe1_io_pipe_phv_out_header_2; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_3 = pipe1_io_pipe_phv_out_header_3; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_4 = pipe1_io_pipe_phv_out_header_4; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_5 = pipe1_io_pipe_phv_out_header_5; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_6 = pipe1_io_pipe_phv_out_header_6; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_7 = pipe1_io_pipe_phv_out_header_7; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_8 = pipe1_io_pipe_phv_out_header_8; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_9 = pipe1_io_pipe_phv_out_header_9; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_10 = pipe1_io_pipe_phv_out_header_10; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_11 = pipe1_io_pipe_phv_out_header_11; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_12 = pipe1_io_pipe_phv_out_header_12; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_13 = pipe1_io_pipe_phv_out_header_13; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_14 = pipe1_io_pipe_phv_out_header_14; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_15 = pipe1_io_pipe_phv_out_header_15; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_parse_current_state = pipe1_io_pipe_phv_out_parse_current_state; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_parse_current_offset = pipe1_io_pipe_phv_out_parse_current_offset; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_parse_transition_field = pipe1_io_pipe_phv_out_parse_transition_field; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_next_processor_id = pipe1_io_pipe_phv_out_next_processor_id; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_next_config_id = pipe1_io_pipe_phv_out_next_config_id; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_is_valid_processor = pipe1_io_pipe_phv_out_is_valid_processor; // @[hash.scala 112:27]
  assign pipe2_io_key_in = pipe1_io_key_out; // @[hash.scala 113:27]
  assign pipe2_io_sum_in = pipe1_io_sum_out; // @[hash.scala 114:27]
  assign pipe3_clock = clock;
  assign pipe3_io_pipe_phv_in_data_0 = pipe2_io_pipe_phv_out_data_0; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_1 = pipe2_io_pipe_phv_out_data_1; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_2 = pipe2_io_pipe_phv_out_data_2; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_3 = pipe2_io_pipe_phv_out_data_3; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_4 = pipe2_io_pipe_phv_out_data_4; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_5 = pipe2_io_pipe_phv_out_data_5; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_6 = pipe2_io_pipe_phv_out_data_6; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_7 = pipe2_io_pipe_phv_out_data_7; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_8 = pipe2_io_pipe_phv_out_data_8; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_9 = pipe2_io_pipe_phv_out_data_9; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_10 = pipe2_io_pipe_phv_out_data_10; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_11 = pipe2_io_pipe_phv_out_data_11; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_12 = pipe2_io_pipe_phv_out_data_12; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_13 = pipe2_io_pipe_phv_out_data_13; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_14 = pipe2_io_pipe_phv_out_data_14; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_15 = pipe2_io_pipe_phv_out_data_15; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_16 = pipe2_io_pipe_phv_out_data_16; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_17 = pipe2_io_pipe_phv_out_data_17; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_18 = pipe2_io_pipe_phv_out_data_18; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_19 = pipe2_io_pipe_phv_out_data_19; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_20 = pipe2_io_pipe_phv_out_data_20; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_21 = pipe2_io_pipe_phv_out_data_21; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_22 = pipe2_io_pipe_phv_out_data_22; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_23 = pipe2_io_pipe_phv_out_data_23; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_24 = pipe2_io_pipe_phv_out_data_24; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_25 = pipe2_io_pipe_phv_out_data_25; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_26 = pipe2_io_pipe_phv_out_data_26; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_27 = pipe2_io_pipe_phv_out_data_27; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_28 = pipe2_io_pipe_phv_out_data_28; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_29 = pipe2_io_pipe_phv_out_data_29; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_30 = pipe2_io_pipe_phv_out_data_30; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_31 = pipe2_io_pipe_phv_out_data_31; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_32 = pipe2_io_pipe_phv_out_data_32; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_33 = pipe2_io_pipe_phv_out_data_33; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_34 = pipe2_io_pipe_phv_out_data_34; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_35 = pipe2_io_pipe_phv_out_data_35; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_36 = pipe2_io_pipe_phv_out_data_36; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_37 = pipe2_io_pipe_phv_out_data_37; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_38 = pipe2_io_pipe_phv_out_data_38; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_39 = pipe2_io_pipe_phv_out_data_39; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_40 = pipe2_io_pipe_phv_out_data_40; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_41 = pipe2_io_pipe_phv_out_data_41; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_42 = pipe2_io_pipe_phv_out_data_42; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_43 = pipe2_io_pipe_phv_out_data_43; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_44 = pipe2_io_pipe_phv_out_data_44; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_45 = pipe2_io_pipe_phv_out_data_45; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_46 = pipe2_io_pipe_phv_out_data_46; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_47 = pipe2_io_pipe_phv_out_data_47; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_48 = pipe2_io_pipe_phv_out_data_48; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_49 = pipe2_io_pipe_phv_out_data_49; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_50 = pipe2_io_pipe_phv_out_data_50; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_51 = pipe2_io_pipe_phv_out_data_51; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_52 = pipe2_io_pipe_phv_out_data_52; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_53 = pipe2_io_pipe_phv_out_data_53; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_54 = pipe2_io_pipe_phv_out_data_54; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_55 = pipe2_io_pipe_phv_out_data_55; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_56 = pipe2_io_pipe_phv_out_data_56; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_57 = pipe2_io_pipe_phv_out_data_57; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_58 = pipe2_io_pipe_phv_out_data_58; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_59 = pipe2_io_pipe_phv_out_data_59; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_60 = pipe2_io_pipe_phv_out_data_60; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_61 = pipe2_io_pipe_phv_out_data_61; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_62 = pipe2_io_pipe_phv_out_data_62; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_63 = pipe2_io_pipe_phv_out_data_63; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_64 = pipe2_io_pipe_phv_out_data_64; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_65 = pipe2_io_pipe_phv_out_data_65; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_66 = pipe2_io_pipe_phv_out_data_66; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_67 = pipe2_io_pipe_phv_out_data_67; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_68 = pipe2_io_pipe_phv_out_data_68; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_69 = pipe2_io_pipe_phv_out_data_69; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_70 = pipe2_io_pipe_phv_out_data_70; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_71 = pipe2_io_pipe_phv_out_data_71; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_72 = pipe2_io_pipe_phv_out_data_72; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_73 = pipe2_io_pipe_phv_out_data_73; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_74 = pipe2_io_pipe_phv_out_data_74; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_75 = pipe2_io_pipe_phv_out_data_75; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_76 = pipe2_io_pipe_phv_out_data_76; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_77 = pipe2_io_pipe_phv_out_data_77; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_78 = pipe2_io_pipe_phv_out_data_78; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_79 = pipe2_io_pipe_phv_out_data_79; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_80 = pipe2_io_pipe_phv_out_data_80; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_81 = pipe2_io_pipe_phv_out_data_81; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_82 = pipe2_io_pipe_phv_out_data_82; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_83 = pipe2_io_pipe_phv_out_data_83; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_84 = pipe2_io_pipe_phv_out_data_84; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_85 = pipe2_io_pipe_phv_out_data_85; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_86 = pipe2_io_pipe_phv_out_data_86; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_87 = pipe2_io_pipe_phv_out_data_87; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_88 = pipe2_io_pipe_phv_out_data_88; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_89 = pipe2_io_pipe_phv_out_data_89; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_90 = pipe2_io_pipe_phv_out_data_90; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_91 = pipe2_io_pipe_phv_out_data_91; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_92 = pipe2_io_pipe_phv_out_data_92; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_93 = pipe2_io_pipe_phv_out_data_93; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_94 = pipe2_io_pipe_phv_out_data_94; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_95 = pipe2_io_pipe_phv_out_data_95; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_0 = pipe2_io_pipe_phv_out_header_0; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_1 = pipe2_io_pipe_phv_out_header_1; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_2 = pipe2_io_pipe_phv_out_header_2; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_3 = pipe2_io_pipe_phv_out_header_3; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_4 = pipe2_io_pipe_phv_out_header_4; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_5 = pipe2_io_pipe_phv_out_header_5; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_6 = pipe2_io_pipe_phv_out_header_6; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_7 = pipe2_io_pipe_phv_out_header_7; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_8 = pipe2_io_pipe_phv_out_header_8; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_9 = pipe2_io_pipe_phv_out_header_9; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_10 = pipe2_io_pipe_phv_out_header_10; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_11 = pipe2_io_pipe_phv_out_header_11; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_12 = pipe2_io_pipe_phv_out_header_12; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_13 = pipe2_io_pipe_phv_out_header_13; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_14 = pipe2_io_pipe_phv_out_header_14; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_15 = pipe2_io_pipe_phv_out_header_15; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_parse_current_state = pipe2_io_pipe_phv_out_parse_current_state; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_parse_current_offset = pipe2_io_pipe_phv_out_parse_current_offset; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_parse_transition_field = pipe2_io_pipe_phv_out_parse_transition_field; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_next_processor_id = pipe2_io_pipe_phv_out_next_processor_id; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_next_config_id = pipe2_io_pipe_phv_out_next_config_id; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_is_valid_processor = pipe2_io_pipe_phv_out_is_valid_processor; // @[hash.scala 116:27]
  assign pipe3_io_key_in = pipe2_io_key_out; // @[hash.scala 117:27]
  assign pipe3_io_sum_in = pipe2_io_sum_out; // @[hash.scala 118:27]
  assign pipe4_clock = clock;
  assign pipe4_io_pipe_phv_in_data_0 = pipe3_io_pipe_phv_out_data_0; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_1 = pipe3_io_pipe_phv_out_data_1; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_2 = pipe3_io_pipe_phv_out_data_2; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_3 = pipe3_io_pipe_phv_out_data_3; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_4 = pipe3_io_pipe_phv_out_data_4; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_5 = pipe3_io_pipe_phv_out_data_5; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_6 = pipe3_io_pipe_phv_out_data_6; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_7 = pipe3_io_pipe_phv_out_data_7; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_8 = pipe3_io_pipe_phv_out_data_8; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_9 = pipe3_io_pipe_phv_out_data_9; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_10 = pipe3_io_pipe_phv_out_data_10; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_11 = pipe3_io_pipe_phv_out_data_11; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_12 = pipe3_io_pipe_phv_out_data_12; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_13 = pipe3_io_pipe_phv_out_data_13; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_14 = pipe3_io_pipe_phv_out_data_14; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_15 = pipe3_io_pipe_phv_out_data_15; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_16 = pipe3_io_pipe_phv_out_data_16; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_17 = pipe3_io_pipe_phv_out_data_17; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_18 = pipe3_io_pipe_phv_out_data_18; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_19 = pipe3_io_pipe_phv_out_data_19; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_20 = pipe3_io_pipe_phv_out_data_20; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_21 = pipe3_io_pipe_phv_out_data_21; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_22 = pipe3_io_pipe_phv_out_data_22; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_23 = pipe3_io_pipe_phv_out_data_23; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_24 = pipe3_io_pipe_phv_out_data_24; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_25 = pipe3_io_pipe_phv_out_data_25; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_26 = pipe3_io_pipe_phv_out_data_26; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_27 = pipe3_io_pipe_phv_out_data_27; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_28 = pipe3_io_pipe_phv_out_data_28; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_29 = pipe3_io_pipe_phv_out_data_29; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_30 = pipe3_io_pipe_phv_out_data_30; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_31 = pipe3_io_pipe_phv_out_data_31; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_32 = pipe3_io_pipe_phv_out_data_32; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_33 = pipe3_io_pipe_phv_out_data_33; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_34 = pipe3_io_pipe_phv_out_data_34; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_35 = pipe3_io_pipe_phv_out_data_35; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_36 = pipe3_io_pipe_phv_out_data_36; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_37 = pipe3_io_pipe_phv_out_data_37; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_38 = pipe3_io_pipe_phv_out_data_38; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_39 = pipe3_io_pipe_phv_out_data_39; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_40 = pipe3_io_pipe_phv_out_data_40; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_41 = pipe3_io_pipe_phv_out_data_41; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_42 = pipe3_io_pipe_phv_out_data_42; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_43 = pipe3_io_pipe_phv_out_data_43; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_44 = pipe3_io_pipe_phv_out_data_44; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_45 = pipe3_io_pipe_phv_out_data_45; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_46 = pipe3_io_pipe_phv_out_data_46; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_47 = pipe3_io_pipe_phv_out_data_47; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_48 = pipe3_io_pipe_phv_out_data_48; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_49 = pipe3_io_pipe_phv_out_data_49; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_50 = pipe3_io_pipe_phv_out_data_50; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_51 = pipe3_io_pipe_phv_out_data_51; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_52 = pipe3_io_pipe_phv_out_data_52; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_53 = pipe3_io_pipe_phv_out_data_53; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_54 = pipe3_io_pipe_phv_out_data_54; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_55 = pipe3_io_pipe_phv_out_data_55; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_56 = pipe3_io_pipe_phv_out_data_56; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_57 = pipe3_io_pipe_phv_out_data_57; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_58 = pipe3_io_pipe_phv_out_data_58; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_59 = pipe3_io_pipe_phv_out_data_59; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_60 = pipe3_io_pipe_phv_out_data_60; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_61 = pipe3_io_pipe_phv_out_data_61; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_62 = pipe3_io_pipe_phv_out_data_62; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_63 = pipe3_io_pipe_phv_out_data_63; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_64 = pipe3_io_pipe_phv_out_data_64; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_65 = pipe3_io_pipe_phv_out_data_65; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_66 = pipe3_io_pipe_phv_out_data_66; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_67 = pipe3_io_pipe_phv_out_data_67; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_68 = pipe3_io_pipe_phv_out_data_68; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_69 = pipe3_io_pipe_phv_out_data_69; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_70 = pipe3_io_pipe_phv_out_data_70; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_71 = pipe3_io_pipe_phv_out_data_71; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_72 = pipe3_io_pipe_phv_out_data_72; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_73 = pipe3_io_pipe_phv_out_data_73; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_74 = pipe3_io_pipe_phv_out_data_74; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_75 = pipe3_io_pipe_phv_out_data_75; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_76 = pipe3_io_pipe_phv_out_data_76; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_77 = pipe3_io_pipe_phv_out_data_77; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_78 = pipe3_io_pipe_phv_out_data_78; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_79 = pipe3_io_pipe_phv_out_data_79; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_80 = pipe3_io_pipe_phv_out_data_80; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_81 = pipe3_io_pipe_phv_out_data_81; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_82 = pipe3_io_pipe_phv_out_data_82; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_83 = pipe3_io_pipe_phv_out_data_83; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_84 = pipe3_io_pipe_phv_out_data_84; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_85 = pipe3_io_pipe_phv_out_data_85; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_86 = pipe3_io_pipe_phv_out_data_86; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_87 = pipe3_io_pipe_phv_out_data_87; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_88 = pipe3_io_pipe_phv_out_data_88; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_89 = pipe3_io_pipe_phv_out_data_89; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_90 = pipe3_io_pipe_phv_out_data_90; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_91 = pipe3_io_pipe_phv_out_data_91; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_92 = pipe3_io_pipe_phv_out_data_92; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_93 = pipe3_io_pipe_phv_out_data_93; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_94 = pipe3_io_pipe_phv_out_data_94; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_95 = pipe3_io_pipe_phv_out_data_95; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_0 = pipe3_io_pipe_phv_out_header_0; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_1 = pipe3_io_pipe_phv_out_header_1; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_2 = pipe3_io_pipe_phv_out_header_2; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_3 = pipe3_io_pipe_phv_out_header_3; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_4 = pipe3_io_pipe_phv_out_header_4; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_5 = pipe3_io_pipe_phv_out_header_5; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_6 = pipe3_io_pipe_phv_out_header_6; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_7 = pipe3_io_pipe_phv_out_header_7; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_8 = pipe3_io_pipe_phv_out_header_8; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_9 = pipe3_io_pipe_phv_out_header_9; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_10 = pipe3_io_pipe_phv_out_header_10; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_11 = pipe3_io_pipe_phv_out_header_11; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_12 = pipe3_io_pipe_phv_out_header_12; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_13 = pipe3_io_pipe_phv_out_header_13; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_14 = pipe3_io_pipe_phv_out_header_14; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_15 = pipe3_io_pipe_phv_out_header_15; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_parse_current_state = pipe3_io_pipe_phv_out_parse_current_state; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_parse_current_offset = pipe3_io_pipe_phv_out_parse_current_offset; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_parse_transition_field = pipe3_io_pipe_phv_out_parse_transition_field; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_next_processor_id = pipe3_io_pipe_phv_out_next_processor_id; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_next_config_id = pipe3_io_pipe_phv_out_next_config_id; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_is_valid_processor = pipe3_io_pipe_phv_out_is_valid_processor; // @[hash.scala 120:27]
  assign pipe4_io_hash_depth_0 = hash_depth_0; // @[hash.scala 124:27]
  assign pipe4_io_hash_depth_1 = hash_depth_1; // @[hash.scala 124:27]
  assign pipe4_io_key_in = pipe3_io_key_out; // @[hash.scala 121:27]
  assign pipe4_io_sum_in = pipe3_io_sum_out; // @[hash.scala 122:27]
  assign pipe5_clock = clock;
  assign pipe5_io_pipe_phv_in_data_0 = pipe4_io_pipe_phv_out_data_0; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_1 = pipe4_io_pipe_phv_out_data_1; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_2 = pipe4_io_pipe_phv_out_data_2; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_3 = pipe4_io_pipe_phv_out_data_3; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_4 = pipe4_io_pipe_phv_out_data_4; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_5 = pipe4_io_pipe_phv_out_data_5; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_6 = pipe4_io_pipe_phv_out_data_6; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_7 = pipe4_io_pipe_phv_out_data_7; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_8 = pipe4_io_pipe_phv_out_data_8; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_9 = pipe4_io_pipe_phv_out_data_9; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_10 = pipe4_io_pipe_phv_out_data_10; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_11 = pipe4_io_pipe_phv_out_data_11; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_12 = pipe4_io_pipe_phv_out_data_12; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_13 = pipe4_io_pipe_phv_out_data_13; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_14 = pipe4_io_pipe_phv_out_data_14; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_15 = pipe4_io_pipe_phv_out_data_15; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_16 = pipe4_io_pipe_phv_out_data_16; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_17 = pipe4_io_pipe_phv_out_data_17; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_18 = pipe4_io_pipe_phv_out_data_18; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_19 = pipe4_io_pipe_phv_out_data_19; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_20 = pipe4_io_pipe_phv_out_data_20; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_21 = pipe4_io_pipe_phv_out_data_21; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_22 = pipe4_io_pipe_phv_out_data_22; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_23 = pipe4_io_pipe_phv_out_data_23; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_24 = pipe4_io_pipe_phv_out_data_24; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_25 = pipe4_io_pipe_phv_out_data_25; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_26 = pipe4_io_pipe_phv_out_data_26; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_27 = pipe4_io_pipe_phv_out_data_27; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_28 = pipe4_io_pipe_phv_out_data_28; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_29 = pipe4_io_pipe_phv_out_data_29; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_30 = pipe4_io_pipe_phv_out_data_30; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_31 = pipe4_io_pipe_phv_out_data_31; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_32 = pipe4_io_pipe_phv_out_data_32; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_33 = pipe4_io_pipe_phv_out_data_33; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_34 = pipe4_io_pipe_phv_out_data_34; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_35 = pipe4_io_pipe_phv_out_data_35; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_36 = pipe4_io_pipe_phv_out_data_36; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_37 = pipe4_io_pipe_phv_out_data_37; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_38 = pipe4_io_pipe_phv_out_data_38; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_39 = pipe4_io_pipe_phv_out_data_39; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_40 = pipe4_io_pipe_phv_out_data_40; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_41 = pipe4_io_pipe_phv_out_data_41; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_42 = pipe4_io_pipe_phv_out_data_42; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_43 = pipe4_io_pipe_phv_out_data_43; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_44 = pipe4_io_pipe_phv_out_data_44; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_45 = pipe4_io_pipe_phv_out_data_45; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_46 = pipe4_io_pipe_phv_out_data_46; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_47 = pipe4_io_pipe_phv_out_data_47; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_48 = pipe4_io_pipe_phv_out_data_48; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_49 = pipe4_io_pipe_phv_out_data_49; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_50 = pipe4_io_pipe_phv_out_data_50; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_51 = pipe4_io_pipe_phv_out_data_51; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_52 = pipe4_io_pipe_phv_out_data_52; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_53 = pipe4_io_pipe_phv_out_data_53; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_54 = pipe4_io_pipe_phv_out_data_54; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_55 = pipe4_io_pipe_phv_out_data_55; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_56 = pipe4_io_pipe_phv_out_data_56; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_57 = pipe4_io_pipe_phv_out_data_57; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_58 = pipe4_io_pipe_phv_out_data_58; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_59 = pipe4_io_pipe_phv_out_data_59; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_60 = pipe4_io_pipe_phv_out_data_60; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_61 = pipe4_io_pipe_phv_out_data_61; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_62 = pipe4_io_pipe_phv_out_data_62; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_63 = pipe4_io_pipe_phv_out_data_63; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_64 = pipe4_io_pipe_phv_out_data_64; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_65 = pipe4_io_pipe_phv_out_data_65; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_66 = pipe4_io_pipe_phv_out_data_66; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_67 = pipe4_io_pipe_phv_out_data_67; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_68 = pipe4_io_pipe_phv_out_data_68; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_69 = pipe4_io_pipe_phv_out_data_69; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_70 = pipe4_io_pipe_phv_out_data_70; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_71 = pipe4_io_pipe_phv_out_data_71; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_72 = pipe4_io_pipe_phv_out_data_72; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_73 = pipe4_io_pipe_phv_out_data_73; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_74 = pipe4_io_pipe_phv_out_data_74; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_75 = pipe4_io_pipe_phv_out_data_75; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_76 = pipe4_io_pipe_phv_out_data_76; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_77 = pipe4_io_pipe_phv_out_data_77; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_78 = pipe4_io_pipe_phv_out_data_78; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_79 = pipe4_io_pipe_phv_out_data_79; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_80 = pipe4_io_pipe_phv_out_data_80; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_81 = pipe4_io_pipe_phv_out_data_81; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_82 = pipe4_io_pipe_phv_out_data_82; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_83 = pipe4_io_pipe_phv_out_data_83; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_84 = pipe4_io_pipe_phv_out_data_84; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_85 = pipe4_io_pipe_phv_out_data_85; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_86 = pipe4_io_pipe_phv_out_data_86; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_87 = pipe4_io_pipe_phv_out_data_87; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_88 = pipe4_io_pipe_phv_out_data_88; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_89 = pipe4_io_pipe_phv_out_data_89; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_90 = pipe4_io_pipe_phv_out_data_90; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_91 = pipe4_io_pipe_phv_out_data_91; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_92 = pipe4_io_pipe_phv_out_data_92; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_93 = pipe4_io_pipe_phv_out_data_93; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_94 = pipe4_io_pipe_phv_out_data_94; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_95 = pipe4_io_pipe_phv_out_data_95; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_0 = pipe4_io_pipe_phv_out_header_0; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_1 = pipe4_io_pipe_phv_out_header_1; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_2 = pipe4_io_pipe_phv_out_header_2; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_3 = pipe4_io_pipe_phv_out_header_3; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_4 = pipe4_io_pipe_phv_out_header_4; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_5 = pipe4_io_pipe_phv_out_header_5; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_6 = pipe4_io_pipe_phv_out_header_6; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_7 = pipe4_io_pipe_phv_out_header_7; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_8 = pipe4_io_pipe_phv_out_header_8; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_9 = pipe4_io_pipe_phv_out_header_9; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_10 = pipe4_io_pipe_phv_out_header_10; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_11 = pipe4_io_pipe_phv_out_header_11; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_12 = pipe4_io_pipe_phv_out_header_12; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_13 = pipe4_io_pipe_phv_out_header_13; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_14 = pipe4_io_pipe_phv_out_header_14; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_15 = pipe4_io_pipe_phv_out_header_15; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_parse_current_state = pipe4_io_pipe_phv_out_parse_current_state; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_parse_current_offset = pipe4_io_pipe_phv_out_parse_current_offset; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_parse_transition_field = pipe4_io_pipe_phv_out_parse_transition_field; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_next_processor_id = pipe4_io_pipe_phv_out_next_processor_id; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_next_config_id = pipe4_io_pipe_phv_out_next_config_id; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_is_valid_processor = pipe4_io_pipe_phv_out_is_valid_processor; // @[hash.scala 126:27]
  assign pipe5_io_hash_depth_0 = hash_depth_0; // @[hash.scala 130:27]
  assign pipe5_io_hash_depth_1 = hash_depth_1; // @[hash.scala 130:27]
  assign pipe5_io_key_in = pipe4_io_key_out; // @[hash.scala 127:27]
  assign pipe5_io_sum_in = pipe4_io_sum_out; // @[hash.scala 128:27]
  assign pipe5_io_val_in = pipe4_io_val_out; // @[hash.scala 129:27]
  assign pipe6_clock = clock;
  assign pipe6_io_pipe_phv_in_data_0 = pipe5_io_pipe_phv_out_data_0; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_1 = pipe5_io_pipe_phv_out_data_1; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_2 = pipe5_io_pipe_phv_out_data_2; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_3 = pipe5_io_pipe_phv_out_data_3; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_4 = pipe5_io_pipe_phv_out_data_4; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_5 = pipe5_io_pipe_phv_out_data_5; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_6 = pipe5_io_pipe_phv_out_data_6; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_7 = pipe5_io_pipe_phv_out_data_7; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_8 = pipe5_io_pipe_phv_out_data_8; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_9 = pipe5_io_pipe_phv_out_data_9; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_10 = pipe5_io_pipe_phv_out_data_10; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_11 = pipe5_io_pipe_phv_out_data_11; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_12 = pipe5_io_pipe_phv_out_data_12; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_13 = pipe5_io_pipe_phv_out_data_13; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_14 = pipe5_io_pipe_phv_out_data_14; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_15 = pipe5_io_pipe_phv_out_data_15; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_16 = pipe5_io_pipe_phv_out_data_16; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_17 = pipe5_io_pipe_phv_out_data_17; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_18 = pipe5_io_pipe_phv_out_data_18; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_19 = pipe5_io_pipe_phv_out_data_19; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_20 = pipe5_io_pipe_phv_out_data_20; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_21 = pipe5_io_pipe_phv_out_data_21; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_22 = pipe5_io_pipe_phv_out_data_22; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_23 = pipe5_io_pipe_phv_out_data_23; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_24 = pipe5_io_pipe_phv_out_data_24; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_25 = pipe5_io_pipe_phv_out_data_25; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_26 = pipe5_io_pipe_phv_out_data_26; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_27 = pipe5_io_pipe_phv_out_data_27; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_28 = pipe5_io_pipe_phv_out_data_28; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_29 = pipe5_io_pipe_phv_out_data_29; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_30 = pipe5_io_pipe_phv_out_data_30; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_31 = pipe5_io_pipe_phv_out_data_31; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_32 = pipe5_io_pipe_phv_out_data_32; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_33 = pipe5_io_pipe_phv_out_data_33; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_34 = pipe5_io_pipe_phv_out_data_34; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_35 = pipe5_io_pipe_phv_out_data_35; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_36 = pipe5_io_pipe_phv_out_data_36; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_37 = pipe5_io_pipe_phv_out_data_37; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_38 = pipe5_io_pipe_phv_out_data_38; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_39 = pipe5_io_pipe_phv_out_data_39; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_40 = pipe5_io_pipe_phv_out_data_40; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_41 = pipe5_io_pipe_phv_out_data_41; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_42 = pipe5_io_pipe_phv_out_data_42; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_43 = pipe5_io_pipe_phv_out_data_43; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_44 = pipe5_io_pipe_phv_out_data_44; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_45 = pipe5_io_pipe_phv_out_data_45; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_46 = pipe5_io_pipe_phv_out_data_46; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_47 = pipe5_io_pipe_phv_out_data_47; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_48 = pipe5_io_pipe_phv_out_data_48; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_49 = pipe5_io_pipe_phv_out_data_49; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_50 = pipe5_io_pipe_phv_out_data_50; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_51 = pipe5_io_pipe_phv_out_data_51; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_52 = pipe5_io_pipe_phv_out_data_52; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_53 = pipe5_io_pipe_phv_out_data_53; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_54 = pipe5_io_pipe_phv_out_data_54; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_55 = pipe5_io_pipe_phv_out_data_55; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_56 = pipe5_io_pipe_phv_out_data_56; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_57 = pipe5_io_pipe_phv_out_data_57; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_58 = pipe5_io_pipe_phv_out_data_58; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_59 = pipe5_io_pipe_phv_out_data_59; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_60 = pipe5_io_pipe_phv_out_data_60; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_61 = pipe5_io_pipe_phv_out_data_61; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_62 = pipe5_io_pipe_phv_out_data_62; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_63 = pipe5_io_pipe_phv_out_data_63; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_64 = pipe5_io_pipe_phv_out_data_64; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_65 = pipe5_io_pipe_phv_out_data_65; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_66 = pipe5_io_pipe_phv_out_data_66; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_67 = pipe5_io_pipe_phv_out_data_67; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_68 = pipe5_io_pipe_phv_out_data_68; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_69 = pipe5_io_pipe_phv_out_data_69; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_70 = pipe5_io_pipe_phv_out_data_70; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_71 = pipe5_io_pipe_phv_out_data_71; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_72 = pipe5_io_pipe_phv_out_data_72; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_73 = pipe5_io_pipe_phv_out_data_73; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_74 = pipe5_io_pipe_phv_out_data_74; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_75 = pipe5_io_pipe_phv_out_data_75; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_76 = pipe5_io_pipe_phv_out_data_76; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_77 = pipe5_io_pipe_phv_out_data_77; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_78 = pipe5_io_pipe_phv_out_data_78; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_79 = pipe5_io_pipe_phv_out_data_79; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_80 = pipe5_io_pipe_phv_out_data_80; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_81 = pipe5_io_pipe_phv_out_data_81; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_82 = pipe5_io_pipe_phv_out_data_82; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_83 = pipe5_io_pipe_phv_out_data_83; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_84 = pipe5_io_pipe_phv_out_data_84; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_85 = pipe5_io_pipe_phv_out_data_85; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_86 = pipe5_io_pipe_phv_out_data_86; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_87 = pipe5_io_pipe_phv_out_data_87; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_88 = pipe5_io_pipe_phv_out_data_88; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_89 = pipe5_io_pipe_phv_out_data_89; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_90 = pipe5_io_pipe_phv_out_data_90; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_91 = pipe5_io_pipe_phv_out_data_91; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_92 = pipe5_io_pipe_phv_out_data_92; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_93 = pipe5_io_pipe_phv_out_data_93; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_94 = pipe5_io_pipe_phv_out_data_94; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_95 = pipe5_io_pipe_phv_out_data_95; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_0 = pipe5_io_pipe_phv_out_header_0; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_1 = pipe5_io_pipe_phv_out_header_1; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_2 = pipe5_io_pipe_phv_out_header_2; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_3 = pipe5_io_pipe_phv_out_header_3; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_4 = pipe5_io_pipe_phv_out_header_4; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_5 = pipe5_io_pipe_phv_out_header_5; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_6 = pipe5_io_pipe_phv_out_header_6; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_7 = pipe5_io_pipe_phv_out_header_7; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_8 = pipe5_io_pipe_phv_out_header_8; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_9 = pipe5_io_pipe_phv_out_header_9; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_10 = pipe5_io_pipe_phv_out_header_10; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_11 = pipe5_io_pipe_phv_out_header_11; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_12 = pipe5_io_pipe_phv_out_header_12; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_13 = pipe5_io_pipe_phv_out_header_13; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_14 = pipe5_io_pipe_phv_out_header_14; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_15 = pipe5_io_pipe_phv_out_header_15; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_parse_current_state = pipe5_io_pipe_phv_out_parse_current_state; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_parse_current_offset = pipe5_io_pipe_phv_out_parse_current_offset; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_parse_transition_field = pipe5_io_pipe_phv_out_parse_transition_field; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_next_processor_id = pipe5_io_pipe_phv_out_next_processor_id; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_next_config_id = pipe5_io_pipe_phv_out_next_config_id; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_is_valid_processor = pipe5_io_pipe_phv_out_is_valid_processor; // @[hash.scala 132:27]
  assign pipe6_io_hash_depth_0 = hash_depth_0; // @[hash.scala 136:27]
  assign pipe6_io_hash_depth_1 = hash_depth_1; // @[hash.scala 136:27]
  assign pipe6_io_key_in = pipe5_io_key_out; // @[hash.scala 133:27]
  assign pipe6_io_sum_in = pipe5_io_sum_out; // @[hash.scala 134:27]
  assign pipe6_io_val_in = pipe5_io_val_out; // @[hash.scala 135:27]
  always @(posedge clock) begin
    if (io_mod_hash_depth_mod) begin // @[hash.scala 19:34]
      if (~io_mod_config_id) begin // @[hash.scala 20:38]
        hash_depth_0 <= io_mod_hash_depth; // @[hash.scala 20:38]
      end
    end
    if (io_mod_hash_depth_mod) begin // @[hash.scala 19:34]
      if (io_mod_config_id) begin // @[hash.scala 20:38]
        hash_depth_1 <= io_mod_hash_depth; // @[hash.scala 20:38]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  hash_depth_0 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  hash_depth_1 = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MatchGetCs(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input  [3:0]  io_table_config_0_table_width,
  input  [3:0]  io_table_config_0_table_depth,
  input  [3:0]  io_table_config_1_table_width,
  input  [3:0]  io_table_config_1_table_depth,
  input  [63:0] io_key_in,
  output [63:0] io_key_out,
  input  [7:0]  io_addr_in,
  output [7:0]  io_addr_out,
  input  [2:0]  io_cs_in,
  output [2:0]  io_cs_out,
  output        io_cs_vec_out_0,
  output        io_cs_vec_out_1,
  output        io_cs_vec_out_2,
  output        io_cs_vec_out_3,
  output        io_cs_vec_out_4,
  output        io_cs_vec_out_5,
  output        io_cs_vec_out_6,
  output        io_cs_vec_out_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[matcher.scala 102:22]
  reg [7:0] phv_data_1; // @[matcher.scala 102:22]
  reg [7:0] phv_data_2; // @[matcher.scala 102:22]
  reg [7:0] phv_data_3; // @[matcher.scala 102:22]
  reg [7:0] phv_data_4; // @[matcher.scala 102:22]
  reg [7:0] phv_data_5; // @[matcher.scala 102:22]
  reg [7:0] phv_data_6; // @[matcher.scala 102:22]
  reg [7:0] phv_data_7; // @[matcher.scala 102:22]
  reg [7:0] phv_data_8; // @[matcher.scala 102:22]
  reg [7:0] phv_data_9; // @[matcher.scala 102:22]
  reg [7:0] phv_data_10; // @[matcher.scala 102:22]
  reg [7:0] phv_data_11; // @[matcher.scala 102:22]
  reg [7:0] phv_data_12; // @[matcher.scala 102:22]
  reg [7:0] phv_data_13; // @[matcher.scala 102:22]
  reg [7:0] phv_data_14; // @[matcher.scala 102:22]
  reg [7:0] phv_data_15; // @[matcher.scala 102:22]
  reg [7:0] phv_data_16; // @[matcher.scala 102:22]
  reg [7:0] phv_data_17; // @[matcher.scala 102:22]
  reg [7:0] phv_data_18; // @[matcher.scala 102:22]
  reg [7:0] phv_data_19; // @[matcher.scala 102:22]
  reg [7:0] phv_data_20; // @[matcher.scala 102:22]
  reg [7:0] phv_data_21; // @[matcher.scala 102:22]
  reg [7:0] phv_data_22; // @[matcher.scala 102:22]
  reg [7:0] phv_data_23; // @[matcher.scala 102:22]
  reg [7:0] phv_data_24; // @[matcher.scala 102:22]
  reg [7:0] phv_data_25; // @[matcher.scala 102:22]
  reg [7:0] phv_data_26; // @[matcher.scala 102:22]
  reg [7:0] phv_data_27; // @[matcher.scala 102:22]
  reg [7:0] phv_data_28; // @[matcher.scala 102:22]
  reg [7:0] phv_data_29; // @[matcher.scala 102:22]
  reg [7:0] phv_data_30; // @[matcher.scala 102:22]
  reg [7:0] phv_data_31; // @[matcher.scala 102:22]
  reg [7:0] phv_data_32; // @[matcher.scala 102:22]
  reg [7:0] phv_data_33; // @[matcher.scala 102:22]
  reg [7:0] phv_data_34; // @[matcher.scala 102:22]
  reg [7:0] phv_data_35; // @[matcher.scala 102:22]
  reg [7:0] phv_data_36; // @[matcher.scala 102:22]
  reg [7:0] phv_data_37; // @[matcher.scala 102:22]
  reg [7:0] phv_data_38; // @[matcher.scala 102:22]
  reg [7:0] phv_data_39; // @[matcher.scala 102:22]
  reg [7:0] phv_data_40; // @[matcher.scala 102:22]
  reg [7:0] phv_data_41; // @[matcher.scala 102:22]
  reg [7:0] phv_data_42; // @[matcher.scala 102:22]
  reg [7:0] phv_data_43; // @[matcher.scala 102:22]
  reg [7:0] phv_data_44; // @[matcher.scala 102:22]
  reg [7:0] phv_data_45; // @[matcher.scala 102:22]
  reg [7:0] phv_data_46; // @[matcher.scala 102:22]
  reg [7:0] phv_data_47; // @[matcher.scala 102:22]
  reg [7:0] phv_data_48; // @[matcher.scala 102:22]
  reg [7:0] phv_data_49; // @[matcher.scala 102:22]
  reg [7:0] phv_data_50; // @[matcher.scala 102:22]
  reg [7:0] phv_data_51; // @[matcher.scala 102:22]
  reg [7:0] phv_data_52; // @[matcher.scala 102:22]
  reg [7:0] phv_data_53; // @[matcher.scala 102:22]
  reg [7:0] phv_data_54; // @[matcher.scala 102:22]
  reg [7:0] phv_data_55; // @[matcher.scala 102:22]
  reg [7:0] phv_data_56; // @[matcher.scala 102:22]
  reg [7:0] phv_data_57; // @[matcher.scala 102:22]
  reg [7:0] phv_data_58; // @[matcher.scala 102:22]
  reg [7:0] phv_data_59; // @[matcher.scala 102:22]
  reg [7:0] phv_data_60; // @[matcher.scala 102:22]
  reg [7:0] phv_data_61; // @[matcher.scala 102:22]
  reg [7:0] phv_data_62; // @[matcher.scala 102:22]
  reg [7:0] phv_data_63; // @[matcher.scala 102:22]
  reg [7:0] phv_data_64; // @[matcher.scala 102:22]
  reg [7:0] phv_data_65; // @[matcher.scala 102:22]
  reg [7:0] phv_data_66; // @[matcher.scala 102:22]
  reg [7:0] phv_data_67; // @[matcher.scala 102:22]
  reg [7:0] phv_data_68; // @[matcher.scala 102:22]
  reg [7:0] phv_data_69; // @[matcher.scala 102:22]
  reg [7:0] phv_data_70; // @[matcher.scala 102:22]
  reg [7:0] phv_data_71; // @[matcher.scala 102:22]
  reg [7:0] phv_data_72; // @[matcher.scala 102:22]
  reg [7:0] phv_data_73; // @[matcher.scala 102:22]
  reg [7:0] phv_data_74; // @[matcher.scala 102:22]
  reg [7:0] phv_data_75; // @[matcher.scala 102:22]
  reg [7:0] phv_data_76; // @[matcher.scala 102:22]
  reg [7:0] phv_data_77; // @[matcher.scala 102:22]
  reg [7:0] phv_data_78; // @[matcher.scala 102:22]
  reg [7:0] phv_data_79; // @[matcher.scala 102:22]
  reg [7:0] phv_data_80; // @[matcher.scala 102:22]
  reg [7:0] phv_data_81; // @[matcher.scala 102:22]
  reg [7:0] phv_data_82; // @[matcher.scala 102:22]
  reg [7:0] phv_data_83; // @[matcher.scala 102:22]
  reg [7:0] phv_data_84; // @[matcher.scala 102:22]
  reg [7:0] phv_data_85; // @[matcher.scala 102:22]
  reg [7:0] phv_data_86; // @[matcher.scala 102:22]
  reg [7:0] phv_data_87; // @[matcher.scala 102:22]
  reg [7:0] phv_data_88; // @[matcher.scala 102:22]
  reg [7:0] phv_data_89; // @[matcher.scala 102:22]
  reg [7:0] phv_data_90; // @[matcher.scala 102:22]
  reg [7:0] phv_data_91; // @[matcher.scala 102:22]
  reg [7:0] phv_data_92; // @[matcher.scala 102:22]
  reg [7:0] phv_data_93; // @[matcher.scala 102:22]
  reg [7:0] phv_data_94; // @[matcher.scala 102:22]
  reg [7:0] phv_data_95; // @[matcher.scala 102:22]
  reg [15:0] phv_header_0; // @[matcher.scala 102:22]
  reg [15:0] phv_header_1; // @[matcher.scala 102:22]
  reg [15:0] phv_header_2; // @[matcher.scala 102:22]
  reg [15:0] phv_header_3; // @[matcher.scala 102:22]
  reg [15:0] phv_header_4; // @[matcher.scala 102:22]
  reg [15:0] phv_header_5; // @[matcher.scala 102:22]
  reg [15:0] phv_header_6; // @[matcher.scala 102:22]
  reg [15:0] phv_header_7; // @[matcher.scala 102:22]
  reg [15:0] phv_header_8; // @[matcher.scala 102:22]
  reg [15:0] phv_header_9; // @[matcher.scala 102:22]
  reg [15:0] phv_header_10; // @[matcher.scala 102:22]
  reg [15:0] phv_header_11; // @[matcher.scala 102:22]
  reg [15:0] phv_header_12; // @[matcher.scala 102:22]
  reg [15:0] phv_header_13; // @[matcher.scala 102:22]
  reg [15:0] phv_header_14; // @[matcher.scala 102:22]
  reg [15:0] phv_header_15; // @[matcher.scala 102:22]
  reg [7:0] phv_parse_current_state; // @[matcher.scala 102:22]
  reg [7:0] phv_parse_current_offset; // @[matcher.scala 102:22]
  reg [15:0] phv_parse_transition_field; // @[matcher.scala 102:22]
  reg [1:0] phv_next_processor_id; // @[matcher.scala 102:22]
  reg  phv_next_config_id; // @[matcher.scala 102:22]
  reg  phv_is_valid_processor; // @[matcher.scala 102:22]
  reg [63:0] key; // @[matcher.scala 106:22]
  reg [7:0] addr; // @[matcher.scala 110:23]
  reg [2:0] cs; // @[matcher.scala 114:21]
  wire  _T = 3'h0 == cs; // @[matcher.scala 121:55]
  wire [3:0] _GEN_19 = phv_next_config_id ? io_table_config_1_table_width : io_table_config_0_table_width; // @[matcher.scala 124:84 matcher.scala 124:84]
  wire [3:0] _GEN_20 = phv_next_config_id ? io_table_config_1_table_depth : io_table_config_0_table_depth; // @[matcher.scala 124:84 matcher.scala 124:84]
  wire  width_extend = _GEN_19 == 4'h2; // @[matcher.scala 124:84]
  wire [3:0] _GEN_44 = {{1'd0}, cs}; // @[matcher.scala 125:39]
  wire [3:0] extended_cs = _GEN_44 + _GEN_20; // @[matcher.scala 125:39]
  wire  _GEN_21 = width_extend & 4'h0 == extended_cs | _T; // @[matcher.scala 126:88 matcher.scala 127:38]
  wire  _T_3 = 3'h1 == cs; // @[matcher.scala 121:55]
  wire  _GEN_24 = width_extend & 4'h1 == extended_cs | _T_3; // @[matcher.scala 126:88 matcher.scala 127:38]
  wire  _T_6 = 3'h2 == cs; // @[matcher.scala 121:55]
  wire  _GEN_27 = width_extend & 4'h2 == extended_cs | _T_6; // @[matcher.scala 126:88 matcher.scala 127:38]
  wire  _T_9 = 3'h3 == cs; // @[matcher.scala 121:55]
  wire  _GEN_30 = width_extend & 4'h3 == extended_cs | _T_9; // @[matcher.scala 126:88 matcher.scala 127:38]
  wire  _T_12 = 3'h4 == cs; // @[matcher.scala 121:55]
  wire  _GEN_33 = width_extend & 4'h4 == extended_cs | _T_12; // @[matcher.scala 126:88 matcher.scala 127:38]
  wire  _T_15 = 3'h5 == cs; // @[matcher.scala 121:55]
  wire  _GEN_36 = width_extend & 4'h5 == extended_cs | _T_15; // @[matcher.scala 126:88 matcher.scala 127:38]
  wire  _T_18 = 3'h6 == cs; // @[matcher.scala 121:55]
  wire  _GEN_39 = width_extend & 4'h6 == extended_cs | _T_18; // @[matcher.scala 126:88 matcher.scala 127:38]
  wire  _T_21 = 3'h7 == cs; // @[matcher.scala 121:55]
  wire  _GEN_42 = width_extend & 4'h7 == extended_cs | _T_21; // @[matcher.scala 126:88 matcher.scala 127:38]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[matcher.scala 104:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[matcher.scala 104:25]
  assign io_key_out = key; // @[matcher.scala 108:20]
  assign io_addr_out = addr; // @[matcher.scala 112:21]
  assign io_cs_out = cs; // @[matcher.scala 116:19]
  assign io_cs_vec_out_0 = phv_is_valid_processor & _GEN_21; // @[matcher.scala 120:43 matcher.scala 119:30]
  assign io_cs_vec_out_1 = phv_is_valid_processor & _GEN_24; // @[matcher.scala 120:43 matcher.scala 119:30]
  assign io_cs_vec_out_2 = phv_is_valid_processor & _GEN_27; // @[matcher.scala 120:43 matcher.scala 119:30]
  assign io_cs_vec_out_3 = phv_is_valid_processor & _GEN_30; // @[matcher.scala 120:43 matcher.scala 119:30]
  assign io_cs_vec_out_4 = phv_is_valid_processor & _GEN_33; // @[matcher.scala 120:43 matcher.scala 119:30]
  assign io_cs_vec_out_5 = phv_is_valid_processor & _GEN_36; // @[matcher.scala 120:43 matcher.scala 119:30]
  assign io_cs_vec_out_6 = phv_is_valid_processor & _GEN_39; // @[matcher.scala 120:43 matcher.scala 119:30]
  assign io_cs_vec_out_7 = phv_is_valid_processor & _GEN_42; // @[matcher.scala 120:43 matcher.scala 119:30]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[matcher.scala 103:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[matcher.scala 103:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[matcher.scala 103:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[matcher.scala 103:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[matcher.scala 103:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[matcher.scala 103:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[matcher.scala 103:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[matcher.scala 103:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[matcher.scala 103:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[matcher.scala 103:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[matcher.scala 103:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[matcher.scala 103:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[matcher.scala 103:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[matcher.scala 103:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[matcher.scala 103:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[matcher.scala 103:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[matcher.scala 103:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[matcher.scala 103:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[matcher.scala 103:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[matcher.scala 103:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[matcher.scala 103:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[matcher.scala 103:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[matcher.scala 103:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[matcher.scala 103:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[matcher.scala 103:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[matcher.scala 103:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[matcher.scala 103:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[matcher.scala 103:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[matcher.scala 103:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[matcher.scala 103:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[matcher.scala 103:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[matcher.scala 103:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[matcher.scala 103:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[matcher.scala 103:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[matcher.scala 103:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[matcher.scala 103:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[matcher.scala 103:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[matcher.scala 103:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[matcher.scala 103:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[matcher.scala 103:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[matcher.scala 103:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[matcher.scala 103:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[matcher.scala 103:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[matcher.scala 103:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[matcher.scala 103:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[matcher.scala 103:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[matcher.scala 103:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[matcher.scala 103:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[matcher.scala 103:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[matcher.scala 103:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[matcher.scala 103:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[matcher.scala 103:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[matcher.scala 103:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[matcher.scala 103:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[matcher.scala 103:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[matcher.scala 103:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[matcher.scala 103:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[matcher.scala 103:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[matcher.scala 103:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[matcher.scala 103:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[matcher.scala 103:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[matcher.scala 103:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[matcher.scala 103:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[matcher.scala 103:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[matcher.scala 103:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[matcher.scala 103:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[matcher.scala 103:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[matcher.scala 103:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[matcher.scala 103:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[matcher.scala 103:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[matcher.scala 103:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[matcher.scala 103:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[matcher.scala 103:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[matcher.scala 103:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[matcher.scala 103:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[matcher.scala 103:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[matcher.scala 103:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[matcher.scala 103:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[matcher.scala 103:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[matcher.scala 103:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[matcher.scala 103:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[matcher.scala 103:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[matcher.scala 103:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[matcher.scala 103:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[matcher.scala 103:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[matcher.scala 103:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[matcher.scala 103:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[matcher.scala 103:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[matcher.scala 103:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[matcher.scala 103:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[matcher.scala 103:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[matcher.scala 103:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[matcher.scala 103:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[matcher.scala 103:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[matcher.scala 103:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[matcher.scala 103:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[matcher.scala 103:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[matcher.scala 103:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[matcher.scala 103:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[matcher.scala 103:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[matcher.scala 103:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[matcher.scala 103:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[matcher.scala 103:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[matcher.scala 103:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[matcher.scala 103:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[matcher.scala 103:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[matcher.scala 103:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[matcher.scala 103:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[matcher.scala 103:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[matcher.scala 103:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[matcher.scala 103:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[matcher.scala 103:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[matcher.scala 103:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[matcher.scala 103:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[matcher.scala 103:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[matcher.scala 103:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[matcher.scala 103:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[matcher.scala 103:13]
    key <= io_key_in; // @[matcher.scala 107:13]
    addr <= io_addr_in; // @[matcher.scala 111:14]
    cs <= io_cs_in; // @[matcher.scala 115:12]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  phv_next_config_id = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_117[0:0];
  _RAND_118 = {2{`RANDOM}};
  key = _RAND_118[63:0];
  _RAND_119 = {1{`RANDOM}};
  addr = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  cs = _RAND_120[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MatchReadData(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input  [63:0] io_key_in,
  output [63:0] io_key_out,
  input  [2:0]  io_cs_in,
  output [2:0]  io_cs_out,
  input  [7:0]  io_addr_in,
  input         io_cs_vec_in_0,
  input         io_cs_vec_in_1,
  input         io_cs_vec_in_2,
  input         io_cs_vec_in_3,
  input         io_cs_vec_in_4,
  input         io_cs_vec_in_5,
  input         io_cs_vec_in_6,
  input         io_cs_vec_in_7,
  output [63:0] io_data_out_0,
  output [63:0] io_data_out_1,
  output [63:0] io_data_out_2,
  output [63:0] io_data_out_3,
  output [63:0] io_data_out_4,
  output [63:0] io_data_out_5,
  output [63:0] io_data_out_6,
  output [63:0] io_data_out_7,
  output        io_mem_cluster_0_en,
  output [7:0]  io_mem_cluster_0_addr,
  input  [63:0] io_mem_cluster_0_data,
  output        io_mem_cluster_1_en,
  output [7:0]  io_mem_cluster_1_addr,
  input  [63:0] io_mem_cluster_1_data,
  output        io_mem_cluster_2_en,
  output [7:0]  io_mem_cluster_2_addr,
  input  [63:0] io_mem_cluster_2_data,
  output        io_mem_cluster_3_en,
  output [7:0]  io_mem_cluster_3_addr,
  input  [63:0] io_mem_cluster_3_data,
  output        io_mem_cluster_4_en,
  output [7:0]  io_mem_cluster_4_addr,
  input  [63:0] io_mem_cluster_4_data,
  output        io_mem_cluster_5_en,
  output [7:0]  io_mem_cluster_5_addr,
  input  [63:0] io_mem_cluster_5_data,
  output        io_mem_cluster_6_en,
  output [7:0]  io_mem_cluster_6_addr,
  input  [63:0] io_mem_cluster_6_data,
  output        io_mem_cluster_7_en,
  output [7:0]  io_mem_cluster_7_addr,
  input  [63:0] io_mem_cluster_7_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [31:0] _RAND_119;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[matcher.scala 148:22]
  reg [7:0] phv_data_1; // @[matcher.scala 148:22]
  reg [7:0] phv_data_2; // @[matcher.scala 148:22]
  reg [7:0] phv_data_3; // @[matcher.scala 148:22]
  reg [7:0] phv_data_4; // @[matcher.scala 148:22]
  reg [7:0] phv_data_5; // @[matcher.scala 148:22]
  reg [7:0] phv_data_6; // @[matcher.scala 148:22]
  reg [7:0] phv_data_7; // @[matcher.scala 148:22]
  reg [7:0] phv_data_8; // @[matcher.scala 148:22]
  reg [7:0] phv_data_9; // @[matcher.scala 148:22]
  reg [7:0] phv_data_10; // @[matcher.scala 148:22]
  reg [7:0] phv_data_11; // @[matcher.scala 148:22]
  reg [7:0] phv_data_12; // @[matcher.scala 148:22]
  reg [7:0] phv_data_13; // @[matcher.scala 148:22]
  reg [7:0] phv_data_14; // @[matcher.scala 148:22]
  reg [7:0] phv_data_15; // @[matcher.scala 148:22]
  reg [7:0] phv_data_16; // @[matcher.scala 148:22]
  reg [7:0] phv_data_17; // @[matcher.scala 148:22]
  reg [7:0] phv_data_18; // @[matcher.scala 148:22]
  reg [7:0] phv_data_19; // @[matcher.scala 148:22]
  reg [7:0] phv_data_20; // @[matcher.scala 148:22]
  reg [7:0] phv_data_21; // @[matcher.scala 148:22]
  reg [7:0] phv_data_22; // @[matcher.scala 148:22]
  reg [7:0] phv_data_23; // @[matcher.scala 148:22]
  reg [7:0] phv_data_24; // @[matcher.scala 148:22]
  reg [7:0] phv_data_25; // @[matcher.scala 148:22]
  reg [7:0] phv_data_26; // @[matcher.scala 148:22]
  reg [7:0] phv_data_27; // @[matcher.scala 148:22]
  reg [7:0] phv_data_28; // @[matcher.scala 148:22]
  reg [7:0] phv_data_29; // @[matcher.scala 148:22]
  reg [7:0] phv_data_30; // @[matcher.scala 148:22]
  reg [7:0] phv_data_31; // @[matcher.scala 148:22]
  reg [7:0] phv_data_32; // @[matcher.scala 148:22]
  reg [7:0] phv_data_33; // @[matcher.scala 148:22]
  reg [7:0] phv_data_34; // @[matcher.scala 148:22]
  reg [7:0] phv_data_35; // @[matcher.scala 148:22]
  reg [7:0] phv_data_36; // @[matcher.scala 148:22]
  reg [7:0] phv_data_37; // @[matcher.scala 148:22]
  reg [7:0] phv_data_38; // @[matcher.scala 148:22]
  reg [7:0] phv_data_39; // @[matcher.scala 148:22]
  reg [7:0] phv_data_40; // @[matcher.scala 148:22]
  reg [7:0] phv_data_41; // @[matcher.scala 148:22]
  reg [7:0] phv_data_42; // @[matcher.scala 148:22]
  reg [7:0] phv_data_43; // @[matcher.scala 148:22]
  reg [7:0] phv_data_44; // @[matcher.scala 148:22]
  reg [7:0] phv_data_45; // @[matcher.scala 148:22]
  reg [7:0] phv_data_46; // @[matcher.scala 148:22]
  reg [7:0] phv_data_47; // @[matcher.scala 148:22]
  reg [7:0] phv_data_48; // @[matcher.scala 148:22]
  reg [7:0] phv_data_49; // @[matcher.scala 148:22]
  reg [7:0] phv_data_50; // @[matcher.scala 148:22]
  reg [7:0] phv_data_51; // @[matcher.scala 148:22]
  reg [7:0] phv_data_52; // @[matcher.scala 148:22]
  reg [7:0] phv_data_53; // @[matcher.scala 148:22]
  reg [7:0] phv_data_54; // @[matcher.scala 148:22]
  reg [7:0] phv_data_55; // @[matcher.scala 148:22]
  reg [7:0] phv_data_56; // @[matcher.scala 148:22]
  reg [7:0] phv_data_57; // @[matcher.scala 148:22]
  reg [7:0] phv_data_58; // @[matcher.scala 148:22]
  reg [7:0] phv_data_59; // @[matcher.scala 148:22]
  reg [7:0] phv_data_60; // @[matcher.scala 148:22]
  reg [7:0] phv_data_61; // @[matcher.scala 148:22]
  reg [7:0] phv_data_62; // @[matcher.scala 148:22]
  reg [7:0] phv_data_63; // @[matcher.scala 148:22]
  reg [7:0] phv_data_64; // @[matcher.scala 148:22]
  reg [7:0] phv_data_65; // @[matcher.scala 148:22]
  reg [7:0] phv_data_66; // @[matcher.scala 148:22]
  reg [7:0] phv_data_67; // @[matcher.scala 148:22]
  reg [7:0] phv_data_68; // @[matcher.scala 148:22]
  reg [7:0] phv_data_69; // @[matcher.scala 148:22]
  reg [7:0] phv_data_70; // @[matcher.scala 148:22]
  reg [7:0] phv_data_71; // @[matcher.scala 148:22]
  reg [7:0] phv_data_72; // @[matcher.scala 148:22]
  reg [7:0] phv_data_73; // @[matcher.scala 148:22]
  reg [7:0] phv_data_74; // @[matcher.scala 148:22]
  reg [7:0] phv_data_75; // @[matcher.scala 148:22]
  reg [7:0] phv_data_76; // @[matcher.scala 148:22]
  reg [7:0] phv_data_77; // @[matcher.scala 148:22]
  reg [7:0] phv_data_78; // @[matcher.scala 148:22]
  reg [7:0] phv_data_79; // @[matcher.scala 148:22]
  reg [7:0] phv_data_80; // @[matcher.scala 148:22]
  reg [7:0] phv_data_81; // @[matcher.scala 148:22]
  reg [7:0] phv_data_82; // @[matcher.scala 148:22]
  reg [7:0] phv_data_83; // @[matcher.scala 148:22]
  reg [7:0] phv_data_84; // @[matcher.scala 148:22]
  reg [7:0] phv_data_85; // @[matcher.scala 148:22]
  reg [7:0] phv_data_86; // @[matcher.scala 148:22]
  reg [7:0] phv_data_87; // @[matcher.scala 148:22]
  reg [7:0] phv_data_88; // @[matcher.scala 148:22]
  reg [7:0] phv_data_89; // @[matcher.scala 148:22]
  reg [7:0] phv_data_90; // @[matcher.scala 148:22]
  reg [7:0] phv_data_91; // @[matcher.scala 148:22]
  reg [7:0] phv_data_92; // @[matcher.scala 148:22]
  reg [7:0] phv_data_93; // @[matcher.scala 148:22]
  reg [7:0] phv_data_94; // @[matcher.scala 148:22]
  reg [7:0] phv_data_95; // @[matcher.scala 148:22]
  reg [15:0] phv_header_0; // @[matcher.scala 148:22]
  reg [15:0] phv_header_1; // @[matcher.scala 148:22]
  reg [15:0] phv_header_2; // @[matcher.scala 148:22]
  reg [15:0] phv_header_3; // @[matcher.scala 148:22]
  reg [15:0] phv_header_4; // @[matcher.scala 148:22]
  reg [15:0] phv_header_5; // @[matcher.scala 148:22]
  reg [15:0] phv_header_6; // @[matcher.scala 148:22]
  reg [15:0] phv_header_7; // @[matcher.scala 148:22]
  reg [15:0] phv_header_8; // @[matcher.scala 148:22]
  reg [15:0] phv_header_9; // @[matcher.scala 148:22]
  reg [15:0] phv_header_10; // @[matcher.scala 148:22]
  reg [15:0] phv_header_11; // @[matcher.scala 148:22]
  reg [15:0] phv_header_12; // @[matcher.scala 148:22]
  reg [15:0] phv_header_13; // @[matcher.scala 148:22]
  reg [15:0] phv_header_14; // @[matcher.scala 148:22]
  reg [15:0] phv_header_15; // @[matcher.scala 148:22]
  reg [7:0] phv_parse_current_state; // @[matcher.scala 148:22]
  reg [7:0] phv_parse_current_offset; // @[matcher.scala 148:22]
  reg [15:0] phv_parse_transition_field; // @[matcher.scala 148:22]
  reg [1:0] phv_next_processor_id; // @[matcher.scala 148:22]
  reg  phv_next_config_id; // @[matcher.scala 148:22]
  reg  phv_is_valid_processor; // @[matcher.scala 148:22]
  reg [63:0] key; // @[matcher.scala 152:22]
  reg [2:0] cs; // @[matcher.scala 156:21]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[matcher.scala 150:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[matcher.scala 150:25]
  assign io_key_out = key; // @[matcher.scala 154:20]
  assign io_cs_out = cs; // @[matcher.scala 158:19]
  assign io_data_out_0 = io_mem_cluster_0_data; // @[matcher.scala 163:36]
  assign io_data_out_1 = io_mem_cluster_1_data; // @[matcher.scala 163:36]
  assign io_data_out_2 = io_mem_cluster_2_data; // @[matcher.scala 163:36]
  assign io_data_out_3 = io_mem_cluster_3_data; // @[matcher.scala 163:36]
  assign io_data_out_4 = io_mem_cluster_4_data; // @[matcher.scala 163:36]
  assign io_data_out_5 = io_mem_cluster_5_data; // @[matcher.scala 163:36]
  assign io_data_out_6 = io_mem_cluster_6_data; // @[matcher.scala 163:36]
  assign io_data_out_7 = io_mem_cluster_7_data; // @[matcher.scala 163:36]
  assign io_mem_cluster_0_en = io_cs_vec_in_0 & io_pipe_phv_in_is_valid_processor; // @[matcher.scala 161:55]
  assign io_mem_cluster_0_addr = io_addr_in; // @[matcher.scala 162:36]
  assign io_mem_cluster_1_en = io_cs_vec_in_1 & io_pipe_phv_in_is_valid_processor; // @[matcher.scala 161:55]
  assign io_mem_cluster_1_addr = io_addr_in; // @[matcher.scala 162:36]
  assign io_mem_cluster_2_en = io_cs_vec_in_2 & io_pipe_phv_in_is_valid_processor; // @[matcher.scala 161:55]
  assign io_mem_cluster_2_addr = io_addr_in; // @[matcher.scala 162:36]
  assign io_mem_cluster_3_en = io_cs_vec_in_3 & io_pipe_phv_in_is_valid_processor; // @[matcher.scala 161:55]
  assign io_mem_cluster_3_addr = io_addr_in; // @[matcher.scala 162:36]
  assign io_mem_cluster_4_en = io_cs_vec_in_4 & io_pipe_phv_in_is_valid_processor; // @[matcher.scala 161:55]
  assign io_mem_cluster_4_addr = io_addr_in; // @[matcher.scala 162:36]
  assign io_mem_cluster_5_en = io_cs_vec_in_5 & io_pipe_phv_in_is_valid_processor; // @[matcher.scala 161:55]
  assign io_mem_cluster_5_addr = io_addr_in; // @[matcher.scala 162:36]
  assign io_mem_cluster_6_en = io_cs_vec_in_6 & io_pipe_phv_in_is_valid_processor; // @[matcher.scala 161:55]
  assign io_mem_cluster_6_addr = io_addr_in; // @[matcher.scala 162:36]
  assign io_mem_cluster_7_en = io_cs_vec_in_7 & io_pipe_phv_in_is_valid_processor; // @[matcher.scala 161:55]
  assign io_mem_cluster_7_addr = io_addr_in; // @[matcher.scala 162:36]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[matcher.scala 149:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[matcher.scala 149:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[matcher.scala 149:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[matcher.scala 149:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[matcher.scala 149:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[matcher.scala 149:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[matcher.scala 149:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[matcher.scala 149:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[matcher.scala 149:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[matcher.scala 149:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[matcher.scala 149:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[matcher.scala 149:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[matcher.scala 149:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[matcher.scala 149:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[matcher.scala 149:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[matcher.scala 149:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[matcher.scala 149:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[matcher.scala 149:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[matcher.scala 149:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[matcher.scala 149:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[matcher.scala 149:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[matcher.scala 149:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[matcher.scala 149:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[matcher.scala 149:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[matcher.scala 149:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[matcher.scala 149:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[matcher.scala 149:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[matcher.scala 149:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[matcher.scala 149:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[matcher.scala 149:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[matcher.scala 149:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[matcher.scala 149:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[matcher.scala 149:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[matcher.scala 149:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[matcher.scala 149:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[matcher.scala 149:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[matcher.scala 149:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[matcher.scala 149:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[matcher.scala 149:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[matcher.scala 149:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[matcher.scala 149:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[matcher.scala 149:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[matcher.scala 149:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[matcher.scala 149:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[matcher.scala 149:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[matcher.scala 149:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[matcher.scala 149:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[matcher.scala 149:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[matcher.scala 149:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[matcher.scala 149:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[matcher.scala 149:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[matcher.scala 149:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[matcher.scala 149:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[matcher.scala 149:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[matcher.scala 149:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[matcher.scala 149:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[matcher.scala 149:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[matcher.scala 149:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[matcher.scala 149:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[matcher.scala 149:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[matcher.scala 149:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[matcher.scala 149:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[matcher.scala 149:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[matcher.scala 149:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[matcher.scala 149:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[matcher.scala 149:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[matcher.scala 149:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[matcher.scala 149:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[matcher.scala 149:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[matcher.scala 149:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[matcher.scala 149:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[matcher.scala 149:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[matcher.scala 149:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[matcher.scala 149:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[matcher.scala 149:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[matcher.scala 149:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[matcher.scala 149:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[matcher.scala 149:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[matcher.scala 149:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[matcher.scala 149:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[matcher.scala 149:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[matcher.scala 149:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[matcher.scala 149:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[matcher.scala 149:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[matcher.scala 149:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[matcher.scala 149:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[matcher.scala 149:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[matcher.scala 149:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[matcher.scala 149:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[matcher.scala 149:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[matcher.scala 149:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[matcher.scala 149:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[matcher.scala 149:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[matcher.scala 149:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[matcher.scala 149:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[matcher.scala 149:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[matcher.scala 149:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[matcher.scala 149:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[matcher.scala 149:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[matcher.scala 149:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[matcher.scala 149:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[matcher.scala 149:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[matcher.scala 149:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[matcher.scala 149:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[matcher.scala 149:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[matcher.scala 149:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[matcher.scala 149:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[matcher.scala 149:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[matcher.scala 149:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[matcher.scala 149:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[matcher.scala 149:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[matcher.scala 149:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[matcher.scala 149:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[matcher.scala 149:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[matcher.scala 149:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[matcher.scala 149:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[matcher.scala 149:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[matcher.scala 149:13]
    key <= io_key_in; // @[matcher.scala 153:13]
    cs <= io_cs_in; // @[matcher.scala 157:12]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  phv_next_config_id = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_117[0:0];
  _RAND_118 = {2{`RANDOM}};
  key = _RAND_118[63:0];
  _RAND_119 = {1{`RANDOM}};
  cs = _RAND_119[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MatchDataReshape(
  input          clock,
  input  [7:0]   io_pipe_phv_in_data_0,
  input  [7:0]   io_pipe_phv_in_data_1,
  input  [7:0]   io_pipe_phv_in_data_2,
  input  [7:0]   io_pipe_phv_in_data_3,
  input  [7:0]   io_pipe_phv_in_data_4,
  input  [7:0]   io_pipe_phv_in_data_5,
  input  [7:0]   io_pipe_phv_in_data_6,
  input  [7:0]   io_pipe_phv_in_data_7,
  input  [7:0]   io_pipe_phv_in_data_8,
  input  [7:0]   io_pipe_phv_in_data_9,
  input  [7:0]   io_pipe_phv_in_data_10,
  input  [7:0]   io_pipe_phv_in_data_11,
  input  [7:0]   io_pipe_phv_in_data_12,
  input  [7:0]   io_pipe_phv_in_data_13,
  input  [7:0]   io_pipe_phv_in_data_14,
  input  [7:0]   io_pipe_phv_in_data_15,
  input  [7:0]   io_pipe_phv_in_data_16,
  input  [7:0]   io_pipe_phv_in_data_17,
  input  [7:0]   io_pipe_phv_in_data_18,
  input  [7:0]   io_pipe_phv_in_data_19,
  input  [7:0]   io_pipe_phv_in_data_20,
  input  [7:0]   io_pipe_phv_in_data_21,
  input  [7:0]   io_pipe_phv_in_data_22,
  input  [7:0]   io_pipe_phv_in_data_23,
  input  [7:0]   io_pipe_phv_in_data_24,
  input  [7:0]   io_pipe_phv_in_data_25,
  input  [7:0]   io_pipe_phv_in_data_26,
  input  [7:0]   io_pipe_phv_in_data_27,
  input  [7:0]   io_pipe_phv_in_data_28,
  input  [7:0]   io_pipe_phv_in_data_29,
  input  [7:0]   io_pipe_phv_in_data_30,
  input  [7:0]   io_pipe_phv_in_data_31,
  input  [7:0]   io_pipe_phv_in_data_32,
  input  [7:0]   io_pipe_phv_in_data_33,
  input  [7:0]   io_pipe_phv_in_data_34,
  input  [7:0]   io_pipe_phv_in_data_35,
  input  [7:0]   io_pipe_phv_in_data_36,
  input  [7:0]   io_pipe_phv_in_data_37,
  input  [7:0]   io_pipe_phv_in_data_38,
  input  [7:0]   io_pipe_phv_in_data_39,
  input  [7:0]   io_pipe_phv_in_data_40,
  input  [7:0]   io_pipe_phv_in_data_41,
  input  [7:0]   io_pipe_phv_in_data_42,
  input  [7:0]   io_pipe_phv_in_data_43,
  input  [7:0]   io_pipe_phv_in_data_44,
  input  [7:0]   io_pipe_phv_in_data_45,
  input  [7:0]   io_pipe_phv_in_data_46,
  input  [7:0]   io_pipe_phv_in_data_47,
  input  [7:0]   io_pipe_phv_in_data_48,
  input  [7:0]   io_pipe_phv_in_data_49,
  input  [7:0]   io_pipe_phv_in_data_50,
  input  [7:0]   io_pipe_phv_in_data_51,
  input  [7:0]   io_pipe_phv_in_data_52,
  input  [7:0]   io_pipe_phv_in_data_53,
  input  [7:0]   io_pipe_phv_in_data_54,
  input  [7:0]   io_pipe_phv_in_data_55,
  input  [7:0]   io_pipe_phv_in_data_56,
  input  [7:0]   io_pipe_phv_in_data_57,
  input  [7:0]   io_pipe_phv_in_data_58,
  input  [7:0]   io_pipe_phv_in_data_59,
  input  [7:0]   io_pipe_phv_in_data_60,
  input  [7:0]   io_pipe_phv_in_data_61,
  input  [7:0]   io_pipe_phv_in_data_62,
  input  [7:0]   io_pipe_phv_in_data_63,
  input  [7:0]   io_pipe_phv_in_data_64,
  input  [7:0]   io_pipe_phv_in_data_65,
  input  [7:0]   io_pipe_phv_in_data_66,
  input  [7:0]   io_pipe_phv_in_data_67,
  input  [7:0]   io_pipe_phv_in_data_68,
  input  [7:0]   io_pipe_phv_in_data_69,
  input  [7:0]   io_pipe_phv_in_data_70,
  input  [7:0]   io_pipe_phv_in_data_71,
  input  [7:0]   io_pipe_phv_in_data_72,
  input  [7:0]   io_pipe_phv_in_data_73,
  input  [7:0]   io_pipe_phv_in_data_74,
  input  [7:0]   io_pipe_phv_in_data_75,
  input  [7:0]   io_pipe_phv_in_data_76,
  input  [7:0]   io_pipe_phv_in_data_77,
  input  [7:0]   io_pipe_phv_in_data_78,
  input  [7:0]   io_pipe_phv_in_data_79,
  input  [7:0]   io_pipe_phv_in_data_80,
  input  [7:0]   io_pipe_phv_in_data_81,
  input  [7:0]   io_pipe_phv_in_data_82,
  input  [7:0]   io_pipe_phv_in_data_83,
  input  [7:0]   io_pipe_phv_in_data_84,
  input  [7:0]   io_pipe_phv_in_data_85,
  input  [7:0]   io_pipe_phv_in_data_86,
  input  [7:0]   io_pipe_phv_in_data_87,
  input  [7:0]   io_pipe_phv_in_data_88,
  input  [7:0]   io_pipe_phv_in_data_89,
  input  [7:0]   io_pipe_phv_in_data_90,
  input  [7:0]   io_pipe_phv_in_data_91,
  input  [7:0]   io_pipe_phv_in_data_92,
  input  [7:0]   io_pipe_phv_in_data_93,
  input  [7:0]   io_pipe_phv_in_data_94,
  input  [7:0]   io_pipe_phv_in_data_95,
  input  [15:0]  io_pipe_phv_in_header_0,
  input  [15:0]  io_pipe_phv_in_header_1,
  input  [15:0]  io_pipe_phv_in_header_2,
  input  [15:0]  io_pipe_phv_in_header_3,
  input  [15:0]  io_pipe_phv_in_header_4,
  input  [15:0]  io_pipe_phv_in_header_5,
  input  [15:0]  io_pipe_phv_in_header_6,
  input  [15:0]  io_pipe_phv_in_header_7,
  input  [15:0]  io_pipe_phv_in_header_8,
  input  [15:0]  io_pipe_phv_in_header_9,
  input  [15:0]  io_pipe_phv_in_header_10,
  input  [15:0]  io_pipe_phv_in_header_11,
  input  [15:0]  io_pipe_phv_in_header_12,
  input  [15:0]  io_pipe_phv_in_header_13,
  input  [15:0]  io_pipe_phv_in_header_14,
  input  [15:0]  io_pipe_phv_in_header_15,
  input  [7:0]   io_pipe_phv_in_parse_current_state,
  input  [7:0]   io_pipe_phv_in_parse_current_offset,
  input  [15:0]  io_pipe_phv_in_parse_transition_field,
  input  [1:0]   io_pipe_phv_in_next_processor_id,
  input          io_pipe_phv_in_next_config_id,
  input          io_pipe_phv_in_is_valid_processor,
  output [7:0]   io_pipe_phv_out_data_0,
  output [7:0]   io_pipe_phv_out_data_1,
  output [7:0]   io_pipe_phv_out_data_2,
  output [7:0]   io_pipe_phv_out_data_3,
  output [7:0]   io_pipe_phv_out_data_4,
  output [7:0]   io_pipe_phv_out_data_5,
  output [7:0]   io_pipe_phv_out_data_6,
  output [7:0]   io_pipe_phv_out_data_7,
  output [7:0]   io_pipe_phv_out_data_8,
  output [7:0]   io_pipe_phv_out_data_9,
  output [7:0]   io_pipe_phv_out_data_10,
  output [7:0]   io_pipe_phv_out_data_11,
  output [7:0]   io_pipe_phv_out_data_12,
  output [7:0]   io_pipe_phv_out_data_13,
  output [7:0]   io_pipe_phv_out_data_14,
  output [7:0]   io_pipe_phv_out_data_15,
  output [7:0]   io_pipe_phv_out_data_16,
  output [7:0]   io_pipe_phv_out_data_17,
  output [7:0]   io_pipe_phv_out_data_18,
  output [7:0]   io_pipe_phv_out_data_19,
  output [7:0]   io_pipe_phv_out_data_20,
  output [7:0]   io_pipe_phv_out_data_21,
  output [7:0]   io_pipe_phv_out_data_22,
  output [7:0]   io_pipe_phv_out_data_23,
  output [7:0]   io_pipe_phv_out_data_24,
  output [7:0]   io_pipe_phv_out_data_25,
  output [7:0]   io_pipe_phv_out_data_26,
  output [7:0]   io_pipe_phv_out_data_27,
  output [7:0]   io_pipe_phv_out_data_28,
  output [7:0]   io_pipe_phv_out_data_29,
  output [7:0]   io_pipe_phv_out_data_30,
  output [7:0]   io_pipe_phv_out_data_31,
  output [7:0]   io_pipe_phv_out_data_32,
  output [7:0]   io_pipe_phv_out_data_33,
  output [7:0]   io_pipe_phv_out_data_34,
  output [7:0]   io_pipe_phv_out_data_35,
  output [7:0]   io_pipe_phv_out_data_36,
  output [7:0]   io_pipe_phv_out_data_37,
  output [7:0]   io_pipe_phv_out_data_38,
  output [7:0]   io_pipe_phv_out_data_39,
  output [7:0]   io_pipe_phv_out_data_40,
  output [7:0]   io_pipe_phv_out_data_41,
  output [7:0]   io_pipe_phv_out_data_42,
  output [7:0]   io_pipe_phv_out_data_43,
  output [7:0]   io_pipe_phv_out_data_44,
  output [7:0]   io_pipe_phv_out_data_45,
  output [7:0]   io_pipe_phv_out_data_46,
  output [7:0]   io_pipe_phv_out_data_47,
  output [7:0]   io_pipe_phv_out_data_48,
  output [7:0]   io_pipe_phv_out_data_49,
  output [7:0]   io_pipe_phv_out_data_50,
  output [7:0]   io_pipe_phv_out_data_51,
  output [7:0]   io_pipe_phv_out_data_52,
  output [7:0]   io_pipe_phv_out_data_53,
  output [7:0]   io_pipe_phv_out_data_54,
  output [7:0]   io_pipe_phv_out_data_55,
  output [7:0]   io_pipe_phv_out_data_56,
  output [7:0]   io_pipe_phv_out_data_57,
  output [7:0]   io_pipe_phv_out_data_58,
  output [7:0]   io_pipe_phv_out_data_59,
  output [7:0]   io_pipe_phv_out_data_60,
  output [7:0]   io_pipe_phv_out_data_61,
  output [7:0]   io_pipe_phv_out_data_62,
  output [7:0]   io_pipe_phv_out_data_63,
  output [7:0]   io_pipe_phv_out_data_64,
  output [7:0]   io_pipe_phv_out_data_65,
  output [7:0]   io_pipe_phv_out_data_66,
  output [7:0]   io_pipe_phv_out_data_67,
  output [7:0]   io_pipe_phv_out_data_68,
  output [7:0]   io_pipe_phv_out_data_69,
  output [7:0]   io_pipe_phv_out_data_70,
  output [7:0]   io_pipe_phv_out_data_71,
  output [7:0]   io_pipe_phv_out_data_72,
  output [7:0]   io_pipe_phv_out_data_73,
  output [7:0]   io_pipe_phv_out_data_74,
  output [7:0]   io_pipe_phv_out_data_75,
  output [7:0]   io_pipe_phv_out_data_76,
  output [7:0]   io_pipe_phv_out_data_77,
  output [7:0]   io_pipe_phv_out_data_78,
  output [7:0]   io_pipe_phv_out_data_79,
  output [7:0]   io_pipe_phv_out_data_80,
  output [7:0]   io_pipe_phv_out_data_81,
  output [7:0]   io_pipe_phv_out_data_82,
  output [7:0]   io_pipe_phv_out_data_83,
  output [7:0]   io_pipe_phv_out_data_84,
  output [7:0]   io_pipe_phv_out_data_85,
  output [7:0]   io_pipe_phv_out_data_86,
  output [7:0]   io_pipe_phv_out_data_87,
  output [7:0]   io_pipe_phv_out_data_88,
  output [7:0]   io_pipe_phv_out_data_89,
  output [7:0]   io_pipe_phv_out_data_90,
  output [7:0]   io_pipe_phv_out_data_91,
  output [7:0]   io_pipe_phv_out_data_92,
  output [7:0]   io_pipe_phv_out_data_93,
  output [7:0]   io_pipe_phv_out_data_94,
  output [7:0]   io_pipe_phv_out_data_95,
  output [15:0]  io_pipe_phv_out_header_0,
  output [15:0]  io_pipe_phv_out_header_1,
  output [15:0]  io_pipe_phv_out_header_2,
  output [15:0]  io_pipe_phv_out_header_3,
  output [15:0]  io_pipe_phv_out_header_4,
  output [15:0]  io_pipe_phv_out_header_5,
  output [15:0]  io_pipe_phv_out_header_6,
  output [15:0]  io_pipe_phv_out_header_7,
  output [15:0]  io_pipe_phv_out_header_8,
  output [15:0]  io_pipe_phv_out_header_9,
  output [15:0]  io_pipe_phv_out_header_10,
  output [15:0]  io_pipe_phv_out_header_11,
  output [15:0]  io_pipe_phv_out_header_12,
  output [15:0]  io_pipe_phv_out_header_13,
  output [15:0]  io_pipe_phv_out_header_14,
  output [15:0]  io_pipe_phv_out_header_15,
  output [7:0]   io_pipe_phv_out_parse_current_state,
  output [7:0]   io_pipe_phv_out_parse_current_offset,
  output [15:0]  io_pipe_phv_out_parse_transition_field,
  output [1:0]   io_pipe_phv_out_next_processor_id,
  output         io_pipe_phv_out_next_config_id,
  output         io_pipe_phv_out_is_valid_processor,
  input  [3:0]   io_table_config_0_table_width,
  input  [3:0]   io_table_config_0_table_depth,
  input  [3:0]   io_table_config_1_table_width,
  input  [3:0]   io_table_config_1_table_depth,
  input  [63:0]  io_key_in,
  output [63:0]  io_key_out,
  input  [2:0]   io_cs_in,
  input  [63:0]  io_data_in_0,
  input  [63:0]  io_data_in_1,
  input  [63:0]  io_data_in_2,
  input  [63:0]  io_data_in_3,
  input  [63:0]  io_data_in_4,
  input  [63:0]  io_data_in_5,
  input  [63:0]  io_data_in_6,
  input  [63:0]  io_data_in_7,
  output [127:0] io_data_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [127:0] _RAND_119;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[matcher.scala 180:22]
  reg [7:0] phv_data_1; // @[matcher.scala 180:22]
  reg [7:0] phv_data_2; // @[matcher.scala 180:22]
  reg [7:0] phv_data_3; // @[matcher.scala 180:22]
  reg [7:0] phv_data_4; // @[matcher.scala 180:22]
  reg [7:0] phv_data_5; // @[matcher.scala 180:22]
  reg [7:0] phv_data_6; // @[matcher.scala 180:22]
  reg [7:0] phv_data_7; // @[matcher.scala 180:22]
  reg [7:0] phv_data_8; // @[matcher.scala 180:22]
  reg [7:0] phv_data_9; // @[matcher.scala 180:22]
  reg [7:0] phv_data_10; // @[matcher.scala 180:22]
  reg [7:0] phv_data_11; // @[matcher.scala 180:22]
  reg [7:0] phv_data_12; // @[matcher.scala 180:22]
  reg [7:0] phv_data_13; // @[matcher.scala 180:22]
  reg [7:0] phv_data_14; // @[matcher.scala 180:22]
  reg [7:0] phv_data_15; // @[matcher.scala 180:22]
  reg [7:0] phv_data_16; // @[matcher.scala 180:22]
  reg [7:0] phv_data_17; // @[matcher.scala 180:22]
  reg [7:0] phv_data_18; // @[matcher.scala 180:22]
  reg [7:0] phv_data_19; // @[matcher.scala 180:22]
  reg [7:0] phv_data_20; // @[matcher.scala 180:22]
  reg [7:0] phv_data_21; // @[matcher.scala 180:22]
  reg [7:0] phv_data_22; // @[matcher.scala 180:22]
  reg [7:0] phv_data_23; // @[matcher.scala 180:22]
  reg [7:0] phv_data_24; // @[matcher.scala 180:22]
  reg [7:0] phv_data_25; // @[matcher.scala 180:22]
  reg [7:0] phv_data_26; // @[matcher.scala 180:22]
  reg [7:0] phv_data_27; // @[matcher.scala 180:22]
  reg [7:0] phv_data_28; // @[matcher.scala 180:22]
  reg [7:0] phv_data_29; // @[matcher.scala 180:22]
  reg [7:0] phv_data_30; // @[matcher.scala 180:22]
  reg [7:0] phv_data_31; // @[matcher.scala 180:22]
  reg [7:0] phv_data_32; // @[matcher.scala 180:22]
  reg [7:0] phv_data_33; // @[matcher.scala 180:22]
  reg [7:0] phv_data_34; // @[matcher.scala 180:22]
  reg [7:0] phv_data_35; // @[matcher.scala 180:22]
  reg [7:0] phv_data_36; // @[matcher.scala 180:22]
  reg [7:0] phv_data_37; // @[matcher.scala 180:22]
  reg [7:0] phv_data_38; // @[matcher.scala 180:22]
  reg [7:0] phv_data_39; // @[matcher.scala 180:22]
  reg [7:0] phv_data_40; // @[matcher.scala 180:22]
  reg [7:0] phv_data_41; // @[matcher.scala 180:22]
  reg [7:0] phv_data_42; // @[matcher.scala 180:22]
  reg [7:0] phv_data_43; // @[matcher.scala 180:22]
  reg [7:0] phv_data_44; // @[matcher.scala 180:22]
  reg [7:0] phv_data_45; // @[matcher.scala 180:22]
  reg [7:0] phv_data_46; // @[matcher.scala 180:22]
  reg [7:0] phv_data_47; // @[matcher.scala 180:22]
  reg [7:0] phv_data_48; // @[matcher.scala 180:22]
  reg [7:0] phv_data_49; // @[matcher.scala 180:22]
  reg [7:0] phv_data_50; // @[matcher.scala 180:22]
  reg [7:0] phv_data_51; // @[matcher.scala 180:22]
  reg [7:0] phv_data_52; // @[matcher.scala 180:22]
  reg [7:0] phv_data_53; // @[matcher.scala 180:22]
  reg [7:0] phv_data_54; // @[matcher.scala 180:22]
  reg [7:0] phv_data_55; // @[matcher.scala 180:22]
  reg [7:0] phv_data_56; // @[matcher.scala 180:22]
  reg [7:0] phv_data_57; // @[matcher.scala 180:22]
  reg [7:0] phv_data_58; // @[matcher.scala 180:22]
  reg [7:0] phv_data_59; // @[matcher.scala 180:22]
  reg [7:0] phv_data_60; // @[matcher.scala 180:22]
  reg [7:0] phv_data_61; // @[matcher.scala 180:22]
  reg [7:0] phv_data_62; // @[matcher.scala 180:22]
  reg [7:0] phv_data_63; // @[matcher.scala 180:22]
  reg [7:0] phv_data_64; // @[matcher.scala 180:22]
  reg [7:0] phv_data_65; // @[matcher.scala 180:22]
  reg [7:0] phv_data_66; // @[matcher.scala 180:22]
  reg [7:0] phv_data_67; // @[matcher.scala 180:22]
  reg [7:0] phv_data_68; // @[matcher.scala 180:22]
  reg [7:0] phv_data_69; // @[matcher.scala 180:22]
  reg [7:0] phv_data_70; // @[matcher.scala 180:22]
  reg [7:0] phv_data_71; // @[matcher.scala 180:22]
  reg [7:0] phv_data_72; // @[matcher.scala 180:22]
  reg [7:0] phv_data_73; // @[matcher.scala 180:22]
  reg [7:0] phv_data_74; // @[matcher.scala 180:22]
  reg [7:0] phv_data_75; // @[matcher.scala 180:22]
  reg [7:0] phv_data_76; // @[matcher.scala 180:22]
  reg [7:0] phv_data_77; // @[matcher.scala 180:22]
  reg [7:0] phv_data_78; // @[matcher.scala 180:22]
  reg [7:0] phv_data_79; // @[matcher.scala 180:22]
  reg [7:0] phv_data_80; // @[matcher.scala 180:22]
  reg [7:0] phv_data_81; // @[matcher.scala 180:22]
  reg [7:0] phv_data_82; // @[matcher.scala 180:22]
  reg [7:0] phv_data_83; // @[matcher.scala 180:22]
  reg [7:0] phv_data_84; // @[matcher.scala 180:22]
  reg [7:0] phv_data_85; // @[matcher.scala 180:22]
  reg [7:0] phv_data_86; // @[matcher.scala 180:22]
  reg [7:0] phv_data_87; // @[matcher.scala 180:22]
  reg [7:0] phv_data_88; // @[matcher.scala 180:22]
  reg [7:0] phv_data_89; // @[matcher.scala 180:22]
  reg [7:0] phv_data_90; // @[matcher.scala 180:22]
  reg [7:0] phv_data_91; // @[matcher.scala 180:22]
  reg [7:0] phv_data_92; // @[matcher.scala 180:22]
  reg [7:0] phv_data_93; // @[matcher.scala 180:22]
  reg [7:0] phv_data_94; // @[matcher.scala 180:22]
  reg [7:0] phv_data_95; // @[matcher.scala 180:22]
  reg [15:0] phv_header_0; // @[matcher.scala 180:22]
  reg [15:0] phv_header_1; // @[matcher.scala 180:22]
  reg [15:0] phv_header_2; // @[matcher.scala 180:22]
  reg [15:0] phv_header_3; // @[matcher.scala 180:22]
  reg [15:0] phv_header_4; // @[matcher.scala 180:22]
  reg [15:0] phv_header_5; // @[matcher.scala 180:22]
  reg [15:0] phv_header_6; // @[matcher.scala 180:22]
  reg [15:0] phv_header_7; // @[matcher.scala 180:22]
  reg [15:0] phv_header_8; // @[matcher.scala 180:22]
  reg [15:0] phv_header_9; // @[matcher.scala 180:22]
  reg [15:0] phv_header_10; // @[matcher.scala 180:22]
  reg [15:0] phv_header_11; // @[matcher.scala 180:22]
  reg [15:0] phv_header_12; // @[matcher.scala 180:22]
  reg [15:0] phv_header_13; // @[matcher.scala 180:22]
  reg [15:0] phv_header_14; // @[matcher.scala 180:22]
  reg [15:0] phv_header_15; // @[matcher.scala 180:22]
  reg [7:0] phv_parse_current_state; // @[matcher.scala 180:22]
  reg [7:0] phv_parse_current_offset; // @[matcher.scala 180:22]
  reg [15:0] phv_parse_transition_field; // @[matcher.scala 180:22]
  reg [1:0] phv_next_processor_id; // @[matcher.scala 180:22]
  reg  phv_next_config_id; // @[matcher.scala 180:22]
  reg  phv_is_valid_processor; // @[matcher.scala 180:22]
  reg [63:0] key; // @[matcher.scala 184:22]
  reg [127:0] data; // @[matcher.scala 188:23]
  wire [63:0] _GEN_0 = io_cs_in == 3'h0 ? io_data_in_0 : 64'h0; // @[matcher.scala 198:69 matcher.scala 199:27 matcher.scala 194:19]
  wire [3:0] _GEN_19 = io_pipe_phv_in_next_config_id ? io_table_config_1_table_width : io_table_config_0_table_width; // @[matcher.scala 201:61 matcher.scala 201:61]
  wire [3:0] _GEN_20 = io_pipe_phv_in_next_config_id ? io_table_config_1_table_depth : io_table_config_0_table_depth; // @[matcher.scala 201:61 matcher.scala 201:61]
  wire  width_extend = _GEN_19 == 4'h2; // @[matcher.scala 201:61]
  wire [3:0] _GEN_37 = {{1'd0}, io_cs_in}; // @[matcher.scala 202:48]
  wire [3:0] _T_2 = _GEN_37 + _GEN_20; // @[matcher.scala 202:48]
  wire [63:0] _GEN_21 = width_extend & _T_2 == 4'h0 ? io_data_in_0 : 64'h0; // @[matcher.scala 202:112 matcher.scala 203:27 matcher.scala 195:19]
  wire [63:0] _GEN_22 = io_cs_in == 3'h1 ? io_data_in_1 : _GEN_0; // @[matcher.scala 198:69 matcher.scala 199:27]
  wire [63:0] _GEN_23 = width_extend & _T_2 == 4'h1 ? io_data_in_1 : _GEN_21; // @[matcher.scala 202:112 matcher.scala 203:27]
  wire [63:0] _GEN_24 = io_cs_in == 3'h2 ? io_data_in_2 : _GEN_22; // @[matcher.scala 198:69 matcher.scala 199:27]
  wire [63:0] _GEN_25 = width_extend & _T_2 == 4'h2 ? io_data_in_2 : _GEN_23; // @[matcher.scala 202:112 matcher.scala 203:27]
  wire [63:0] _GEN_26 = io_cs_in == 3'h3 ? io_data_in_3 : _GEN_24; // @[matcher.scala 198:69 matcher.scala 199:27]
  wire [63:0] _GEN_27 = width_extend & _T_2 == 4'h3 ? io_data_in_3 : _GEN_25; // @[matcher.scala 202:112 matcher.scala 203:27]
  wire [63:0] _GEN_28 = io_cs_in == 3'h4 ? io_data_in_4 : _GEN_26; // @[matcher.scala 198:69 matcher.scala 199:27]
  wire [63:0] _GEN_29 = width_extend & _T_2 == 4'h4 ? io_data_in_4 : _GEN_27; // @[matcher.scala 202:112 matcher.scala 203:27]
  wire [63:0] _GEN_30 = io_cs_in == 3'h5 ? io_data_in_5 : _GEN_28; // @[matcher.scala 198:69 matcher.scala 199:27]
  wire [63:0] _GEN_31 = width_extend & _T_2 == 4'h5 ? io_data_in_5 : _GEN_29; // @[matcher.scala 202:112 matcher.scala 203:27]
  wire [63:0] _GEN_32 = io_cs_in == 3'h6 ? io_data_in_6 : _GEN_30; // @[matcher.scala 198:69 matcher.scala 199:27]
  wire [63:0] _GEN_33 = width_extend & _T_2 == 4'h6 ? io_data_in_6 : _GEN_31; // @[matcher.scala 202:112 matcher.scala 203:27]
  wire [63:0] data_hi = io_cs_in == 3'h7 ? io_data_in_7 : _GEN_32; // @[matcher.scala 198:69 matcher.scala 199:27]
  wire [63:0] data_lo = width_extend & _T_2 == 4'h7 ? io_data_in_7 : _GEN_33; // @[matcher.scala 202:112 matcher.scala 203:27]
  wire [127:0] _data_T = {data_hi,data_lo}; // @[Cat.scala 30:58]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[matcher.scala 182:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[matcher.scala 182:25]
  assign io_key_out = key; // @[matcher.scala 186:20]
  assign io_data_out = data; // @[matcher.scala 211:21]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[matcher.scala 181:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[matcher.scala 181:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[matcher.scala 181:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[matcher.scala 181:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[matcher.scala 181:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[matcher.scala 181:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[matcher.scala 181:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[matcher.scala 181:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[matcher.scala 181:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[matcher.scala 181:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[matcher.scala 181:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[matcher.scala 181:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[matcher.scala 181:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[matcher.scala 181:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[matcher.scala 181:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[matcher.scala 181:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[matcher.scala 181:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[matcher.scala 181:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[matcher.scala 181:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[matcher.scala 181:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[matcher.scala 181:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[matcher.scala 181:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[matcher.scala 181:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[matcher.scala 181:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[matcher.scala 181:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[matcher.scala 181:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[matcher.scala 181:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[matcher.scala 181:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[matcher.scala 181:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[matcher.scala 181:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[matcher.scala 181:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[matcher.scala 181:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[matcher.scala 181:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[matcher.scala 181:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[matcher.scala 181:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[matcher.scala 181:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[matcher.scala 181:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[matcher.scala 181:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[matcher.scala 181:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[matcher.scala 181:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[matcher.scala 181:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[matcher.scala 181:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[matcher.scala 181:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[matcher.scala 181:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[matcher.scala 181:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[matcher.scala 181:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[matcher.scala 181:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[matcher.scala 181:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[matcher.scala 181:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[matcher.scala 181:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[matcher.scala 181:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[matcher.scala 181:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[matcher.scala 181:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[matcher.scala 181:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[matcher.scala 181:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[matcher.scala 181:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[matcher.scala 181:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[matcher.scala 181:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[matcher.scala 181:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[matcher.scala 181:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[matcher.scala 181:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[matcher.scala 181:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[matcher.scala 181:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[matcher.scala 181:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[matcher.scala 181:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[matcher.scala 181:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[matcher.scala 181:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[matcher.scala 181:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[matcher.scala 181:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[matcher.scala 181:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[matcher.scala 181:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[matcher.scala 181:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[matcher.scala 181:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[matcher.scala 181:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[matcher.scala 181:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[matcher.scala 181:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[matcher.scala 181:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[matcher.scala 181:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[matcher.scala 181:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[matcher.scala 181:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[matcher.scala 181:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[matcher.scala 181:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[matcher.scala 181:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[matcher.scala 181:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[matcher.scala 181:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[matcher.scala 181:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[matcher.scala 181:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[matcher.scala 181:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[matcher.scala 181:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[matcher.scala 181:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[matcher.scala 181:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[matcher.scala 181:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[matcher.scala 181:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[matcher.scala 181:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[matcher.scala 181:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[matcher.scala 181:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[matcher.scala 181:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[matcher.scala 181:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[matcher.scala 181:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[matcher.scala 181:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[matcher.scala 181:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[matcher.scala 181:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[matcher.scala 181:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[matcher.scala 181:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[matcher.scala 181:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[matcher.scala 181:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[matcher.scala 181:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[matcher.scala 181:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[matcher.scala 181:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[matcher.scala 181:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[matcher.scala 181:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[matcher.scala 181:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[matcher.scala 181:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[matcher.scala 181:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[matcher.scala 181:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[matcher.scala 181:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[matcher.scala 181:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[matcher.scala 181:13]
    key <= io_key_in; // @[matcher.scala 185:13]
    if (io_pipe_phv_in_is_valid_processor) begin // @[matcher.scala 191:50]
      data <= _data_T; // @[matcher.scala 206:18]
    end else begin
      data <= 128'h0; // @[matcher.scala 208:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  phv_next_config_id = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_117[0:0];
  _RAND_118 = {2{`RANDOM}};
  key = _RAND_118[63:0];
  _RAND_119 = {4{`RANDOM}};
  data = _RAND_119[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MatchResult(
  input          clock,
  input  [7:0]   io_pipe_phv_in_data_0,
  input  [7:0]   io_pipe_phv_in_data_1,
  input  [7:0]   io_pipe_phv_in_data_2,
  input  [7:0]   io_pipe_phv_in_data_3,
  input  [7:0]   io_pipe_phv_in_data_4,
  input  [7:0]   io_pipe_phv_in_data_5,
  input  [7:0]   io_pipe_phv_in_data_6,
  input  [7:0]   io_pipe_phv_in_data_7,
  input  [7:0]   io_pipe_phv_in_data_8,
  input  [7:0]   io_pipe_phv_in_data_9,
  input  [7:0]   io_pipe_phv_in_data_10,
  input  [7:0]   io_pipe_phv_in_data_11,
  input  [7:0]   io_pipe_phv_in_data_12,
  input  [7:0]   io_pipe_phv_in_data_13,
  input  [7:0]   io_pipe_phv_in_data_14,
  input  [7:0]   io_pipe_phv_in_data_15,
  input  [7:0]   io_pipe_phv_in_data_16,
  input  [7:0]   io_pipe_phv_in_data_17,
  input  [7:0]   io_pipe_phv_in_data_18,
  input  [7:0]   io_pipe_phv_in_data_19,
  input  [7:0]   io_pipe_phv_in_data_20,
  input  [7:0]   io_pipe_phv_in_data_21,
  input  [7:0]   io_pipe_phv_in_data_22,
  input  [7:0]   io_pipe_phv_in_data_23,
  input  [7:0]   io_pipe_phv_in_data_24,
  input  [7:0]   io_pipe_phv_in_data_25,
  input  [7:0]   io_pipe_phv_in_data_26,
  input  [7:0]   io_pipe_phv_in_data_27,
  input  [7:0]   io_pipe_phv_in_data_28,
  input  [7:0]   io_pipe_phv_in_data_29,
  input  [7:0]   io_pipe_phv_in_data_30,
  input  [7:0]   io_pipe_phv_in_data_31,
  input  [7:0]   io_pipe_phv_in_data_32,
  input  [7:0]   io_pipe_phv_in_data_33,
  input  [7:0]   io_pipe_phv_in_data_34,
  input  [7:0]   io_pipe_phv_in_data_35,
  input  [7:0]   io_pipe_phv_in_data_36,
  input  [7:0]   io_pipe_phv_in_data_37,
  input  [7:0]   io_pipe_phv_in_data_38,
  input  [7:0]   io_pipe_phv_in_data_39,
  input  [7:0]   io_pipe_phv_in_data_40,
  input  [7:0]   io_pipe_phv_in_data_41,
  input  [7:0]   io_pipe_phv_in_data_42,
  input  [7:0]   io_pipe_phv_in_data_43,
  input  [7:0]   io_pipe_phv_in_data_44,
  input  [7:0]   io_pipe_phv_in_data_45,
  input  [7:0]   io_pipe_phv_in_data_46,
  input  [7:0]   io_pipe_phv_in_data_47,
  input  [7:0]   io_pipe_phv_in_data_48,
  input  [7:0]   io_pipe_phv_in_data_49,
  input  [7:0]   io_pipe_phv_in_data_50,
  input  [7:0]   io_pipe_phv_in_data_51,
  input  [7:0]   io_pipe_phv_in_data_52,
  input  [7:0]   io_pipe_phv_in_data_53,
  input  [7:0]   io_pipe_phv_in_data_54,
  input  [7:0]   io_pipe_phv_in_data_55,
  input  [7:0]   io_pipe_phv_in_data_56,
  input  [7:0]   io_pipe_phv_in_data_57,
  input  [7:0]   io_pipe_phv_in_data_58,
  input  [7:0]   io_pipe_phv_in_data_59,
  input  [7:0]   io_pipe_phv_in_data_60,
  input  [7:0]   io_pipe_phv_in_data_61,
  input  [7:0]   io_pipe_phv_in_data_62,
  input  [7:0]   io_pipe_phv_in_data_63,
  input  [7:0]   io_pipe_phv_in_data_64,
  input  [7:0]   io_pipe_phv_in_data_65,
  input  [7:0]   io_pipe_phv_in_data_66,
  input  [7:0]   io_pipe_phv_in_data_67,
  input  [7:0]   io_pipe_phv_in_data_68,
  input  [7:0]   io_pipe_phv_in_data_69,
  input  [7:0]   io_pipe_phv_in_data_70,
  input  [7:0]   io_pipe_phv_in_data_71,
  input  [7:0]   io_pipe_phv_in_data_72,
  input  [7:0]   io_pipe_phv_in_data_73,
  input  [7:0]   io_pipe_phv_in_data_74,
  input  [7:0]   io_pipe_phv_in_data_75,
  input  [7:0]   io_pipe_phv_in_data_76,
  input  [7:0]   io_pipe_phv_in_data_77,
  input  [7:0]   io_pipe_phv_in_data_78,
  input  [7:0]   io_pipe_phv_in_data_79,
  input  [7:0]   io_pipe_phv_in_data_80,
  input  [7:0]   io_pipe_phv_in_data_81,
  input  [7:0]   io_pipe_phv_in_data_82,
  input  [7:0]   io_pipe_phv_in_data_83,
  input  [7:0]   io_pipe_phv_in_data_84,
  input  [7:0]   io_pipe_phv_in_data_85,
  input  [7:0]   io_pipe_phv_in_data_86,
  input  [7:0]   io_pipe_phv_in_data_87,
  input  [7:0]   io_pipe_phv_in_data_88,
  input  [7:0]   io_pipe_phv_in_data_89,
  input  [7:0]   io_pipe_phv_in_data_90,
  input  [7:0]   io_pipe_phv_in_data_91,
  input  [7:0]   io_pipe_phv_in_data_92,
  input  [7:0]   io_pipe_phv_in_data_93,
  input  [7:0]   io_pipe_phv_in_data_94,
  input  [7:0]   io_pipe_phv_in_data_95,
  input  [15:0]  io_pipe_phv_in_header_0,
  input  [15:0]  io_pipe_phv_in_header_1,
  input  [15:0]  io_pipe_phv_in_header_2,
  input  [15:0]  io_pipe_phv_in_header_3,
  input  [15:0]  io_pipe_phv_in_header_4,
  input  [15:0]  io_pipe_phv_in_header_5,
  input  [15:0]  io_pipe_phv_in_header_6,
  input  [15:0]  io_pipe_phv_in_header_7,
  input  [15:0]  io_pipe_phv_in_header_8,
  input  [15:0]  io_pipe_phv_in_header_9,
  input  [15:0]  io_pipe_phv_in_header_10,
  input  [15:0]  io_pipe_phv_in_header_11,
  input  [15:0]  io_pipe_phv_in_header_12,
  input  [15:0]  io_pipe_phv_in_header_13,
  input  [15:0]  io_pipe_phv_in_header_14,
  input  [15:0]  io_pipe_phv_in_header_15,
  input  [7:0]   io_pipe_phv_in_parse_current_state,
  input  [7:0]   io_pipe_phv_in_parse_current_offset,
  input  [15:0]  io_pipe_phv_in_parse_transition_field,
  input  [1:0]   io_pipe_phv_in_next_processor_id,
  input          io_pipe_phv_in_next_config_id,
  input          io_pipe_phv_in_is_valid_processor,
  output [7:0]   io_pipe_phv_out_data_0,
  output [7:0]   io_pipe_phv_out_data_1,
  output [7:0]   io_pipe_phv_out_data_2,
  output [7:0]   io_pipe_phv_out_data_3,
  output [7:0]   io_pipe_phv_out_data_4,
  output [7:0]   io_pipe_phv_out_data_5,
  output [7:0]   io_pipe_phv_out_data_6,
  output [7:0]   io_pipe_phv_out_data_7,
  output [7:0]   io_pipe_phv_out_data_8,
  output [7:0]   io_pipe_phv_out_data_9,
  output [7:0]   io_pipe_phv_out_data_10,
  output [7:0]   io_pipe_phv_out_data_11,
  output [7:0]   io_pipe_phv_out_data_12,
  output [7:0]   io_pipe_phv_out_data_13,
  output [7:0]   io_pipe_phv_out_data_14,
  output [7:0]   io_pipe_phv_out_data_15,
  output [7:0]   io_pipe_phv_out_data_16,
  output [7:0]   io_pipe_phv_out_data_17,
  output [7:0]   io_pipe_phv_out_data_18,
  output [7:0]   io_pipe_phv_out_data_19,
  output [7:0]   io_pipe_phv_out_data_20,
  output [7:0]   io_pipe_phv_out_data_21,
  output [7:0]   io_pipe_phv_out_data_22,
  output [7:0]   io_pipe_phv_out_data_23,
  output [7:0]   io_pipe_phv_out_data_24,
  output [7:0]   io_pipe_phv_out_data_25,
  output [7:0]   io_pipe_phv_out_data_26,
  output [7:0]   io_pipe_phv_out_data_27,
  output [7:0]   io_pipe_phv_out_data_28,
  output [7:0]   io_pipe_phv_out_data_29,
  output [7:0]   io_pipe_phv_out_data_30,
  output [7:0]   io_pipe_phv_out_data_31,
  output [7:0]   io_pipe_phv_out_data_32,
  output [7:0]   io_pipe_phv_out_data_33,
  output [7:0]   io_pipe_phv_out_data_34,
  output [7:0]   io_pipe_phv_out_data_35,
  output [7:0]   io_pipe_phv_out_data_36,
  output [7:0]   io_pipe_phv_out_data_37,
  output [7:0]   io_pipe_phv_out_data_38,
  output [7:0]   io_pipe_phv_out_data_39,
  output [7:0]   io_pipe_phv_out_data_40,
  output [7:0]   io_pipe_phv_out_data_41,
  output [7:0]   io_pipe_phv_out_data_42,
  output [7:0]   io_pipe_phv_out_data_43,
  output [7:0]   io_pipe_phv_out_data_44,
  output [7:0]   io_pipe_phv_out_data_45,
  output [7:0]   io_pipe_phv_out_data_46,
  output [7:0]   io_pipe_phv_out_data_47,
  output [7:0]   io_pipe_phv_out_data_48,
  output [7:0]   io_pipe_phv_out_data_49,
  output [7:0]   io_pipe_phv_out_data_50,
  output [7:0]   io_pipe_phv_out_data_51,
  output [7:0]   io_pipe_phv_out_data_52,
  output [7:0]   io_pipe_phv_out_data_53,
  output [7:0]   io_pipe_phv_out_data_54,
  output [7:0]   io_pipe_phv_out_data_55,
  output [7:0]   io_pipe_phv_out_data_56,
  output [7:0]   io_pipe_phv_out_data_57,
  output [7:0]   io_pipe_phv_out_data_58,
  output [7:0]   io_pipe_phv_out_data_59,
  output [7:0]   io_pipe_phv_out_data_60,
  output [7:0]   io_pipe_phv_out_data_61,
  output [7:0]   io_pipe_phv_out_data_62,
  output [7:0]   io_pipe_phv_out_data_63,
  output [7:0]   io_pipe_phv_out_data_64,
  output [7:0]   io_pipe_phv_out_data_65,
  output [7:0]   io_pipe_phv_out_data_66,
  output [7:0]   io_pipe_phv_out_data_67,
  output [7:0]   io_pipe_phv_out_data_68,
  output [7:0]   io_pipe_phv_out_data_69,
  output [7:0]   io_pipe_phv_out_data_70,
  output [7:0]   io_pipe_phv_out_data_71,
  output [7:0]   io_pipe_phv_out_data_72,
  output [7:0]   io_pipe_phv_out_data_73,
  output [7:0]   io_pipe_phv_out_data_74,
  output [7:0]   io_pipe_phv_out_data_75,
  output [7:0]   io_pipe_phv_out_data_76,
  output [7:0]   io_pipe_phv_out_data_77,
  output [7:0]   io_pipe_phv_out_data_78,
  output [7:0]   io_pipe_phv_out_data_79,
  output [7:0]   io_pipe_phv_out_data_80,
  output [7:0]   io_pipe_phv_out_data_81,
  output [7:0]   io_pipe_phv_out_data_82,
  output [7:0]   io_pipe_phv_out_data_83,
  output [7:0]   io_pipe_phv_out_data_84,
  output [7:0]   io_pipe_phv_out_data_85,
  output [7:0]   io_pipe_phv_out_data_86,
  output [7:0]   io_pipe_phv_out_data_87,
  output [7:0]   io_pipe_phv_out_data_88,
  output [7:0]   io_pipe_phv_out_data_89,
  output [7:0]   io_pipe_phv_out_data_90,
  output [7:0]   io_pipe_phv_out_data_91,
  output [7:0]   io_pipe_phv_out_data_92,
  output [7:0]   io_pipe_phv_out_data_93,
  output [7:0]   io_pipe_phv_out_data_94,
  output [7:0]   io_pipe_phv_out_data_95,
  output [15:0]  io_pipe_phv_out_header_0,
  output [15:0]  io_pipe_phv_out_header_1,
  output [15:0]  io_pipe_phv_out_header_2,
  output [15:0]  io_pipe_phv_out_header_3,
  output [15:0]  io_pipe_phv_out_header_4,
  output [15:0]  io_pipe_phv_out_header_5,
  output [15:0]  io_pipe_phv_out_header_6,
  output [15:0]  io_pipe_phv_out_header_7,
  output [15:0]  io_pipe_phv_out_header_8,
  output [15:0]  io_pipe_phv_out_header_9,
  output [15:0]  io_pipe_phv_out_header_10,
  output [15:0]  io_pipe_phv_out_header_11,
  output [15:0]  io_pipe_phv_out_header_12,
  output [15:0]  io_pipe_phv_out_header_13,
  output [15:0]  io_pipe_phv_out_header_14,
  output [15:0]  io_pipe_phv_out_header_15,
  output [7:0]   io_pipe_phv_out_parse_current_state,
  output [7:0]   io_pipe_phv_out_parse_current_offset,
  output [15:0]  io_pipe_phv_out_parse_transition_field,
  output [1:0]   io_pipe_phv_out_next_processor_id,
  output         io_pipe_phv_out_next_config_id,
  output         io_pipe_phv_out_is_valid_processor,
  input  [3:0]   io_key_config_0_key_length,
  input  [3:0]   io_key_config_1_key_length,
  input  [63:0]  io_key_in,
  input  [127:0] io_data_in,
  output         io_hit,
  output [63:0]  io_match_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [127:0] _RAND_119;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[matcher.scala 226:22]
  reg [7:0] phv_data_1; // @[matcher.scala 226:22]
  reg [7:0] phv_data_2; // @[matcher.scala 226:22]
  reg [7:0] phv_data_3; // @[matcher.scala 226:22]
  reg [7:0] phv_data_4; // @[matcher.scala 226:22]
  reg [7:0] phv_data_5; // @[matcher.scala 226:22]
  reg [7:0] phv_data_6; // @[matcher.scala 226:22]
  reg [7:0] phv_data_7; // @[matcher.scala 226:22]
  reg [7:0] phv_data_8; // @[matcher.scala 226:22]
  reg [7:0] phv_data_9; // @[matcher.scala 226:22]
  reg [7:0] phv_data_10; // @[matcher.scala 226:22]
  reg [7:0] phv_data_11; // @[matcher.scala 226:22]
  reg [7:0] phv_data_12; // @[matcher.scala 226:22]
  reg [7:0] phv_data_13; // @[matcher.scala 226:22]
  reg [7:0] phv_data_14; // @[matcher.scala 226:22]
  reg [7:0] phv_data_15; // @[matcher.scala 226:22]
  reg [7:0] phv_data_16; // @[matcher.scala 226:22]
  reg [7:0] phv_data_17; // @[matcher.scala 226:22]
  reg [7:0] phv_data_18; // @[matcher.scala 226:22]
  reg [7:0] phv_data_19; // @[matcher.scala 226:22]
  reg [7:0] phv_data_20; // @[matcher.scala 226:22]
  reg [7:0] phv_data_21; // @[matcher.scala 226:22]
  reg [7:0] phv_data_22; // @[matcher.scala 226:22]
  reg [7:0] phv_data_23; // @[matcher.scala 226:22]
  reg [7:0] phv_data_24; // @[matcher.scala 226:22]
  reg [7:0] phv_data_25; // @[matcher.scala 226:22]
  reg [7:0] phv_data_26; // @[matcher.scala 226:22]
  reg [7:0] phv_data_27; // @[matcher.scala 226:22]
  reg [7:0] phv_data_28; // @[matcher.scala 226:22]
  reg [7:0] phv_data_29; // @[matcher.scala 226:22]
  reg [7:0] phv_data_30; // @[matcher.scala 226:22]
  reg [7:0] phv_data_31; // @[matcher.scala 226:22]
  reg [7:0] phv_data_32; // @[matcher.scala 226:22]
  reg [7:0] phv_data_33; // @[matcher.scala 226:22]
  reg [7:0] phv_data_34; // @[matcher.scala 226:22]
  reg [7:0] phv_data_35; // @[matcher.scala 226:22]
  reg [7:0] phv_data_36; // @[matcher.scala 226:22]
  reg [7:0] phv_data_37; // @[matcher.scala 226:22]
  reg [7:0] phv_data_38; // @[matcher.scala 226:22]
  reg [7:0] phv_data_39; // @[matcher.scala 226:22]
  reg [7:0] phv_data_40; // @[matcher.scala 226:22]
  reg [7:0] phv_data_41; // @[matcher.scala 226:22]
  reg [7:0] phv_data_42; // @[matcher.scala 226:22]
  reg [7:0] phv_data_43; // @[matcher.scala 226:22]
  reg [7:0] phv_data_44; // @[matcher.scala 226:22]
  reg [7:0] phv_data_45; // @[matcher.scala 226:22]
  reg [7:0] phv_data_46; // @[matcher.scala 226:22]
  reg [7:0] phv_data_47; // @[matcher.scala 226:22]
  reg [7:0] phv_data_48; // @[matcher.scala 226:22]
  reg [7:0] phv_data_49; // @[matcher.scala 226:22]
  reg [7:0] phv_data_50; // @[matcher.scala 226:22]
  reg [7:0] phv_data_51; // @[matcher.scala 226:22]
  reg [7:0] phv_data_52; // @[matcher.scala 226:22]
  reg [7:0] phv_data_53; // @[matcher.scala 226:22]
  reg [7:0] phv_data_54; // @[matcher.scala 226:22]
  reg [7:0] phv_data_55; // @[matcher.scala 226:22]
  reg [7:0] phv_data_56; // @[matcher.scala 226:22]
  reg [7:0] phv_data_57; // @[matcher.scala 226:22]
  reg [7:0] phv_data_58; // @[matcher.scala 226:22]
  reg [7:0] phv_data_59; // @[matcher.scala 226:22]
  reg [7:0] phv_data_60; // @[matcher.scala 226:22]
  reg [7:0] phv_data_61; // @[matcher.scala 226:22]
  reg [7:0] phv_data_62; // @[matcher.scala 226:22]
  reg [7:0] phv_data_63; // @[matcher.scala 226:22]
  reg [7:0] phv_data_64; // @[matcher.scala 226:22]
  reg [7:0] phv_data_65; // @[matcher.scala 226:22]
  reg [7:0] phv_data_66; // @[matcher.scala 226:22]
  reg [7:0] phv_data_67; // @[matcher.scala 226:22]
  reg [7:0] phv_data_68; // @[matcher.scala 226:22]
  reg [7:0] phv_data_69; // @[matcher.scala 226:22]
  reg [7:0] phv_data_70; // @[matcher.scala 226:22]
  reg [7:0] phv_data_71; // @[matcher.scala 226:22]
  reg [7:0] phv_data_72; // @[matcher.scala 226:22]
  reg [7:0] phv_data_73; // @[matcher.scala 226:22]
  reg [7:0] phv_data_74; // @[matcher.scala 226:22]
  reg [7:0] phv_data_75; // @[matcher.scala 226:22]
  reg [7:0] phv_data_76; // @[matcher.scala 226:22]
  reg [7:0] phv_data_77; // @[matcher.scala 226:22]
  reg [7:0] phv_data_78; // @[matcher.scala 226:22]
  reg [7:0] phv_data_79; // @[matcher.scala 226:22]
  reg [7:0] phv_data_80; // @[matcher.scala 226:22]
  reg [7:0] phv_data_81; // @[matcher.scala 226:22]
  reg [7:0] phv_data_82; // @[matcher.scala 226:22]
  reg [7:0] phv_data_83; // @[matcher.scala 226:22]
  reg [7:0] phv_data_84; // @[matcher.scala 226:22]
  reg [7:0] phv_data_85; // @[matcher.scala 226:22]
  reg [7:0] phv_data_86; // @[matcher.scala 226:22]
  reg [7:0] phv_data_87; // @[matcher.scala 226:22]
  reg [7:0] phv_data_88; // @[matcher.scala 226:22]
  reg [7:0] phv_data_89; // @[matcher.scala 226:22]
  reg [7:0] phv_data_90; // @[matcher.scala 226:22]
  reg [7:0] phv_data_91; // @[matcher.scala 226:22]
  reg [7:0] phv_data_92; // @[matcher.scala 226:22]
  reg [7:0] phv_data_93; // @[matcher.scala 226:22]
  reg [7:0] phv_data_94; // @[matcher.scala 226:22]
  reg [7:0] phv_data_95; // @[matcher.scala 226:22]
  reg [15:0] phv_header_0; // @[matcher.scala 226:22]
  reg [15:0] phv_header_1; // @[matcher.scala 226:22]
  reg [15:0] phv_header_2; // @[matcher.scala 226:22]
  reg [15:0] phv_header_3; // @[matcher.scala 226:22]
  reg [15:0] phv_header_4; // @[matcher.scala 226:22]
  reg [15:0] phv_header_5; // @[matcher.scala 226:22]
  reg [15:0] phv_header_6; // @[matcher.scala 226:22]
  reg [15:0] phv_header_7; // @[matcher.scala 226:22]
  reg [15:0] phv_header_8; // @[matcher.scala 226:22]
  reg [15:0] phv_header_9; // @[matcher.scala 226:22]
  reg [15:0] phv_header_10; // @[matcher.scala 226:22]
  reg [15:0] phv_header_11; // @[matcher.scala 226:22]
  reg [15:0] phv_header_12; // @[matcher.scala 226:22]
  reg [15:0] phv_header_13; // @[matcher.scala 226:22]
  reg [15:0] phv_header_14; // @[matcher.scala 226:22]
  reg [15:0] phv_header_15; // @[matcher.scala 226:22]
  reg [7:0] phv_parse_current_state; // @[matcher.scala 226:22]
  reg [7:0] phv_parse_current_offset; // @[matcher.scala 226:22]
  reg [15:0] phv_parse_transition_field; // @[matcher.scala 226:22]
  reg [1:0] phv_next_processor_id; // @[matcher.scala 226:22]
  reg  phv_next_config_id; // @[matcher.scala 226:22]
  reg  phv_is_valid_processor; // @[matcher.scala 226:22]
  reg [63:0] key; // @[matcher.scala 230:22]
  reg [127:0] data; // @[matcher.scala 232:23]
  wire [7:0] key_byte = key[63:56]; // @[matcher.scala 240:35]
  wire [7:0] data_byte = data[127:120]; // @[matcher.scala 241:37]
  wire [3:0] _GEN_6 = phv_next_config_id ? io_key_config_1_key_length : io_key_config_0_key_length; // @[matcher.scala 242:65 matcher.scala 242:65]
  wire  key_equal_0 = 4'h0 < _GEN_6 ? key_byte == data_byte : 1'h1; // @[matcher.scala 242:90 matcher.scala 243:34 matcher.scala 245:34]
  wire [7:0] key_byte_1 = key[55:48]; // @[matcher.scala 240:35]
  wire [7:0] data_byte_1 = data[119:112]; // @[matcher.scala 241:37]
  wire  key_equal_1 = 4'h1 < _GEN_6 ? key_byte_1 == data_byte_1 : 1'h1; // @[matcher.scala 242:90 matcher.scala 243:34 matcher.scala 245:34]
  wire [7:0] key_byte_2 = key[47:40]; // @[matcher.scala 240:35]
  wire [7:0] data_byte_2 = data[111:104]; // @[matcher.scala 241:37]
  wire  key_equal_2 = 4'h2 < _GEN_6 ? key_byte_2 == data_byte_2 : 1'h1; // @[matcher.scala 242:90 matcher.scala 243:34 matcher.scala 245:34]
  wire [7:0] key_byte_3 = key[39:32]; // @[matcher.scala 240:35]
  wire [7:0] data_byte_3 = data[103:96]; // @[matcher.scala 241:37]
  wire  key_equal_3 = 4'h3 < _GEN_6 ? key_byte_3 == data_byte_3 : 1'h1; // @[matcher.scala 242:90 matcher.scala 243:34 matcher.scala 245:34]
  wire [7:0] key_byte_4 = key[31:24]; // @[matcher.scala 240:35]
  wire [7:0] data_byte_4 = data[95:88]; // @[matcher.scala 241:37]
  wire  key_equal_4 = 4'h4 < _GEN_6 ? key_byte_4 == data_byte_4 : 1'h1; // @[matcher.scala 242:90 matcher.scala 243:34 matcher.scala 245:34]
  wire [7:0] key_byte_5 = key[23:16]; // @[matcher.scala 240:35]
  wire [7:0] data_byte_5 = data[87:80]; // @[matcher.scala 241:37]
  wire  key_equal_5 = 4'h5 < _GEN_6 ? key_byte_5 == data_byte_5 : 1'h1; // @[matcher.scala 242:90 matcher.scala 243:34 matcher.scala 245:34]
  wire [7:0] key_byte_6 = key[15:8]; // @[matcher.scala 240:35]
  wire [7:0] data_byte_6 = data[79:72]; // @[matcher.scala 241:37]
  wire  key_equal_6 = 4'h6 < _GEN_6 ? key_byte_6 == data_byte_6 : 1'h1; // @[matcher.scala 242:90 matcher.scala 243:34 matcher.scala 245:34]
  wire [7:0] key_byte_7 = key[7:0]; // @[matcher.scala 240:35]
  wire [7:0] data_byte_7 = data[71:64]; // @[matcher.scala 241:37]
  wire  key_equal_7 = 4'h7 < _GEN_6 ? key_byte_7 == data_byte_7 : 1'h1; // @[matcher.scala 242:90 matcher.scala 243:34 matcher.scala 245:34]
  wire [63:0] _GEN_16 = 4'h1 == _GEN_6 ? data[119:56] : 64'h0; // @[matcher.scala 252:92 matcher.scala 253:36 matcher.scala 250:28]
  wire [63:0] _GEN_17 = 4'h2 == _GEN_6 ? data[111:48] : _GEN_16; // @[matcher.scala 252:92 matcher.scala 253:36]
  wire [63:0] _GEN_18 = 4'h3 == _GEN_6 ? data[103:40] : _GEN_17; // @[matcher.scala 252:92 matcher.scala 253:36]
  wire [63:0] _GEN_19 = 4'h4 == _GEN_6 ? data[95:32] : _GEN_18; // @[matcher.scala 252:92 matcher.scala 253:36]
  wire [63:0] _GEN_20 = 4'h5 == _GEN_6 ? data[87:24] : _GEN_19; // @[matcher.scala 252:92 matcher.scala 253:36]
  wire [63:0] _GEN_21 = 4'h6 == _GEN_6 ? data[79:16] : _GEN_20; // @[matcher.scala 252:92 matcher.scala 253:36]
  wire [63:0] _GEN_22 = 4'h7 == _GEN_6 ? data[71:8] : _GEN_21; // @[matcher.scala 252:92 matcher.scala 253:36]
  wire [63:0] _GEN_23 = 4'h8 == _GEN_6 ? data[63:0] : _GEN_22; // @[matcher.scala 252:92 matcher.scala 253:36]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[matcher.scala 228:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[matcher.scala 228:25]
  assign io_hit = phv_is_valid_processor & (key_equal_0 & key_equal_1 & key_equal_2 & key_equal_3 & key_equal_4 &
    key_equal_5 & key_equal_6 & key_equal_7); // @[matcher.scala 235:39 matcher.scala 249:20 matcher.scala 257:20]
  assign io_match_value = phv_is_valid_processor ? _GEN_23 : 64'h0; // @[matcher.scala 235:39 matcher.scala 258:28]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[matcher.scala 227:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[matcher.scala 227:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[matcher.scala 227:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[matcher.scala 227:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[matcher.scala 227:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[matcher.scala 227:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[matcher.scala 227:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[matcher.scala 227:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[matcher.scala 227:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[matcher.scala 227:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[matcher.scala 227:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[matcher.scala 227:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[matcher.scala 227:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[matcher.scala 227:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[matcher.scala 227:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[matcher.scala 227:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[matcher.scala 227:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[matcher.scala 227:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[matcher.scala 227:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[matcher.scala 227:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[matcher.scala 227:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[matcher.scala 227:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[matcher.scala 227:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[matcher.scala 227:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[matcher.scala 227:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[matcher.scala 227:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[matcher.scala 227:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[matcher.scala 227:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[matcher.scala 227:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[matcher.scala 227:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[matcher.scala 227:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[matcher.scala 227:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[matcher.scala 227:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[matcher.scala 227:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[matcher.scala 227:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[matcher.scala 227:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[matcher.scala 227:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[matcher.scala 227:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[matcher.scala 227:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[matcher.scala 227:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[matcher.scala 227:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[matcher.scala 227:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[matcher.scala 227:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[matcher.scala 227:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[matcher.scala 227:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[matcher.scala 227:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[matcher.scala 227:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[matcher.scala 227:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[matcher.scala 227:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[matcher.scala 227:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[matcher.scala 227:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[matcher.scala 227:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[matcher.scala 227:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[matcher.scala 227:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[matcher.scala 227:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[matcher.scala 227:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[matcher.scala 227:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[matcher.scala 227:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[matcher.scala 227:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[matcher.scala 227:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[matcher.scala 227:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[matcher.scala 227:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[matcher.scala 227:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[matcher.scala 227:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[matcher.scala 227:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[matcher.scala 227:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[matcher.scala 227:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[matcher.scala 227:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[matcher.scala 227:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[matcher.scala 227:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[matcher.scala 227:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[matcher.scala 227:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[matcher.scala 227:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[matcher.scala 227:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[matcher.scala 227:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[matcher.scala 227:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[matcher.scala 227:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[matcher.scala 227:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[matcher.scala 227:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[matcher.scala 227:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[matcher.scala 227:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[matcher.scala 227:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[matcher.scala 227:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[matcher.scala 227:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[matcher.scala 227:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[matcher.scala 227:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[matcher.scala 227:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[matcher.scala 227:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[matcher.scala 227:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[matcher.scala 227:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[matcher.scala 227:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[matcher.scala 227:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[matcher.scala 227:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[matcher.scala 227:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[matcher.scala 227:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[matcher.scala 227:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[matcher.scala 227:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[matcher.scala 227:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[matcher.scala 227:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[matcher.scala 227:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[matcher.scala 227:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[matcher.scala 227:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[matcher.scala 227:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[matcher.scala 227:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[matcher.scala 227:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[matcher.scala 227:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[matcher.scala 227:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[matcher.scala 227:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[matcher.scala 227:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[matcher.scala 227:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[matcher.scala 227:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[matcher.scala 227:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[matcher.scala 227:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[matcher.scala 227:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[matcher.scala 227:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[matcher.scala 227:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[matcher.scala 227:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[matcher.scala 227:13]
    key <= io_key_in; // @[matcher.scala 231:13]
    data <= io_data_in; // @[matcher.scala 233:14]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  phv_next_config_id = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_117[0:0];
  _RAND_118 = {2{`RANDOM}};
  key = _RAND_118[63:0];
  _RAND_119 = {4{`RANDOM}};
  data = _RAND_119[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Matcher(
  input         clock,
  input         reset,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input         io_mod_en,
  input         io_mod_config_id,
  input  [7:0]  io_mod_key_mod_header_id,
  input  [7:0]  io_mod_key_mod_internal_offset,
  input  [3:0]  io_mod_key_mod_key_length,
  input  [3:0]  io_mod_key_mod_val_length,
  input  [2:0]  io_mod_table_mod_sram_id_table_0,
  input  [2:0]  io_mod_table_mod_sram_id_table_1,
  input  [2:0]  io_mod_table_mod_sram_id_table_2,
  input  [2:0]  io_mod_table_mod_sram_id_table_3,
  input  [2:0]  io_mod_table_mod_sram_id_table_4,
  input  [2:0]  io_mod_table_mod_sram_id_table_5,
  input  [2:0]  io_mod_table_mod_sram_id_table_6,
  input  [2:0]  io_mod_table_mod_sram_id_table_7,
  input  [3:0]  io_mod_table_mod_table_width,
  input  [3:0]  io_mod_table_mod_table_depth,
  output        io_hit,
  output [63:0] io_match_value,
  output        io_mem_cluster_0_en,
  output [7:0]  io_mem_cluster_0_addr,
  input  [63:0] io_mem_cluster_0_data,
  output        io_mem_cluster_1_en,
  output [7:0]  io_mem_cluster_1_addr,
  input  [63:0] io_mem_cluster_1_data,
  output        io_mem_cluster_2_en,
  output [7:0]  io_mem_cluster_2_addr,
  input  [63:0] io_mem_cluster_2_data,
  output        io_mem_cluster_3_en,
  output [7:0]  io_mem_cluster_3_addr,
  input  [63:0] io_mem_cluster_3_data,
  output        io_mem_cluster_4_en,
  output [7:0]  io_mem_cluster_4_addr,
  input  [63:0] io_mem_cluster_4_data,
  output        io_mem_cluster_5_en,
  output [7:0]  io_mem_cluster_5_addr,
  input  [63:0] io_mem_cluster_5_data,
  output        io_mem_cluster_6_en,
  output [7:0]  io_mem_cluster_6_addr,
  input  [63:0] io_mem_cluster_6_data,
  output        io_mem_cluster_7_en,
  output [7:0]  io_mem_cluster_7_addr,
  input  [63:0] io_mem_cluster_7_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  pipe1_clock; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_0; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_1; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_2; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_3; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_4; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_5; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_6; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_7; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_8; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_9; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_10; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_11; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_12; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_13; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_14; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_15; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_16; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_17; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_18; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_19; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_20; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_21; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_22; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_23; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_24; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_25; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_26; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_27; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_28; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_29; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_30; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_31; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_32; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_33; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_34; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_35; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_36; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_37; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_38; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_39; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_40; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_41; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_42; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_43; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_44; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_45; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_46; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_47; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_48; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_49; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_50; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_51; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_52; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_53; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_54; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_55; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_56; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_57; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_58; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_59; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_60; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_61; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_62; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_63; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_64; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_65; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_66; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_67; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_68; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_69; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_70; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_71; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_72; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_73; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_74; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_75; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_76; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_77; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_78; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_79; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_80; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_81; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_82; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_83; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_84; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_85; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_86; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_87; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_88; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_89; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_90; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_91; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_92; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_93; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_94; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_95; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_0; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_1; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_2; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_3; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_4; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_5; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_6; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_7; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_8; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_9; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_10; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_11; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_12; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_13; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_14; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_15; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_state; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 263:23]
  wire [1:0] pipe1_io_pipe_phv_in_next_processor_id; // @[matcher.scala 263:23]
  wire  pipe1_io_pipe_phv_in_next_config_id; // @[matcher.scala 263:23]
  wire  pipe1_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_0; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_1; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_2; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_3; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_4; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_5; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_6; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_7; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_8; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_9; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_10; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_11; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_12; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_13; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_14; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_15; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_16; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_17; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_18; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_19; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_20; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_21; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_22; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_23; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_24; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_25; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_26; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_27; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_28; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_29; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_30; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_31; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_32; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_33; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_34; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_35; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_36; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_37; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_38; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_39; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_40; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_41; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_42; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_43; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_44; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_45; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_46; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_47; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_48; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_49; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_50; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_51; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_52; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_53; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_54; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_55; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_56; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_57; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_58; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_59; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_60; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_61; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_62; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_63; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_64; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_65; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_66; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_67; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_68; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_69; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_70; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_71; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_72; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_73; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_74; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_75; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_76; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_77; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_78; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_79; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_80; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_81; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_82; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_83; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_84; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_85; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_86; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_87; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_88; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_89; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_90; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_91; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_92; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_93; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_94; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_95; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_0; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_1; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_2; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_3; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_4; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_5; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_6; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_7; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_8; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_9; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_10; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_11; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_12; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_13; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_14; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_15; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_state; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 263:23]
  wire [15:0] pipe1_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 263:23]
  wire [1:0] pipe1_io_pipe_phv_out_next_processor_id; // @[matcher.scala 263:23]
  wire  pipe1_io_pipe_phv_out_next_config_id; // @[matcher.scala 263:23]
  wire  pipe1_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_key_config_0_header_id; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_key_config_0_internal_offset; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_key_config_1_header_id; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_key_config_1_internal_offset; // @[matcher.scala 263:23]
  wire [7:0] pipe1_io_key_offset; // @[matcher.scala 263:23]
  wire  pipe2_clock; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_0; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_1; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_2; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_3; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_4; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_5; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_6; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_7; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_8; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_9; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_10; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_11; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_12; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_13; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_14; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_15; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_16; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_17; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_18; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_19; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_20; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_21; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_22; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_23; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_24; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_25; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_26; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_27; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_28; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_29; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_30; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_31; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_32; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_33; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_34; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_35; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_36; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_37; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_38; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_39; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_40; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_41; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_42; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_43; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_44; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_45; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_46; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_47; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_48; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_49; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_50; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_51; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_52; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_53; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_54; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_55; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_56; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_57; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_58; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_59; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_60; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_61; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_62; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_63; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_64; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_65; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_66; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_67; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_68; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_69; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_70; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_71; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_72; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_73; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_74; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_75; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_76; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_77; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_78; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_79; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_80; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_81; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_82; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_83; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_84; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_85; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_86; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_87; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_88; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_89; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_90; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_91; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_92; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_93; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_94; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_95; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_0; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_1; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_2; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_3; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_4; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_5; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_6; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_7; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_8; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_9; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_10; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_11; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_12; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_13; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_14; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_15; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_state; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 264:23]
  wire [1:0] pipe2_io_pipe_phv_in_next_processor_id; // @[matcher.scala 264:23]
  wire  pipe2_io_pipe_phv_in_next_config_id; // @[matcher.scala 264:23]
  wire  pipe2_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_0; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_1; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_2; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_3; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_4; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_5; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_6; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_7; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_8; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_9; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_10; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_11; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_12; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_13; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_14; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_15; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_16; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_17; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_18; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_19; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_20; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_21; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_22; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_23; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_24; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_25; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_26; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_27; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_28; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_29; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_30; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_31; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_32; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_33; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_34; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_35; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_36; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_37; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_38; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_39; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_40; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_41; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_42; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_43; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_44; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_45; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_46; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_47; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_48; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_49; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_50; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_51; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_52; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_53; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_54; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_55; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_56; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_57; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_58; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_59; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_60; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_61; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_62; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_63; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_64; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_65; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_66; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_67; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_68; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_69; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_70; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_71; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_72; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_73; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_74; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_75; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_76; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_77; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_78; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_79; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_80; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_81; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_82; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_83; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_84; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_85; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_86; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_87; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_88; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_89; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_90; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_91; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_92; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_93; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_94; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_95; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_0; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_1; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_2; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_3; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_4; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_5; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_6; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_7; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_8; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_9; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_10; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_11; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_12; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_13; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_14; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_15; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_state; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 264:23]
  wire [15:0] pipe2_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 264:23]
  wire [1:0] pipe2_io_pipe_phv_out_next_processor_id; // @[matcher.scala 264:23]
  wire  pipe2_io_pipe_phv_out_next_config_id; // @[matcher.scala 264:23]
  wire  pipe2_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 264:23]
  wire [3:0] pipe2_io_key_config_0_key_length; // @[matcher.scala 264:23]
  wire [3:0] pipe2_io_key_config_1_key_length; // @[matcher.scala 264:23]
  wire [7:0] pipe2_io_key_offset; // @[matcher.scala 264:23]
  wire [63:0] pipe2_io_match_key; // @[matcher.scala 264:23]
  wire  pipe3to8_clock; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_0; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_1; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_2; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_3; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_4; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_5; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_6; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_7; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_8; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_9; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_10; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_11; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_12; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_13; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_14; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_15; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_16; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_17; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_18; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_19; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_20; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_21; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_22; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_23; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_24; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_25; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_26; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_27; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_28; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_29; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_30; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_31; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_32; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_33; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_34; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_35; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_36; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_37; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_38; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_39; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_40; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_41; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_42; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_43; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_44; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_45; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_46; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_47; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_48; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_49; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_50; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_51; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_52; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_53; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_54; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_55; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_56; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_57; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_58; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_59; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_60; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_61; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_62; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_63; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_64; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_65; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_66; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_67; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_68; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_69; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_70; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_71; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_72; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_73; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_74; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_75; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_76; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_77; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_78; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_79; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_80; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_81; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_82; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_83; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_84; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_85; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_86; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_87; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_88; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_89; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_90; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_91; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_92; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_93; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_94; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_95; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_0; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_1; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_2; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_3; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_4; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_5; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_6; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_7; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_8; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_9; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_10; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_11; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_12; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_13; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_14; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_15; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_parse_current_state; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 265:26]
  wire [1:0] pipe3to8_io_pipe_phv_in_next_processor_id; // @[matcher.scala 265:26]
  wire  pipe3to8_io_pipe_phv_in_next_config_id; // @[matcher.scala 265:26]
  wire  pipe3to8_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_0; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_1; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_2; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_3; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_4; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_5; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_6; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_7; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_8; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_9; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_10; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_11; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_12; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_13; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_14; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_15; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_16; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_17; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_18; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_19; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_20; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_21; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_22; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_23; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_24; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_25; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_26; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_27; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_28; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_29; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_30; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_31; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_32; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_33; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_34; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_35; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_36; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_37; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_38; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_39; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_40; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_41; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_42; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_43; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_44; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_45; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_46; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_47; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_48; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_49; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_50; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_51; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_52; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_53; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_54; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_55; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_56; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_57; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_58; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_59; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_60; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_61; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_62; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_63; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_64; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_65; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_66; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_67; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_68; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_69; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_70; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_71; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_72; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_73; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_74; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_75; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_76; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_77; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_78; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_79; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_80; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_81; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_82; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_83; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_84; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_85; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_86; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_87; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_88; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_89; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_90; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_91; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_92; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_93; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_94; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_95; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_0; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_1; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_2; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_3; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_4; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_5; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_6; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_7; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_8; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_9; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_10; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_11; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_12; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_13; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_14; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_15; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_parse_current_state; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 265:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 265:26]
  wire [1:0] pipe3to8_io_pipe_phv_out_next_processor_id; // @[matcher.scala 265:26]
  wire  pipe3to8_io_pipe_phv_out_next_config_id; // @[matcher.scala 265:26]
  wire  pipe3to8_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 265:26]
  wire  pipe3to8_io_mod_hash_depth_mod; // @[matcher.scala 265:26]
  wire  pipe3to8_io_mod_config_id; // @[matcher.scala 265:26]
  wire [2:0] pipe3to8_io_mod_hash_depth; // @[matcher.scala 265:26]
  wire [63:0] pipe3to8_io_key_in; // @[matcher.scala 265:26]
  wire [63:0] pipe3to8_io_key_out; // @[matcher.scala 265:26]
  wire [7:0] pipe3to8_io_hash_val; // @[matcher.scala 265:26]
  wire [2:0] pipe3to8_io_hash_val_cs; // @[matcher.scala 265:26]
  wire  pipe9_clock; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_0; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_1; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_2; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_3; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_4; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_5; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_6; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_7; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_8; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_9; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_10; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_11; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_12; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_13; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_14; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_15; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_16; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_17; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_18; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_19; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_20; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_21; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_22; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_23; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_24; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_25; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_26; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_27; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_28; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_29; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_30; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_31; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_32; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_33; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_34; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_35; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_36; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_37; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_38; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_39; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_40; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_41; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_42; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_43; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_44; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_45; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_46; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_47; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_48; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_49; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_50; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_51; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_52; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_53; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_54; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_55; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_56; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_57; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_58; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_59; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_60; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_61; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_62; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_63; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_64; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_65; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_66; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_67; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_68; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_69; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_70; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_71; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_72; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_73; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_74; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_75; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_76; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_77; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_78; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_79; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_80; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_81; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_82; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_83; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_84; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_85; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_86; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_87; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_88; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_89; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_90; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_91; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_92; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_93; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_94; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_95; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_0; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_1; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_2; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_3; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_4; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_5; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_6; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_7; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_8; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_9; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_10; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_11; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_12; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_13; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_14; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_15; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_parse_current_state; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 266:23]
  wire [1:0] pipe9_io_pipe_phv_in_next_processor_id; // @[matcher.scala 266:23]
  wire  pipe9_io_pipe_phv_in_next_config_id; // @[matcher.scala 266:23]
  wire  pipe9_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_0; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_1; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_2; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_3; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_4; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_5; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_6; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_7; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_8; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_9; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_10; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_11; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_12; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_13; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_14; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_15; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_16; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_17; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_18; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_19; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_20; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_21; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_22; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_23; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_24; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_25; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_26; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_27; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_28; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_29; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_30; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_31; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_32; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_33; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_34; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_35; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_36; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_37; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_38; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_39; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_40; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_41; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_42; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_43; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_44; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_45; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_46; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_47; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_48; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_49; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_50; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_51; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_52; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_53; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_54; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_55; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_56; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_57; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_58; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_59; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_60; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_61; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_62; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_63; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_64; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_65; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_66; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_67; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_68; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_69; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_70; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_71; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_72; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_73; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_74; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_75; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_76; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_77; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_78; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_79; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_80; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_81; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_82; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_83; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_84; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_85; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_86; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_87; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_88; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_89; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_90; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_91; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_92; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_93; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_94; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_95; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_0; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_1; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_2; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_3; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_4; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_5; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_6; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_7; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_8; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_9; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_10; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_11; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_12; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_13; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_14; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_15; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_parse_current_state; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 266:23]
  wire [15:0] pipe9_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 266:23]
  wire [1:0] pipe9_io_pipe_phv_out_next_processor_id; // @[matcher.scala 266:23]
  wire  pipe9_io_pipe_phv_out_next_config_id; // @[matcher.scala 266:23]
  wire  pipe9_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 266:23]
  wire [3:0] pipe9_io_table_config_0_table_width; // @[matcher.scala 266:23]
  wire [3:0] pipe9_io_table_config_0_table_depth; // @[matcher.scala 266:23]
  wire [3:0] pipe9_io_table_config_1_table_width; // @[matcher.scala 266:23]
  wire [3:0] pipe9_io_table_config_1_table_depth; // @[matcher.scala 266:23]
  wire [63:0] pipe9_io_key_in; // @[matcher.scala 266:23]
  wire [63:0] pipe9_io_key_out; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_addr_in; // @[matcher.scala 266:23]
  wire [7:0] pipe9_io_addr_out; // @[matcher.scala 266:23]
  wire [2:0] pipe9_io_cs_in; // @[matcher.scala 266:23]
  wire [2:0] pipe9_io_cs_out; // @[matcher.scala 266:23]
  wire  pipe9_io_cs_vec_out_0; // @[matcher.scala 266:23]
  wire  pipe9_io_cs_vec_out_1; // @[matcher.scala 266:23]
  wire  pipe9_io_cs_vec_out_2; // @[matcher.scala 266:23]
  wire  pipe9_io_cs_vec_out_3; // @[matcher.scala 266:23]
  wire  pipe9_io_cs_vec_out_4; // @[matcher.scala 266:23]
  wire  pipe9_io_cs_vec_out_5; // @[matcher.scala 266:23]
  wire  pipe9_io_cs_vec_out_6; // @[matcher.scala 266:23]
  wire  pipe9_io_cs_vec_out_7; // @[matcher.scala 266:23]
  wire  pipe10_clock; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_0; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_1; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_2; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_3; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_4; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_5; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_6; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_7; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_8; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_9; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_10; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_11; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_12; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_13; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_14; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_15; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_16; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_17; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_18; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_19; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_20; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_21; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_22; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_23; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_24; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_25; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_26; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_27; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_28; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_29; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_30; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_31; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_32; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_33; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_34; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_35; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_36; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_37; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_38; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_39; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_40; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_41; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_42; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_43; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_44; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_45; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_46; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_47; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_48; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_49; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_50; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_51; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_52; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_53; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_54; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_55; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_56; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_57; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_58; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_59; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_60; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_61; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_62; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_63; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_64; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_65; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_66; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_67; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_68; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_69; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_70; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_71; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_72; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_73; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_74; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_75; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_76; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_77; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_78; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_79; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_80; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_81; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_82; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_83; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_84; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_85; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_86; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_87; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_88; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_89; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_90; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_91; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_92; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_93; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_94; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_95; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_0; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_1; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_2; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_3; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_4; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_5; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_6; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_7; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_8; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_9; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_10; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_11; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_12; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_13; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_14; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_15; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_parse_current_state; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 267:24]
  wire [1:0] pipe10_io_pipe_phv_in_next_processor_id; // @[matcher.scala 267:24]
  wire  pipe10_io_pipe_phv_in_next_config_id; // @[matcher.scala 267:24]
  wire  pipe10_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_0; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_1; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_2; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_3; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_4; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_5; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_6; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_7; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_8; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_9; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_10; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_11; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_12; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_13; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_14; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_15; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_16; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_17; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_18; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_19; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_20; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_21; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_22; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_23; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_24; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_25; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_26; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_27; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_28; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_29; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_30; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_31; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_32; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_33; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_34; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_35; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_36; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_37; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_38; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_39; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_40; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_41; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_42; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_43; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_44; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_45; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_46; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_47; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_48; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_49; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_50; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_51; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_52; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_53; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_54; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_55; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_56; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_57; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_58; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_59; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_60; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_61; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_62; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_63; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_64; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_65; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_66; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_67; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_68; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_69; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_70; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_71; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_72; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_73; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_74; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_75; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_76; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_77; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_78; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_79; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_80; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_81; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_82; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_83; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_84; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_85; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_86; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_87; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_88; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_89; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_90; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_91; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_92; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_93; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_94; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_95; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_0; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_1; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_2; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_3; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_4; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_5; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_6; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_7; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_8; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_9; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_10; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_11; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_12; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_13; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_14; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_15; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_parse_current_state; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 267:24]
  wire [15:0] pipe10_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 267:24]
  wire [1:0] pipe10_io_pipe_phv_out_next_processor_id; // @[matcher.scala 267:24]
  wire  pipe10_io_pipe_phv_out_next_config_id; // @[matcher.scala 267:24]
  wire  pipe10_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 267:24]
  wire [63:0] pipe10_io_key_in; // @[matcher.scala 267:24]
  wire [63:0] pipe10_io_key_out; // @[matcher.scala 267:24]
  wire [2:0] pipe10_io_cs_in; // @[matcher.scala 267:24]
  wire [2:0] pipe10_io_cs_out; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_addr_in; // @[matcher.scala 267:24]
  wire  pipe10_io_cs_vec_in_0; // @[matcher.scala 267:24]
  wire  pipe10_io_cs_vec_in_1; // @[matcher.scala 267:24]
  wire  pipe10_io_cs_vec_in_2; // @[matcher.scala 267:24]
  wire  pipe10_io_cs_vec_in_3; // @[matcher.scala 267:24]
  wire  pipe10_io_cs_vec_in_4; // @[matcher.scala 267:24]
  wire  pipe10_io_cs_vec_in_5; // @[matcher.scala 267:24]
  wire  pipe10_io_cs_vec_in_6; // @[matcher.scala 267:24]
  wire  pipe10_io_cs_vec_in_7; // @[matcher.scala 267:24]
  wire [63:0] pipe10_io_data_out_0; // @[matcher.scala 267:24]
  wire [63:0] pipe10_io_data_out_1; // @[matcher.scala 267:24]
  wire [63:0] pipe10_io_data_out_2; // @[matcher.scala 267:24]
  wire [63:0] pipe10_io_data_out_3; // @[matcher.scala 267:24]
  wire [63:0] pipe10_io_data_out_4; // @[matcher.scala 267:24]
  wire [63:0] pipe10_io_data_out_5; // @[matcher.scala 267:24]
  wire [63:0] pipe10_io_data_out_6; // @[matcher.scala 267:24]
  wire [63:0] pipe10_io_data_out_7; // @[matcher.scala 267:24]
  wire  pipe10_io_mem_cluster_0_en; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_mem_cluster_0_addr; // @[matcher.scala 267:24]
  wire [63:0] pipe10_io_mem_cluster_0_data; // @[matcher.scala 267:24]
  wire  pipe10_io_mem_cluster_1_en; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_mem_cluster_1_addr; // @[matcher.scala 267:24]
  wire [63:0] pipe10_io_mem_cluster_1_data; // @[matcher.scala 267:24]
  wire  pipe10_io_mem_cluster_2_en; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_mem_cluster_2_addr; // @[matcher.scala 267:24]
  wire [63:0] pipe10_io_mem_cluster_2_data; // @[matcher.scala 267:24]
  wire  pipe10_io_mem_cluster_3_en; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_mem_cluster_3_addr; // @[matcher.scala 267:24]
  wire [63:0] pipe10_io_mem_cluster_3_data; // @[matcher.scala 267:24]
  wire  pipe10_io_mem_cluster_4_en; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_mem_cluster_4_addr; // @[matcher.scala 267:24]
  wire [63:0] pipe10_io_mem_cluster_4_data; // @[matcher.scala 267:24]
  wire  pipe10_io_mem_cluster_5_en; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_mem_cluster_5_addr; // @[matcher.scala 267:24]
  wire [63:0] pipe10_io_mem_cluster_5_data; // @[matcher.scala 267:24]
  wire  pipe10_io_mem_cluster_6_en; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_mem_cluster_6_addr; // @[matcher.scala 267:24]
  wire [63:0] pipe10_io_mem_cluster_6_data; // @[matcher.scala 267:24]
  wire  pipe10_io_mem_cluster_7_en; // @[matcher.scala 267:24]
  wire [7:0] pipe10_io_mem_cluster_7_addr; // @[matcher.scala 267:24]
  wire [63:0] pipe10_io_mem_cluster_7_data; // @[matcher.scala 267:24]
  wire  pipe11_clock; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_0; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_1; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_2; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_3; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_4; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_5; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_6; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_7; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_8; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_9; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_10; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_11; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_12; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_13; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_14; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_15; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_16; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_17; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_18; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_19; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_20; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_21; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_22; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_23; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_24; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_25; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_26; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_27; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_28; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_29; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_30; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_31; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_32; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_33; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_34; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_35; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_36; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_37; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_38; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_39; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_40; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_41; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_42; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_43; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_44; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_45; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_46; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_47; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_48; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_49; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_50; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_51; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_52; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_53; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_54; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_55; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_56; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_57; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_58; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_59; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_60; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_61; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_62; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_63; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_64; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_65; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_66; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_67; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_68; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_69; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_70; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_71; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_72; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_73; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_74; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_75; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_76; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_77; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_78; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_79; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_80; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_81; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_82; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_83; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_84; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_85; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_86; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_87; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_88; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_89; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_90; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_91; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_92; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_93; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_94; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_95; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_0; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_1; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_2; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_3; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_4; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_5; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_6; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_7; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_8; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_9; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_10; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_11; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_12; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_13; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_14; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_15; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_parse_current_state; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 268:24]
  wire [1:0] pipe11_io_pipe_phv_in_next_processor_id; // @[matcher.scala 268:24]
  wire  pipe11_io_pipe_phv_in_next_config_id; // @[matcher.scala 268:24]
  wire  pipe11_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_0; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_1; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_2; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_3; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_4; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_5; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_6; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_7; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_8; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_9; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_10; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_11; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_12; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_13; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_14; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_15; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_16; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_17; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_18; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_19; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_20; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_21; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_22; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_23; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_24; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_25; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_26; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_27; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_28; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_29; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_30; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_31; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_32; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_33; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_34; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_35; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_36; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_37; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_38; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_39; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_40; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_41; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_42; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_43; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_44; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_45; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_46; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_47; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_48; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_49; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_50; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_51; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_52; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_53; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_54; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_55; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_56; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_57; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_58; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_59; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_60; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_61; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_62; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_63; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_64; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_65; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_66; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_67; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_68; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_69; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_70; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_71; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_72; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_73; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_74; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_75; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_76; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_77; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_78; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_79; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_80; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_81; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_82; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_83; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_84; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_85; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_86; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_87; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_88; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_89; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_90; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_91; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_92; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_93; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_94; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_95; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_0; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_1; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_2; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_3; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_4; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_5; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_6; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_7; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_8; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_9; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_10; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_11; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_12; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_13; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_14; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_15; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_parse_current_state; // @[matcher.scala 268:24]
  wire [7:0] pipe11_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 268:24]
  wire [15:0] pipe11_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 268:24]
  wire [1:0] pipe11_io_pipe_phv_out_next_processor_id; // @[matcher.scala 268:24]
  wire  pipe11_io_pipe_phv_out_next_config_id; // @[matcher.scala 268:24]
  wire  pipe11_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 268:24]
  wire [3:0] pipe11_io_table_config_0_table_width; // @[matcher.scala 268:24]
  wire [3:0] pipe11_io_table_config_0_table_depth; // @[matcher.scala 268:24]
  wire [3:0] pipe11_io_table_config_1_table_width; // @[matcher.scala 268:24]
  wire [3:0] pipe11_io_table_config_1_table_depth; // @[matcher.scala 268:24]
  wire [63:0] pipe11_io_key_in; // @[matcher.scala 268:24]
  wire [63:0] pipe11_io_key_out; // @[matcher.scala 268:24]
  wire [2:0] pipe11_io_cs_in; // @[matcher.scala 268:24]
  wire [63:0] pipe11_io_data_in_0; // @[matcher.scala 268:24]
  wire [63:0] pipe11_io_data_in_1; // @[matcher.scala 268:24]
  wire [63:0] pipe11_io_data_in_2; // @[matcher.scala 268:24]
  wire [63:0] pipe11_io_data_in_3; // @[matcher.scala 268:24]
  wire [63:0] pipe11_io_data_in_4; // @[matcher.scala 268:24]
  wire [63:0] pipe11_io_data_in_5; // @[matcher.scala 268:24]
  wire [63:0] pipe11_io_data_in_6; // @[matcher.scala 268:24]
  wire [63:0] pipe11_io_data_in_7; // @[matcher.scala 268:24]
  wire [127:0] pipe11_io_data_out; // @[matcher.scala 268:24]
  wire  pipe12_clock; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_0; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_1; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_2; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_3; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_4; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_5; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_6; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_7; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_8; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_9; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_10; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_11; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_12; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_13; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_14; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_15; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_16; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_17; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_18; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_19; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_20; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_21; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_22; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_23; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_24; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_25; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_26; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_27; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_28; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_29; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_30; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_31; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_32; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_33; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_34; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_35; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_36; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_37; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_38; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_39; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_40; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_41; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_42; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_43; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_44; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_45; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_46; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_47; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_48; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_49; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_50; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_51; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_52; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_53; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_54; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_55; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_56; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_57; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_58; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_59; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_60; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_61; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_62; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_63; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_64; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_65; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_66; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_67; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_68; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_69; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_70; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_71; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_72; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_73; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_74; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_75; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_76; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_77; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_78; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_79; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_80; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_81; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_82; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_83; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_84; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_85; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_86; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_87; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_88; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_89; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_90; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_91; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_92; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_93; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_94; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_95; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_0; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_1; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_2; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_3; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_4; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_5; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_6; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_7; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_8; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_9; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_10; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_11; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_12; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_13; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_14; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_15; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_parse_current_state; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 269:24]
  wire [1:0] pipe12_io_pipe_phv_in_next_processor_id; // @[matcher.scala 269:24]
  wire  pipe12_io_pipe_phv_in_next_config_id; // @[matcher.scala 269:24]
  wire  pipe12_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_0; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_1; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_2; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_3; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_4; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_5; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_6; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_7; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_8; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_9; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_10; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_11; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_12; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_13; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_14; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_15; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_16; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_17; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_18; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_19; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_20; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_21; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_22; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_23; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_24; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_25; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_26; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_27; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_28; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_29; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_30; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_31; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_32; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_33; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_34; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_35; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_36; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_37; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_38; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_39; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_40; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_41; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_42; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_43; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_44; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_45; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_46; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_47; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_48; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_49; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_50; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_51; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_52; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_53; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_54; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_55; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_56; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_57; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_58; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_59; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_60; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_61; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_62; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_63; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_64; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_65; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_66; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_67; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_68; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_69; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_70; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_71; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_72; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_73; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_74; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_75; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_76; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_77; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_78; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_79; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_80; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_81; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_82; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_83; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_84; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_85; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_86; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_87; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_88; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_89; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_90; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_91; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_92; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_93; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_94; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_95; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_0; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_1; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_2; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_3; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_4; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_5; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_6; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_7; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_8; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_9; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_10; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_11; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_12; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_13; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_14; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_15; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_parse_current_state; // @[matcher.scala 269:24]
  wire [7:0] pipe12_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 269:24]
  wire [15:0] pipe12_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 269:24]
  wire [1:0] pipe12_io_pipe_phv_out_next_processor_id; // @[matcher.scala 269:24]
  wire  pipe12_io_pipe_phv_out_next_config_id; // @[matcher.scala 269:24]
  wire  pipe12_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 269:24]
  wire [3:0] pipe12_io_key_config_0_key_length; // @[matcher.scala 269:24]
  wire [3:0] pipe12_io_key_config_1_key_length; // @[matcher.scala 269:24]
  wire [63:0] pipe12_io_key_in; // @[matcher.scala 269:24]
  wire [127:0] pipe12_io_data_in; // @[matcher.scala 269:24]
  wire  pipe12_io_hit; // @[matcher.scala 269:24]
  wire [63:0] pipe12_io_match_value; // @[matcher.scala 269:24]
  reg [7:0] key_config_0_header_id; // @[matcher.scala 17:25]
  reg [7:0] key_config_0_internal_offset; // @[matcher.scala 17:25]
  reg [3:0] key_config_0_key_length; // @[matcher.scala 17:25]
  reg [7:0] key_config_1_header_id; // @[matcher.scala 17:25]
  reg [7:0] key_config_1_internal_offset; // @[matcher.scala 17:25]
  reg [3:0] key_config_1_key_length; // @[matcher.scala 17:25]
  reg [3:0] table_config_0_table_width; // @[matcher.scala 18:27]
  reg [3:0] table_config_0_table_depth; // @[matcher.scala 18:27]
  reg [3:0] table_config_1_table_width; // @[matcher.scala 18:27]
  reg [3:0] table_config_1_table_depth; // @[matcher.scala 18:27]
  MatchGetOffset pipe1 ( // @[matcher.scala 263:23]
    .clock(pipe1_clock),
    .io_pipe_phv_in_data_0(pipe1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe1_io_pipe_phv_out_is_valid_processor),
    .io_key_config_0_header_id(pipe1_io_key_config_0_header_id),
    .io_key_config_0_internal_offset(pipe1_io_key_config_0_internal_offset),
    .io_key_config_1_header_id(pipe1_io_key_config_1_header_id),
    .io_key_config_1_internal_offset(pipe1_io_key_config_1_internal_offset),
    .io_key_offset(pipe1_io_key_offset)
  );
  MatchGetKey pipe2 ( // @[matcher.scala 264:23]
    .clock(pipe2_clock),
    .io_pipe_phv_in_data_0(pipe2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe2_io_pipe_phv_out_is_valid_processor),
    .io_key_config_0_key_length(pipe2_io_key_config_0_key_length),
    .io_key_config_1_key_length(pipe2_io_key_config_1_key_length),
    .io_key_offset(pipe2_io_key_offset),
    .io_match_key(pipe2_io_match_key)
  );
  Hash pipe3to8 ( // @[matcher.scala 265:26]
    .clock(pipe3to8_clock),
    .io_pipe_phv_in_data_0(pipe3to8_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe3to8_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe3to8_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe3to8_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe3to8_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe3to8_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe3to8_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe3to8_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe3to8_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe3to8_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe3to8_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe3to8_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe3to8_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe3to8_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe3to8_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe3to8_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe3to8_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe3to8_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe3to8_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe3to8_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe3to8_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe3to8_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe3to8_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe3to8_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe3to8_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe3to8_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe3to8_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe3to8_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe3to8_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe3to8_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe3to8_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe3to8_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe3to8_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe3to8_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe3to8_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe3to8_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe3to8_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe3to8_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe3to8_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe3to8_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe3to8_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe3to8_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe3to8_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe3to8_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe3to8_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe3to8_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe3to8_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe3to8_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe3to8_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe3to8_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe3to8_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe3to8_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe3to8_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe3to8_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe3to8_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe3to8_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe3to8_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe3to8_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe3to8_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe3to8_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe3to8_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe3to8_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe3to8_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe3to8_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe3to8_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe3to8_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe3to8_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe3to8_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe3to8_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe3to8_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe3to8_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe3to8_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe3to8_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe3to8_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe3to8_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe3to8_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe3to8_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe3to8_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe3to8_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe3to8_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe3to8_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe3to8_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe3to8_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe3to8_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe3to8_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe3to8_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe3to8_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe3to8_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe3to8_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe3to8_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe3to8_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe3to8_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe3to8_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe3to8_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe3to8_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe3to8_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe3to8_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe3to8_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe3to8_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe3to8_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe3to8_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe3to8_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe3to8_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe3to8_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe3to8_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe3to8_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe3to8_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe3to8_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe3to8_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe3to8_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe3to8_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe3to8_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe3to8_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe3to8_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe3to8_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe3to8_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe3to8_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe3to8_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe3to8_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe3to8_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe3to8_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe3to8_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe3to8_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe3to8_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe3to8_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe3to8_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe3to8_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe3to8_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe3to8_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe3to8_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe3to8_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe3to8_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe3to8_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe3to8_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe3to8_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe3to8_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe3to8_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe3to8_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe3to8_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe3to8_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe3to8_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe3to8_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe3to8_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe3to8_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe3to8_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe3to8_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe3to8_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe3to8_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe3to8_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe3to8_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe3to8_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe3to8_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe3to8_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe3to8_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe3to8_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe3to8_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe3to8_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe3to8_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe3to8_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe3to8_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe3to8_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe3to8_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe3to8_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe3to8_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe3to8_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe3to8_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe3to8_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe3to8_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe3to8_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe3to8_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe3to8_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe3to8_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe3to8_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe3to8_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe3to8_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe3to8_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe3to8_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe3to8_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe3to8_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe3to8_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe3to8_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe3to8_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe3to8_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe3to8_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe3to8_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe3to8_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe3to8_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe3to8_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe3to8_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe3to8_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe3to8_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe3to8_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe3to8_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe3to8_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe3to8_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe3to8_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe3to8_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe3to8_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe3to8_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe3to8_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe3to8_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe3to8_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe3to8_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe3to8_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe3to8_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe3to8_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe3to8_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe3to8_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe3to8_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe3to8_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe3to8_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe3to8_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe3to8_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe3to8_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe3to8_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe3to8_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe3to8_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe3to8_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe3to8_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe3to8_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe3to8_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe3to8_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe3to8_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe3to8_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe3to8_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe3to8_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe3to8_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe3to8_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe3to8_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe3to8_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe3to8_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe3to8_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe3to8_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe3to8_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe3to8_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe3to8_io_pipe_phv_out_is_valid_processor),
    .io_mod_hash_depth_mod(pipe3to8_io_mod_hash_depth_mod),
    .io_mod_config_id(pipe3to8_io_mod_config_id),
    .io_mod_hash_depth(pipe3to8_io_mod_hash_depth),
    .io_key_in(pipe3to8_io_key_in),
    .io_key_out(pipe3to8_io_key_out),
    .io_hash_val(pipe3to8_io_hash_val),
    .io_hash_val_cs(pipe3to8_io_hash_val_cs)
  );
  MatchGetCs pipe9 ( // @[matcher.scala 266:23]
    .clock(pipe9_clock),
    .io_pipe_phv_in_data_0(pipe9_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe9_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe9_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe9_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe9_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe9_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe9_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe9_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe9_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe9_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe9_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe9_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe9_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe9_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe9_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe9_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe9_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe9_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe9_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe9_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe9_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe9_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe9_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe9_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe9_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe9_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe9_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe9_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe9_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe9_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe9_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe9_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe9_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe9_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe9_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe9_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe9_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe9_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe9_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe9_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe9_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe9_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe9_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe9_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe9_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe9_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe9_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe9_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe9_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe9_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe9_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe9_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe9_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe9_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe9_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe9_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe9_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe9_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe9_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe9_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe9_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe9_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe9_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe9_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe9_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe9_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe9_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe9_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe9_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe9_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe9_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe9_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe9_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe9_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe9_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe9_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe9_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe9_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe9_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe9_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe9_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe9_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe9_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe9_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe9_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe9_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe9_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe9_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe9_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe9_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe9_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe9_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe9_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe9_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe9_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe9_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe9_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe9_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe9_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe9_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe9_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe9_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe9_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe9_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe9_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe9_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe9_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe9_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe9_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe9_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe9_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe9_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe9_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe9_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe9_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe9_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe9_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe9_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe9_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe9_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe9_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe9_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe9_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe9_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe9_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe9_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe9_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe9_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe9_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe9_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe9_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe9_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe9_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe9_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe9_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe9_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe9_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe9_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe9_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe9_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe9_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe9_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe9_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe9_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe9_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe9_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe9_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe9_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe9_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe9_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe9_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe9_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe9_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe9_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe9_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe9_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe9_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe9_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe9_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe9_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe9_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe9_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe9_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe9_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe9_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe9_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe9_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe9_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe9_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe9_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe9_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe9_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe9_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe9_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe9_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe9_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe9_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe9_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe9_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe9_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe9_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe9_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe9_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe9_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe9_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe9_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe9_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe9_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe9_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe9_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe9_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe9_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe9_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe9_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe9_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe9_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe9_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe9_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe9_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe9_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe9_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe9_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe9_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe9_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe9_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe9_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe9_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe9_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe9_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe9_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe9_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe9_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe9_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe9_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe9_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe9_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe9_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe9_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe9_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe9_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe9_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe9_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe9_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe9_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe9_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe9_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe9_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe9_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe9_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe9_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe9_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe9_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe9_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe9_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe9_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe9_io_pipe_phv_out_is_valid_processor),
    .io_table_config_0_table_width(pipe9_io_table_config_0_table_width),
    .io_table_config_0_table_depth(pipe9_io_table_config_0_table_depth),
    .io_table_config_1_table_width(pipe9_io_table_config_1_table_width),
    .io_table_config_1_table_depth(pipe9_io_table_config_1_table_depth),
    .io_key_in(pipe9_io_key_in),
    .io_key_out(pipe9_io_key_out),
    .io_addr_in(pipe9_io_addr_in),
    .io_addr_out(pipe9_io_addr_out),
    .io_cs_in(pipe9_io_cs_in),
    .io_cs_out(pipe9_io_cs_out),
    .io_cs_vec_out_0(pipe9_io_cs_vec_out_0),
    .io_cs_vec_out_1(pipe9_io_cs_vec_out_1),
    .io_cs_vec_out_2(pipe9_io_cs_vec_out_2),
    .io_cs_vec_out_3(pipe9_io_cs_vec_out_3),
    .io_cs_vec_out_4(pipe9_io_cs_vec_out_4),
    .io_cs_vec_out_5(pipe9_io_cs_vec_out_5),
    .io_cs_vec_out_6(pipe9_io_cs_vec_out_6),
    .io_cs_vec_out_7(pipe9_io_cs_vec_out_7)
  );
  MatchReadData pipe10 ( // @[matcher.scala 267:24]
    .clock(pipe10_clock),
    .io_pipe_phv_in_data_0(pipe10_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe10_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe10_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe10_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe10_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe10_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe10_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe10_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe10_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe10_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe10_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe10_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe10_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe10_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe10_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe10_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe10_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe10_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe10_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe10_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe10_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe10_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe10_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe10_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe10_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe10_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe10_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe10_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe10_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe10_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe10_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe10_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe10_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe10_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe10_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe10_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe10_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe10_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe10_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe10_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe10_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe10_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe10_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe10_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe10_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe10_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe10_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe10_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe10_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe10_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe10_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe10_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe10_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe10_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe10_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe10_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe10_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe10_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe10_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe10_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe10_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe10_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe10_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe10_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe10_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe10_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe10_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe10_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe10_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe10_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe10_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe10_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe10_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe10_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe10_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe10_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe10_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe10_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe10_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe10_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe10_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe10_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe10_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe10_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe10_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe10_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe10_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe10_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe10_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe10_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe10_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe10_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe10_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe10_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe10_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe10_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe10_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe10_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe10_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe10_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe10_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe10_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe10_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe10_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe10_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe10_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe10_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe10_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe10_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe10_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe10_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe10_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe10_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe10_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe10_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe10_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe10_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe10_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe10_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe10_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe10_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe10_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe10_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe10_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe10_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe10_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe10_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe10_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe10_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe10_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe10_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe10_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe10_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe10_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe10_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe10_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe10_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe10_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe10_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe10_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe10_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe10_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe10_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe10_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe10_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe10_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe10_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe10_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe10_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe10_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe10_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe10_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe10_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe10_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe10_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe10_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe10_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe10_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe10_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe10_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe10_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe10_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe10_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe10_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe10_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe10_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe10_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe10_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe10_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe10_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe10_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe10_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe10_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe10_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe10_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe10_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe10_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe10_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe10_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe10_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe10_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe10_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe10_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe10_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe10_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe10_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe10_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe10_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe10_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe10_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe10_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe10_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe10_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe10_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe10_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe10_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe10_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe10_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe10_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe10_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe10_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe10_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe10_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe10_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe10_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe10_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe10_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe10_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe10_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe10_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe10_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe10_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe10_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe10_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe10_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe10_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe10_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe10_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe10_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe10_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe10_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe10_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe10_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe10_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe10_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe10_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe10_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe10_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe10_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe10_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe10_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe10_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe10_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe10_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe10_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe10_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe10_io_key_in),
    .io_key_out(pipe10_io_key_out),
    .io_cs_in(pipe10_io_cs_in),
    .io_cs_out(pipe10_io_cs_out),
    .io_addr_in(pipe10_io_addr_in),
    .io_cs_vec_in_0(pipe10_io_cs_vec_in_0),
    .io_cs_vec_in_1(pipe10_io_cs_vec_in_1),
    .io_cs_vec_in_2(pipe10_io_cs_vec_in_2),
    .io_cs_vec_in_3(pipe10_io_cs_vec_in_3),
    .io_cs_vec_in_4(pipe10_io_cs_vec_in_4),
    .io_cs_vec_in_5(pipe10_io_cs_vec_in_5),
    .io_cs_vec_in_6(pipe10_io_cs_vec_in_6),
    .io_cs_vec_in_7(pipe10_io_cs_vec_in_7),
    .io_data_out_0(pipe10_io_data_out_0),
    .io_data_out_1(pipe10_io_data_out_1),
    .io_data_out_2(pipe10_io_data_out_2),
    .io_data_out_3(pipe10_io_data_out_3),
    .io_data_out_4(pipe10_io_data_out_4),
    .io_data_out_5(pipe10_io_data_out_5),
    .io_data_out_6(pipe10_io_data_out_6),
    .io_data_out_7(pipe10_io_data_out_7),
    .io_mem_cluster_0_en(pipe10_io_mem_cluster_0_en),
    .io_mem_cluster_0_addr(pipe10_io_mem_cluster_0_addr),
    .io_mem_cluster_0_data(pipe10_io_mem_cluster_0_data),
    .io_mem_cluster_1_en(pipe10_io_mem_cluster_1_en),
    .io_mem_cluster_1_addr(pipe10_io_mem_cluster_1_addr),
    .io_mem_cluster_1_data(pipe10_io_mem_cluster_1_data),
    .io_mem_cluster_2_en(pipe10_io_mem_cluster_2_en),
    .io_mem_cluster_2_addr(pipe10_io_mem_cluster_2_addr),
    .io_mem_cluster_2_data(pipe10_io_mem_cluster_2_data),
    .io_mem_cluster_3_en(pipe10_io_mem_cluster_3_en),
    .io_mem_cluster_3_addr(pipe10_io_mem_cluster_3_addr),
    .io_mem_cluster_3_data(pipe10_io_mem_cluster_3_data),
    .io_mem_cluster_4_en(pipe10_io_mem_cluster_4_en),
    .io_mem_cluster_4_addr(pipe10_io_mem_cluster_4_addr),
    .io_mem_cluster_4_data(pipe10_io_mem_cluster_4_data),
    .io_mem_cluster_5_en(pipe10_io_mem_cluster_5_en),
    .io_mem_cluster_5_addr(pipe10_io_mem_cluster_5_addr),
    .io_mem_cluster_5_data(pipe10_io_mem_cluster_5_data),
    .io_mem_cluster_6_en(pipe10_io_mem_cluster_6_en),
    .io_mem_cluster_6_addr(pipe10_io_mem_cluster_6_addr),
    .io_mem_cluster_6_data(pipe10_io_mem_cluster_6_data),
    .io_mem_cluster_7_en(pipe10_io_mem_cluster_7_en),
    .io_mem_cluster_7_addr(pipe10_io_mem_cluster_7_addr),
    .io_mem_cluster_7_data(pipe10_io_mem_cluster_7_data)
  );
  MatchDataReshape pipe11 ( // @[matcher.scala 268:24]
    .clock(pipe11_clock),
    .io_pipe_phv_in_data_0(pipe11_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe11_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe11_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe11_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe11_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe11_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe11_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe11_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe11_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe11_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe11_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe11_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe11_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe11_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe11_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe11_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe11_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe11_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe11_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe11_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe11_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe11_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe11_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe11_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe11_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe11_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe11_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe11_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe11_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe11_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe11_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe11_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe11_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe11_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe11_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe11_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe11_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe11_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe11_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe11_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe11_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe11_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe11_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe11_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe11_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe11_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe11_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe11_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe11_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe11_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe11_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe11_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe11_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe11_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe11_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe11_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe11_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe11_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe11_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe11_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe11_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe11_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe11_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe11_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe11_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe11_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe11_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe11_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe11_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe11_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe11_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe11_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe11_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe11_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe11_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe11_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe11_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe11_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe11_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe11_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe11_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe11_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe11_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe11_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe11_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe11_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe11_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe11_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe11_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe11_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe11_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe11_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe11_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe11_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe11_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe11_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe11_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe11_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe11_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe11_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe11_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe11_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe11_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe11_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe11_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe11_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe11_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe11_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe11_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe11_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe11_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe11_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe11_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe11_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe11_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe11_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe11_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe11_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe11_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe11_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe11_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe11_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe11_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe11_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe11_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe11_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe11_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe11_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe11_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe11_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe11_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe11_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe11_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe11_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe11_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe11_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe11_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe11_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe11_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe11_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe11_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe11_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe11_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe11_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe11_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe11_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe11_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe11_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe11_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe11_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe11_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe11_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe11_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe11_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe11_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe11_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe11_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe11_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe11_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe11_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe11_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe11_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe11_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe11_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe11_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe11_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe11_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe11_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe11_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe11_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe11_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe11_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe11_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe11_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe11_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe11_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe11_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe11_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe11_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe11_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe11_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe11_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe11_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe11_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe11_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe11_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe11_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe11_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe11_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe11_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe11_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe11_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe11_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe11_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe11_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe11_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe11_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe11_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe11_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe11_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe11_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe11_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe11_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe11_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe11_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe11_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe11_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe11_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe11_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe11_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe11_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe11_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe11_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe11_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe11_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe11_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe11_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe11_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe11_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe11_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe11_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe11_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe11_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe11_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe11_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe11_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe11_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe11_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe11_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe11_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe11_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe11_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe11_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe11_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe11_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe11_io_pipe_phv_out_is_valid_processor),
    .io_table_config_0_table_width(pipe11_io_table_config_0_table_width),
    .io_table_config_0_table_depth(pipe11_io_table_config_0_table_depth),
    .io_table_config_1_table_width(pipe11_io_table_config_1_table_width),
    .io_table_config_1_table_depth(pipe11_io_table_config_1_table_depth),
    .io_key_in(pipe11_io_key_in),
    .io_key_out(pipe11_io_key_out),
    .io_cs_in(pipe11_io_cs_in),
    .io_data_in_0(pipe11_io_data_in_0),
    .io_data_in_1(pipe11_io_data_in_1),
    .io_data_in_2(pipe11_io_data_in_2),
    .io_data_in_3(pipe11_io_data_in_3),
    .io_data_in_4(pipe11_io_data_in_4),
    .io_data_in_5(pipe11_io_data_in_5),
    .io_data_in_6(pipe11_io_data_in_6),
    .io_data_in_7(pipe11_io_data_in_7),
    .io_data_out(pipe11_io_data_out)
  );
  MatchResult pipe12 ( // @[matcher.scala 269:24]
    .clock(pipe12_clock),
    .io_pipe_phv_in_data_0(pipe12_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe12_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe12_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe12_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe12_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe12_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe12_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe12_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe12_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe12_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe12_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe12_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe12_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe12_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe12_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe12_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe12_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe12_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe12_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe12_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe12_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe12_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe12_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe12_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe12_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe12_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe12_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe12_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe12_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe12_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe12_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe12_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe12_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe12_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe12_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe12_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe12_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe12_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe12_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe12_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe12_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe12_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe12_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe12_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe12_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe12_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe12_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe12_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe12_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe12_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe12_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe12_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe12_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe12_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe12_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe12_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe12_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe12_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe12_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe12_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe12_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe12_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe12_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe12_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe12_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe12_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe12_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe12_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe12_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe12_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe12_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe12_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe12_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe12_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe12_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe12_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe12_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe12_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe12_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe12_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe12_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe12_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe12_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe12_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe12_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe12_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe12_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe12_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe12_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe12_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe12_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe12_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe12_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe12_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe12_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe12_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe12_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe12_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe12_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe12_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe12_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe12_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe12_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe12_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe12_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe12_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe12_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe12_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe12_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe12_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe12_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe12_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe12_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe12_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe12_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe12_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe12_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe12_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe12_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe12_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe12_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe12_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe12_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe12_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe12_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe12_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe12_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe12_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe12_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe12_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe12_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe12_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe12_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe12_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe12_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe12_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe12_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe12_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe12_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe12_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe12_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe12_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe12_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe12_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe12_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe12_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe12_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe12_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe12_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe12_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe12_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe12_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe12_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe12_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe12_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe12_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe12_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe12_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe12_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe12_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe12_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe12_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe12_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe12_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe12_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe12_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe12_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe12_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe12_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe12_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe12_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe12_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe12_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe12_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe12_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe12_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe12_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe12_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe12_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe12_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe12_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe12_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe12_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe12_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe12_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe12_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe12_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe12_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe12_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe12_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe12_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe12_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe12_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe12_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe12_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe12_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe12_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe12_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe12_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe12_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe12_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe12_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe12_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe12_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe12_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe12_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe12_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe12_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe12_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe12_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe12_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe12_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe12_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe12_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe12_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe12_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe12_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe12_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe12_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe12_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe12_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe12_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe12_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe12_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe12_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe12_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe12_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe12_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe12_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe12_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe12_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe12_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe12_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe12_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe12_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe12_io_pipe_phv_out_is_valid_processor),
    .io_key_config_0_key_length(pipe12_io_key_config_0_key_length),
    .io_key_config_1_key_length(pipe12_io_key_config_1_key_length),
    .io_key_in(pipe12_io_key_in),
    .io_data_in(pipe12_io_data_in),
    .io_hit(pipe12_io_hit),
    .io_match_value(pipe12_io_match_value)
  );
  assign io_pipe_phv_out_data_0 = pipe12_io_pipe_phv_out_data_0; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_1 = pipe12_io_pipe_phv_out_data_1; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_2 = pipe12_io_pipe_phv_out_data_2; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_3 = pipe12_io_pipe_phv_out_data_3; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_4 = pipe12_io_pipe_phv_out_data_4; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_5 = pipe12_io_pipe_phv_out_data_5; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_6 = pipe12_io_pipe_phv_out_data_6; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_7 = pipe12_io_pipe_phv_out_data_7; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_8 = pipe12_io_pipe_phv_out_data_8; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_9 = pipe12_io_pipe_phv_out_data_9; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_10 = pipe12_io_pipe_phv_out_data_10; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_11 = pipe12_io_pipe_phv_out_data_11; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_12 = pipe12_io_pipe_phv_out_data_12; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_13 = pipe12_io_pipe_phv_out_data_13; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_14 = pipe12_io_pipe_phv_out_data_14; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_15 = pipe12_io_pipe_phv_out_data_15; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_16 = pipe12_io_pipe_phv_out_data_16; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_17 = pipe12_io_pipe_phv_out_data_17; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_18 = pipe12_io_pipe_phv_out_data_18; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_19 = pipe12_io_pipe_phv_out_data_19; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_20 = pipe12_io_pipe_phv_out_data_20; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_21 = pipe12_io_pipe_phv_out_data_21; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_22 = pipe12_io_pipe_phv_out_data_22; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_23 = pipe12_io_pipe_phv_out_data_23; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_24 = pipe12_io_pipe_phv_out_data_24; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_25 = pipe12_io_pipe_phv_out_data_25; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_26 = pipe12_io_pipe_phv_out_data_26; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_27 = pipe12_io_pipe_phv_out_data_27; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_28 = pipe12_io_pipe_phv_out_data_28; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_29 = pipe12_io_pipe_phv_out_data_29; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_30 = pipe12_io_pipe_phv_out_data_30; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_31 = pipe12_io_pipe_phv_out_data_31; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_32 = pipe12_io_pipe_phv_out_data_32; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_33 = pipe12_io_pipe_phv_out_data_33; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_34 = pipe12_io_pipe_phv_out_data_34; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_35 = pipe12_io_pipe_phv_out_data_35; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_36 = pipe12_io_pipe_phv_out_data_36; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_37 = pipe12_io_pipe_phv_out_data_37; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_38 = pipe12_io_pipe_phv_out_data_38; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_39 = pipe12_io_pipe_phv_out_data_39; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_40 = pipe12_io_pipe_phv_out_data_40; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_41 = pipe12_io_pipe_phv_out_data_41; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_42 = pipe12_io_pipe_phv_out_data_42; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_43 = pipe12_io_pipe_phv_out_data_43; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_44 = pipe12_io_pipe_phv_out_data_44; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_45 = pipe12_io_pipe_phv_out_data_45; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_46 = pipe12_io_pipe_phv_out_data_46; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_47 = pipe12_io_pipe_phv_out_data_47; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_48 = pipe12_io_pipe_phv_out_data_48; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_49 = pipe12_io_pipe_phv_out_data_49; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_50 = pipe12_io_pipe_phv_out_data_50; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_51 = pipe12_io_pipe_phv_out_data_51; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_52 = pipe12_io_pipe_phv_out_data_52; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_53 = pipe12_io_pipe_phv_out_data_53; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_54 = pipe12_io_pipe_phv_out_data_54; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_55 = pipe12_io_pipe_phv_out_data_55; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_56 = pipe12_io_pipe_phv_out_data_56; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_57 = pipe12_io_pipe_phv_out_data_57; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_58 = pipe12_io_pipe_phv_out_data_58; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_59 = pipe12_io_pipe_phv_out_data_59; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_60 = pipe12_io_pipe_phv_out_data_60; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_61 = pipe12_io_pipe_phv_out_data_61; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_62 = pipe12_io_pipe_phv_out_data_62; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_63 = pipe12_io_pipe_phv_out_data_63; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_64 = pipe12_io_pipe_phv_out_data_64; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_65 = pipe12_io_pipe_phv_out_data_65; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_66 = pipe12_io_pipe_phv_out_data_66; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_67 = pipe12_io_pipe_phv_out_data_67; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_68 = pipe12_io_pipe_phv_out_data_68; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_69 = pipe12_io_pipe_phv_out_data_69; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_70 = pipe12_io_pipe_phv_out_data_70; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_71 = pipe12_io_pipe_phv_out_data_71; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_72 = pipe12_io_pipe_phv_out_data_72; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_73 = pipe12_io_pipe_phv_out_data_73; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_74 = pipe12_io_pipe_phv_out_data_74; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_75 = pipe12_io_pipe_phv_out_data_75; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_76 = pipe12_io_pipe_phv_out_data_76; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_77 = pipe12_io_pipe_phv_out_data_77; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_78 = pipe12_io_pipe_phv_out_data_78; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_79 = pipe12_io_pipe_phv_out_data_79; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_80 = pipe12_io_pipe_phv_out_data_80; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_81 = pipe12_io_pipe_phv_out_data_81; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_82 = pipe12_io_pipe_phv_out_data_82; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_83 = pipe12_io_pipe_phv_out_data_83; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_84 = pipe12_io_pipe_phv_out_data_84; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_85 = pipe12_io_pipe_phv_out_data_85; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_86 = pipe12_io_pipe_phv_out_data_86; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_87 = pipe12_io_pipe_phv_out_data_87; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_88 = pipe12_io_pipe_phv_out_data_88; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_89 = pipe12_io_pipe_phv_out_data_89; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_90 = pipe12_io_pipe_phv_out_data_90; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_91 = pipe12_io_pipe_phv_out_data_91; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_92 = pipe12_io_pipe_phv_out_data_92; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_93 = pipe12_io_pipe_phv_out_data_93; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_94 = pipe12_io_pipe_phv_out_data_94; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_data_95 = pipe12_io_pipe_phv_out_data_95; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_header_0 = pipe12_io_pipe_phv_out_header_0; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_header_1 = pipe12_io_pipe_phv_out_header_1; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_header_2 = pipe12_io_pipe_phv_out_header_2; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_header_3 = pipe12_io_pipe_phv_out_header_3; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_header_4 = pipe12_io_pipe_phv_out_header_4; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_header_5 = pipe12_io_pipe_phv_out_header_5; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_header_6 = pipe12_io_pipe_phv_out_header_6; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_header_7 = pipe12_io_pipe_phv_out_header_7; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_header_8 = pipe12_io_pipe_phv_out_header_8; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_header_9 = pipe12_io_pipe_phv_out_header_9; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_header_10 = pipe12_io_pipe_phv_out_header_10; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_header_11 = pipe12_io_pipe_phv_out_header_11; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_header_12 = pipe12_io_pipe_phv_out_header_12; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_header_13 = pipe12_io_pipe_phv_out_header_13; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_header_14 = pipe12_io_pipe_phv_out_header_14; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_header_15 = pipe12_io_pipe_phv_out_header_15; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_parse_current_state = pipe12_io_pipe_phv_out_parse_current_state; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_parse_current_offset = pipe12_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_parse_transition_field = pipe12_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_next_processor_id = pipe12_io_pipe_phv_out_next_processor_id; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_next_config_id = pipe12_io_pipe_phv_out_next_config_id; // @[matcher.scala 308:27]
  assign io_pipe_phv_out_is_valid_processor = pipe12_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 308:27]
  assign io_hit = pipe12_io_hit; // @[matcher.scala 309:27]
  assign io_match_value = pipe12_io_match_value; // @[matcher.scala 310:27]
  assign io_mem_cluster_0_en = pipe10_io_mem_cluster_0_en; // @[matcher.scala 295:27]
  assign io_mem_cluster_0_addr = pipe10_io_mem_cluster_0_addr; // @[matcher.scala 295:27]
  assign io_mem_cluster_1_en = pipe10_io_mem_cluster_1_en; // @[matcher.scala 295:27]
  assign io_mem_cluster_1_addr = pipe10_io_mem_cluster_1_addr; // @[matcher.scala 295:27]
  assign io_mem_cluster_2_en = pipe10_io_mem_cluster_2_en; // @[matcher.scala 295:27]
  assign io_mem_cluster_2_addr = pipe10_io_mem_cluster_2_addr; // @[matcher.scala 295:27]
  assign io_mem_cluster_3_en = pipe10_io_mem_cluster_3_en; // @[matcher.scala 295:27]
  assign io_mem_cluster_3_addr = pipe10_io_mem_cluster_3_addr; // @[matcher.scala 295:27]
  assign io_mem_cluster_4_en = pipe10_io_mem_cluster_4_en; // @[matcher.scala 295:27]
  assign io_mem_cluster_4_addr = pipe10_io_mem_cluster_4_addr; // @[matcher.scala 295:27]
  assign io_mem_cluster_5_en = pipe10_io_mem_cluster_5_en; // @[matcher.scala 295:27]
  assign io_mem_cluster_5_addr = pipe10_io_mem_cluster_5_addr; // @[matcher.scala 295:27]
  assign io_mem_cluster_6_en = pipe10_io_mem_cluster_6_en; // @[matcher.scala 295:27]
  assign io_mem_cluster_6_addr = pipe10_io_mem_cluster_6_addr; // @[matcher.scala 295:27]
  assign io_mem_cluster_7_en = pipe10_io_mem_cluster_7_en; // @[matcher.scala 295:27]
  assign io_mem_cluster_7_addr = pipe10_io_mem_cluster_7_addr; // @[matcher.scala 295:27]
  assign pipe1_clock = clock;
  assign pipe1_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[matcher.scala 271:26]
  assign pipe1_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[matcher.scala 271:26]
  assign pipe1_io_key_config_0_header_id = key_config_0_header_id; // @[matcher.scala 272:26]
  assign pipe1_io_key_config_0_internal_offset = key_config_0_internal_offset; // @[matcher.scala 272:26]
  assign pipe1_io_key_config_1_header_id = key_config_1_header_id; // @[matcher.scala 272:26]
  assign pipe1_io_key_config_1_internal_offset = key_config_1_internal_offset; // @[matcher.scala 272:26]
  assign pipe2_clock = clock;
  assign pipe2_io_pipe_phv_in_data_0 = pipe1_io_pipe_phv_out_data_0; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_1 = pipe1_io_pipe_phv_out_data_1; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_2 = pipe1_io_pipe_phv_out_data_2; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_3 = pipe1_io_pipe_phv_out_data_3; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_4 = pipe1_io_pipe_phv_out_data_4; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_5 = pipe1_io_pipe_phv_out_data_5; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_6 = pipe1_io_pipe_phv_out_data_6; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_7 = pipe1_io_pipe_phv_out_data_7; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_8 = pipe1_io_pipe_phv_out_data_8; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_9 = pipe1_io_pipe_phv_out_data_9; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_10 = pipe1_io_pipe_phv_out_data_10; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_11 = pipe1_io_pipe_phv_out_data_11; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_12 = pipe1_io_pipe_phv_out_data_12; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_13 = pipe1_io_pipe_phv_out_data_13; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_14 = pipe1_io_pipe_phv_out_data_14; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_15 = pipe1_io_pipe_phv_out_data_15; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_16 = pipe1_io_pipe_phv_out_data_16; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_17 = pipe1_io_pipe_phv_out_data_17; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_18 = pipe1_io_pipe_phv_out_data_18; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_19 = pipe1_io_pipe_phv_out_data_19; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_20 = pipe1_io_pipe_phv_out_data_20; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_21 = pipe1_io_pipe_phv_out_data_21; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_22 = pipe1_io_pipe_phv_out_data_22; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_23 = pipe1_io_pipe_phv_out_data_23; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_24 = pipe1_io_pipe_phv_out_data_24; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_25 = pipe1_io_pipe_phv_out_data_25; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_26 = pipe1_io_pipe_phv_out_data_26; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_27 = pipe1_io_pipe_phv_out_data_27; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_28 = pipe1_io_pipe_phv_out_data_28; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_29 = pipe1_io_pipe_phv_out_data_29; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_30 = pipe1_io_pipe_phv_out_data_30; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_31 = pipe1_io_pipe_phv_out_data_31; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_32 = pipe1_io_pipe_phv_out_data_32; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_33 = pipe1_io_pipe_phv_out_data_33; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_34 = pipe1_io_pipe_phv_out_data_34; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_35 = pipe1_io_pipe_phv_out_data_35; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_36 = pipe1_io_pipe_phv_out_data_36; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_37 = pipe1_io_pipe_phv_out_data_37; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_38 = pipe1_io_pipe_phv_out_data_38; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_39 = pipe1_io_pipe_phv_out_data_39; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_40 = pipe1_io_pipe_phv_out_data_40; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_41 = pipe1_io_pipe_phv_out_data_41; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_42 = pipe1_io_pipe_phv_out_data_42; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_43 = pipe1_io_pipe_phv_out_data_43; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_44 = pipe1_io_pipe_phv_out_data_44; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_45 = pipe1_io_pipe_phv_out_data_45; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_46 = pipe1_io_pipe_phv_out_data_46; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_47 = pipe1_io_pipe_phv_out_data_47; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_48 = pipe1_io_pipe_phv_out_data_48; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_49 = pipe1_io_pipe_phv_out_data_49; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_50 = pipe1_io_pipe_phv_out_data_50; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_51 = pipe1_io_pipe_phv_out_data_51; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_52 = pipe1_io_pipe_phv_out_data_52; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_53 = pipe1_io_pipe_phv_out_data_53; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_54 = pipe1_io_pipe_phv_out_data_54; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_55 = pipe1_io_pipe_phv_out_data_55; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_56 = pipe1_io_pipe_phv_out_data_56; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_57 = pipe1_io_pipe_phv_out_data_57; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_58 = pipe1_io_pipe_phv_out_data_58; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_59 = pipe1_io_pipe_phv_out_data_59; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_60 = pipe1_io_pipe_phv_out_data_60; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_61 = pipe1_io_pipe_phv_out_data_61; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_62 = pipe1_io_pipe_phv_out_data_62; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_63 = pipe1_io_pipe_phv_out_data_63; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_64 = pipe1_io_pipe_phv_out_data_64; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_65 = pipe1_io_pipe_phv_out_data_65; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_66 = pipe1_io_pipe_phv_out_data_66; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_67 = pipe1_io_pipe_phv_out_data_67; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_68 = pipe1_io_pipe_phv_out_data_68; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_69 = pipe1_io_pipe_phv_out_data_69; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_70 = pipe1_io_pipe_phv_out_data_70; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_71 = pipe1_io_pipe_phv_out_data_71; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_72 = pipe1_io_pipe_phv_out_data_72; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_73 = pipe1_io_pipe_phv_out_data_73; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_74 = pipe1_io_pipe_phv_out_data_74; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_75 = pipe1_io_pipe_phv_out_data_75; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_76 = pipe1_io_pipe_phv_out_data_76; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_77 = pipe1_io_pipe_phv_out_data_77; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_78 = pipe1_io_pipe_phv_out_data_78; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_79 = pipe1_io_pipe_phv_out_data_79; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_80 = pipe1_io_pipe_phv_out_data_80; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_81 = pipe1_io_pipe_phv_out_data_81; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_82 = pipe1_io_pipe_phv_out_data_82; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_83 = pipe1_io_pipe_phv_out_data_83; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_84 = pipe1_io_pipe_phv_out_data_84; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_85 = pipe1_io_pipe_phv_out_data_85; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_86 = pipe1_io_pipe_phv_out_data_86; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_87 = pipe1_io_pipe_phv_out_data_87; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_88 = pipe1_io_pipe_phv_out_data_88; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_89 = pipe1_io_pipe_phv_out_data_89; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_90 = pipe1_io_pipe_phv_out_data_90; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_91 = pipe1_io_pipe_phv_out_data_91; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_92 = pipe1_io_pipe_phv_out_data_92; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_93 = pipe1_io_pipe_phv_out_data_93; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_94 = pipe1_io_pipe_phv_out_data_94; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_data_95 = pipe1_io_pipe_phv_out_data_95; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_header_0 = pipe1_io_pipe_phv_out_header_0; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_header_1 = pipe1_io_pipe_phv_out_header_1; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_header_2 = pipe1_io_pipe_phv_out_header_2; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_header_3 = pipe1_io_pipe_phv_out_header_3; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_header_4 = pipe1_io_pipe_phv_out_header_4; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_header_5 = pipe1_io_pipe_phv_out_header_5; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_header_6 = pipe1_io_pipe_phv_out_header_6; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_header_7 = pipe1_io_pipe_phv_out_header_7; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_header_8 = pipe1_io_pipe_phv_out_header_8; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_header_9 = pipe1_io_pipe_phv_out_header_9; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_header_10 = pipe1_io_pipe_phv_out_header_10; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_header_11 = pipe1_io_pipe_phv_out_header_11; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_header_12 = pipe1_io_pipe_phv_out_header_12; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_header_13 = pipe1_io_pipe_phv_out_header_13; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_header_14 = pipe1_io_pipe_phv_out_header_14; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_header_15 = pipe1_io_pipe_phv_out_header_15; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_parse_current_state = pipe1_io_pipe_phv_out_parse_current_state; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_parse_current_offset = pipe1_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_parse_transition_field = pipe1_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_next_processor_id = pipe1_io_pipe_phv_out_next_processor_id; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_next_config_id = pipe1_io_pipe_phv_out_next_config_id; // @[matcher.scala 274:26]
  assign pipe2_io_pipe_phv_in_is_valid_processor = pipe1_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 274:26]
  assign pipe2_io_key_config_0_key_length = key_config_0_key_length; // @[matcher.scala 276:26]
  assign pipe2_io_key_config_1_key_length = key_config_1_key_length; // @[matcher.scala 276:26]
  assign pipe2_io_key_offset = pipe1_io_key_offset; // @[matcher.scala 275:26]
  assign pipe3to8_clock = clock;
  assign pipe3to8_io_pipe_phv_in_data_0 = pipe2_io_pipe_phv_out_data_0; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_1 = pipe2_io_pipe_phv_out_data_1; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_2 = pipe2_io_pipe_phv_out_data_2; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_3 = pipe2_io_pipe_phv_out_data_3; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_4 = pipe2_io_pipe_phv_out_data_4; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_5 = pipe2_io_pipe_phv_out_data_5; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_6 = pipe2_io_pipe_phv_out_data_6; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_7 = pipe2_io_pipe_phv_out_data_7; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_8 = pipe2_io_pipe_phv_out_data_8; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_9 = pipe2_io_pipe_phv_out_data_9; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_10 = pipe2_io_pipe_phv_out_data_10; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_11 = pipe2_io_pipe_phv_out_data_11; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_12 = pipe2_io_pipe_phv_out_data_12; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_13 = pipe2_io_pipe_phv_out_data_13; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_14 = pipe2_io_pipe_phv_out_data_14; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_15 = pipe2_io_pipe_phv_out_data_15; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_16 = pipe2_io_pipe_phv_out_data_16; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_17 = pipe2_io_pipe_phv_out_data_17; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_18 = pipe2_io_pipe_phv_out_data_18; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_19 = pipe2_io_pipe_phv_out_data_19; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_20 = pipe2_io_pipe_phv_out_data_20; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_21 = pipe2_io_pipe_phv_out_data_21; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_22 = pipe2_io_pipe_phv_out_data_22; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_23 = pipe2_io_pipe_phv_out_data_23; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_24 = pipe2_io_pipe_phv_out_data_24; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_25 = pipe2_io_pipe_phv_out_data_25; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_26 = pipe2_io_pipe_phv_out_data_26; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_27 = pipe2_io_pipe_phv_out_data_27; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_28 = pipe2_io_pipe_phv_out_data_28; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_29 = pipe2_io_pipe_phv_out_data_29; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_30 = pipe2_io_pipe_phv_out_data_30; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_31 = pipe2_io_pipe_phv_out_data_31; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_32 = pipe2_io_pipe_phv_out_data_32; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_33 = pipe2_io_pipe_phv_out_data_33; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_34 = pipe2_io_pipe_phv_out_data_34; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_35 = pipe2_io_pipe_phv_out_data_35; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_36 = pipe2_io_pipe_phv_out_data_36; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_37 = pipe2_io_pipe_phv_out_data_37; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_38 = pipe2_io_pipe_phv_out_data_38; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_39 = pipe2_io_pipe_phv_out_data_39; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_40 = pipe2_io_pipe_phv_out_data_40; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_41 = pipe2_io_pipe_phv_out_data_41; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_42 = pipe2_io_pipe_phv_out_data_42; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_43 = pipe2_io_pipe_phv_out_data_43; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_44 = pipe2_io_pipe_phv_out_data_44; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_45 = pipe2_io_pipe_phv_out_data_45; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_46 = pipe2_io_pipe_phv_out_data_46; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_47 = pipe2_io_pipe_phv_out_data_47; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_48 = pipe2_io_pipe_phv_out_data_48; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_49 = pipe2_io_pipe_phv_out_data_49; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_50 = pipe2_io_pipe_phv_out_data_50; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_51 = pipe2_io_pipe_phv_out_data_51; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_52 = pipe2_io_pipe_phv_out_data_52; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_53 = pipe2_io_pipe_phv_out_data_53; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_54 = pipe2_io_pipe_phv_out_data_54; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_55 = pipe2_io_pipe_phv_out_data_55; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_56 = pipe2_io_pipe_phv_out_data_56; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_57 = pipe2_io_pipe_phv_out_data_57; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_58 = pipe2_io_pipe_phv_out_data_58; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_59 = pipe2_io_pipe_phv_out_data_59; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_60 = pipe2_io_pipe_phv_out_data_60; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_61 = pipe2_io_pipe_phv_out_data_61; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_62 = pipe2_io_pipe_phv_out_data_62; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_63 = pipe2_io_pipe_phv_out_data_63; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_64 = pipe2_io_pipe_phv_out_data_64; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_65 = pipe2_io_pipe_phv_out_data_65; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_66 = pipe2_io_pipe_phv_out_data_66; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_67 = pipe2_io_pipe_phv_out_data_67; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_68 = pipe2_io_pipe_phv_out_data_68; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_69 = pipe2_io_pipe_phv_out_data_69; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_70 = pipe2_io_pipe_phv_out_data_70; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_71 = pipe2_io_pipe_phv_out_data_71; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_72 = pipe2_io_pipe_phv_out_data_72; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_73 = pipe2_io_pipe_phv_out_data_73; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_74 = pipe2_io_pipe_phv_out_data_74; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_75 = pipe2_io_pipe_phv_out_data_75; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_76 = pipe2_io_pipe_phv_out_data_76; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_77 = pipe2_io_pipe_phv_out_data_77; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_78 = pipe2_io_pipe_phv_out_data_78; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_79 = pipe2_io_pipe_phv_out_data_79; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_80 = pipe2_io_pipe_phv_out_data_80; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_81 = pipe2_io_pipe_phv_out_data_81; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_82 = pipe2_io_pipe_phv_out_data_82; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_83 = pipe2_io_pipe_phv_out_data_83; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_84 = pipe2_io_pipe_phv_out_data_84; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_85 = pipe2_io_pipe_phv_out_data_85; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_86 = pipe2_io_pipe_phv_out_data_86; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_87 = pipe2_io_pipe_phv_out_data_87; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_88 = pipe2_io_pipe_phv_out_data_88; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_89 = pipe2_io_pipe_phv_out_data_89; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_90 = pipe2_io_pipe_phv_out_data_90; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_91 = pipe2_io_pipe_phv_out_data_91; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_92 = pipe2_io_pipe_phv_out_data_92; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_93 = pipe2_io_pipe_phv_out_data_93; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_94 = pipe2_io_pipe_phv_out_data_94; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_data_95 = pipe2_io_pipe_phv_out_data_95; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_header_0 = pipe2_io_pipe_phv_out_header_0; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_header_1 = pipe2_io_pipe_phv_out_header_1; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_header_2 = pipe2_io_pipe_phv_out_header_2; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_header_3 = pipe2_io_pipe_phv_out_header_3; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_header_4 = pipe2_io_pipe_phv_out_header_4; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_header_5 = pipe2_io_pipe_phv_out_header_5; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_header_6 = pipe2_io_pipe_phv_out_header_6; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_header_7 = pipe2_io_pipe_phv_out_header_7; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_header_8 = pipe2_io_pipe_phv_out_header_8; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_header_9 = pipe2_io_pipe_phv_out_header_9; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_header_10 = pipe2_io_pipe_phv_out_header_10; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_header_11 = pipe2_io_pipe_phv_out_header_11; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_header_12 = pipe2_io_pipe_phv_out_header_12; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_header_13 = pipe2_io_pipe_phv_out_header_13; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_header_14 = pipe2_io_pipe_phv_out_header_14; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_header_15 = pipe2_io_pipe_phv_out_header_15; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_parse_current_state = pipe2_io_pipe_phv_out_parse_current_state; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_parse_current_offset = pipe2_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_parse_transition_field = pipe2_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_next_processor_id = pipe2_io_pipe_phv_out_next_processor_id; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_next_config_id = pipe2_io_pipe_phv_out_next_config_id; // @[matcher.scala 278:29]
  assign pipe3to8_io_pipe_phv_in_is_valid_processor = pipe2_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 278:29]
  assign pipe3to8_io_mod_hash_depth_mod = io_mod_en; // @[matcher.scala 279:36]
  assign pipe3to8_io_mod_config_id = io_mod_config_id; // @[matcher.scala 280:36]
  assign pipe3to8_io_mod_hash_depth = io_mod_table_mod_table_depth[2:0]; // @[matcher.scala 281:36]
  assign pipe3to8_io_key_in = pipe2_io_match_key; // @[matcher.scala 282:26]
  assign pipe9_clock = clock;
  assign pipe9_io_pipe_phv_in_data_0 = pipe3to8_io_pipe_phv_out_data_0; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_1 = pipe3to8_io_pipe_phv_out_data_1; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_2 = pipe3to8_io_pipe_phv_out_data_2; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_3 = pipe3to8_io_pipe_phv_out_data_3; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_4 = pipe3to8_io_pipe_phv_out_data_4; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_5 = pipe3to8_io_pipe_phv_out_data_5; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_6 = pipe3to8_io_pipe_phv_out_data_6; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_7 = pipe3to8_io_pipe_phv_out_data_7; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_8 = pipe3to8_io_pipe_phv_out_data_8; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_9 = pipe3to8_io_pipe_phv_out_data_9; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_10 = pipe3to8_io_pipe_phv_out_data_10; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_11 = pipe3to8_io_pipe_phv_out_data_11; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_12 = pipe3to8_io_pipe_phv_out_data_12; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_13 = pipe3to8_io_pipe_phv_out_data_13; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_14 = pipe3to8_io_pipe_phv_out_data_14; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_15 = pipe3to8_io_pipe_phv_out_data_15; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_16 = pipe3to8_io_pipe_phv_out_data_16; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_17 = pipe3to8_io_pipe_phv_out_data_17; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_18 = pipe3to8_io_pipe_phv_out_data_18; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_19 = pipe3to8_io_pipe_phv_out_data_19; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_20 = pipe3to8_io_pipe_phv_out_data_20; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_21 = pipe3to8_io_pipe_phv_out_data_21; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_22 = pipe3to8_io_pipe_phv_out_data_22; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_23 = pipe3to8_io_pipe_phv_out_data_23; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_24 = pipe3to8_io_pipe_phv_out_data_24; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_25 = pipe3to8_io_pipe_phv_out_data_25; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_26 = pipe3to8_io_pipe_phv_out_data_26; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_27 = pipe3to8_io_pipe_phv_out_data_27; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_28 = pipe3to8_io_pipe_phv_out_data_28; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_29 = pipe3to8_io_pipe_phv_out_data_29; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_30 = pipe3to8_io_pipe_phv_out_data_30; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_31 = pipe3to8_io_pipe_phv_out_data_31; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_32 = pipe3to8_io_pipe_phv_out_data_32; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_33 = pipe3to8_io_pipe_phv_out_data_33; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_34 = pipe3to8_io_pipe_phv_out_data_34; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_35 = pipe3to8_io_pipe_phv_out_data_35; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_36 = pipe3to8_io_pipe_phv_out_data_36; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_37 = pipe3to8_io_pipe_phv_out_data_37; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_38 = pipe3to8_io_pipe_phv_out_data_38; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_39 = pipe3to8_io_pipe_phv_out_data_39; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_40 = pipe3to8_io_pipe_phv_out_data_40; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_41 = pipe3to8_io_pipe_phv_out_data_41; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_42 = pipe3to8_io_pipe_phv_out_data_42; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_43 = pipe3to8_io_pipe_phv_out_data_43; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_44 = pipe3to8_io_pipe_phv_out_data_44; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_45 = pipe3to8_io_pipe_phv_out_data_45; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_46 = pipe3to8_io_pipe_phv_out_data_46; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_47 = pipe3to8_io_pipe_phv_out_data_47; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_48 = pipe3to8_io_pipe_phv_out_data_48; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_49 = pipe3to8_io_pipe_phv_out_data_49; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_50 = pipe3to8_io_pipe_phv_out_data_50; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_51 = pipe3to8_io_pipe_phv_out_data_51; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_52 = pipe3to8_io_pipe_phv_out_data_52; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_53 = pipe3to8_io_pipe_phv_out_data_53; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_54 = pipe3to8_io_pipe_phv_out_data_54; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_55 = pipe3to8_io_pipe_phv_out_data_55; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_56 = pipe3to8_io_pipe_phv_out_data_56; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_57 = pipe3to8_io_pipe_phv_out_data_57; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_58 = pipe3to8_io_pipe_phv_out_data_58; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_59 = pipe3to8_io_pipe_phv_out_data_59; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_60 = pipe3to8_io_pipe_phv_out_data_60; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_61 = pipe3to8_io_pipe_phv_out_data_61; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_62 = pipe3to8_io_pipe_phv_out_data_62; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_63 = pipe3to8_io_pipe_phv_out_data_63; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_64 = pipe3to8_io_pipe_phv_out_data_64; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_65 = pipe3to8_io_pipe_phv_out_data_65; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_66 = pipe3to8_io_pipe_phv_out_data_66; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_67 = pipe3to8_io_pipe_phv_out_data_67; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_68 = pipe3to8_io_pipe_phv_out_data_68; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_69 = pipe3to8_io_pipe_phv_out_data_69; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_70 = pipe3to8_io_pipe_phv_out_data_70; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_71 = pipe3to8_io_pipe_phv_out_data_71; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_72 = pipe3to8_io_pipe_phv_out_data_72; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_73 = pipe3to8_io_pipe_phv_out_data_73; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_74 = pipe3to8_io_pipe_phv_out_data_74; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_75 = pipe3to8_io_pipe_phv_out_data_75; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_76 = pipe3to8_io_pipe_phv_out_data_76; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_77 = pipe3to8_io_pipe_phv_out_data_77; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_78 = pipe3to8_io_pipe_phv_out_data_78; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_79 = pipe3to8_io_pipe_phv_out_data_79; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_80 = pipe3to8_io_pipe_phv_out_data_80; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_81 = pipe3to8_io_pipe_phv_out_data_81; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_82 = pipe3to8_io_pipe_phv_out_data_82; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_83 = pipe3to8_io_pipe_phv_out_data_83; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_84 = pipe3to8_io_pipe_phv_out_data_84; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_85 = pipe3to8_io_pipe_phv_out_data_85; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_86 = pipe3to8_io_pipe_phv_out_data_86; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_87 = pipe3to8_io_pipe_phv_out_data_87; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_88 = pipe3to8_io_pipe_phv_out_data_88; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_89 = pipe3to8_io_pipe_phv_out_data_89; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_90 = pipe3to8_io_pipe_phv_out_data_90; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_91 = pipe3to8_io_pipe_phv_out_data_91; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_92 = pipe3to8_io_pipe_phv_out_data_92; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_93 = pipe3to8_io_pipe_phv_out_data_93; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_94 = pipe3to8_io_pipe_phv_out_data_94; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_data_95 = pipe3to8_io_pipe_phv_out_data_95; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_header_0 = pipe3to8_io_pipe_phv_out_header_0; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_header_1 = pipe3to8_io_pipe_phv_out_header_1; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_header_2 = pipe3to8_io_pipe_phv_out_header_2; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_header_3 = pipe3to8_io_pipe_phv_out_header_3; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_header_4 = pipe3to8_io_pipe_phv_out_header_4; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_header_5 = pipe3to8_io_pipe_phv_out_header_5; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_header_6 = pipe3to8_io_pipe_phv_out_header_6; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_header_7 = pipe3to8_io_pipe_phv_out_header_7; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_header_8 = pipe3to8_io_pipe_phv_out_header_8; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_header_9 = pipe3to8_io_pipe_phv_out_header_9; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_header_10 = pipe3to8_io_pipe_phv_out_header_10; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_header_11 = pipe3to8_io_pipe_phv_out_header_11; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_header_12 = pipe3to8_io_pipe_phv_out_header_12; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_header_13 = pipe3to8_io_pipe_phv_out_header_13; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_header_14 = pipe3to8_io_pipe_phv_out_header_14; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_header_15 = pipe3to8_io_pipe_phv_out_header_15; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_parse_current_state = pipe3to8_io_pipe_phv_out_parse_current_state; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_parse_current_offset = pipe3to8_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_parse_transition_field = pipe3to8_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_next_processor_id = pipe3to8_io_pipe_phv_out_next_processor_id; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_next_config_id = pipe3to8_io_pipe_phv_out_next_config_id; // @[matcher.scala 284:27]
  assign pipe9_io_pipe_phv_in_is_valid_processor = pipe3to8_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 284:27]
  assign pipe9_io_table_config_0_table_width = table_config_0_table_width; // @[matcher.scala 288:27]
  assign pipe9_io_table_config_0_table_depth = table_config_0_table_depth; // @[matcher.scala 288:27]
  assign pipe9_io_table_config_1_table_width = table_config_1_table_width; // @[matcher.scala 288:27]
  assign pipe9_io_table_config_1_table_depth = table_config_1_table_depth; // @[matcher.scala 288:27]
  assign pipe9_io_key_in = pipe3to8_io_key_out; // @[matcher.scala 285:27]
  assign pipe9_io_addr_in = pipe3to8_io_hash_val; // @[matcher.scala 286:27]
  assign pipe9_io_cs_in = pipe3to8_io_hash_val_cs; // @[matcher.scala 287:27]
  assign pipe10_clock = clock;
  assign pipe10_io_pipe_phv_in_data_0 = pipe9_io_pipe_phv_out_data_0; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_1 = pipe9_io_pipe_phv_out_data_1; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_2 = pipe9_io_pipe_phv_out_data_2; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_3 = pipe9_io_pipe_phv_out_data_3; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_4 = pipe9_io_pipe_phv_out_data_4; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_5 = pipe9_io_pipe_phv_out_data_5; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_6 = pipe9_io_pipe_phv_out_data_6; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_7 = pipe9_io_pipe_phv_out_data_7; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_8 = pipe9_io_pipe_phv_out_data_8; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_9 = pipe9_io_pipe_phv_out_data_9; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_10 = pipe9_io_pipe_phv_out_data_10; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_11 = pipe9_io_pipe_phv_out_data_11; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_12 = pipe9_io_pipe_phv_out_data_12; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_13 = pipe9_io_pipe_phv_out_data_13; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_14 = pipe9_io_pipe_phv_out_data_14; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_15 = pipe9_io_pipe_phv_out_data_15; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_16 = pipe9_io_pipe_phv_out_data_16; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_17 = pipe9_io_pipe_phv_out_data_17; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_18 = pipe9_io_pipe_phv_out_data_18; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_19 = pipe9_io_pipe_phv_out_data_19; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_20 = pipe9_io_pipe_phv_out_data_20; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_21 = pipe9_io_pipe_phv_out_data_21; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_22 = pipe9_io_pipe_phv_out_data_22; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_23 = pipe9_io_pipe_phv_out_data_23; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_24 = pipe9_io_pipe_phv_out_data_24; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_25 = pipe9_io_pipe_phv_out_data_25; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_26 = pipe9_io_pipe_phv_out_data_26; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_27 = pipe9_io_pipe_phv_out_data_27; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_28 = pipe9_io_pipe_phv_out_data_28; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_29 = pipe9_io_pipe_phv_out_data_29; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_30 = pipe9_io_pipe_phv_out_data_30; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_31 = pipe9_io_pipe_phv_out_data_31; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_32 = pipe9_io_pipe_phv_out_data_32; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_33 = pipe9_io_pipe_phv_out_data_33; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_34 = pipe9_io_pipe_phv_out_data_34; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_35 = pipe9_io_pipe_phv_out_data_35; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_36 = pipe9_io_pipe_phv_out_data_36; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_37 = pipe9_io_pipe_phv_out_data_37; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_38 = pipe9_io_pipe_phv_out_data_38; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_39 = pipe9_io_pipe_phv_out_data_39; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_40 = pipe9_io_pipe_phv_out_data_40; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_41 = pipe9_io_pipe_phv_out_data_41; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_42 = pipe9_io_pipe_phv_out_data_42; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_43 = pipe9_io_pipe_phv_out_data_43; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_44 = pipe9_io_pipe_phv_out_data_44; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_45 = pipe9_io_pipe_phv_out_data_45; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_46 = pipe9_io_pipe_phv_out_data_46; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_47 = pipe9_io_pipe_phv_out_data_47; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_48 = pipe9_io_pipe_phv_out_data_48; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_49 = pipe9_io_pipe_phv_out_data_49; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_50 = pipe9_io_pipe_phv_out_data_50; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_51 = pipe9_io_pipe_phv_out_data_51; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_52 = pipe9_io_pipe_phv_out_data_52; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_53 = pipe9_io_pipe_phv_out_data_53; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_54 = pipe9_io_pipe_phv_out_data_54; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_55 = pipe9_io_pipe_phv_out_data_55; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_56 = pipe9_io_pipe_phv_out_data_56; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_57 = pipe9_io_pipe_phv_out_data_57; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_58 = pipe9_io_pipe_phv_out_data_58; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_59 = pipe9_io_pipe_phv_out_data_59; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_60 = pipe9_io_pipe_phv_out_data_60; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_61 = pipe9_io_pipe_phv_out_data_61; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_62 = pipe9_io_pipe_phv_out_data_62; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_63 = pipe9_io_pipe_phv_out_data_63; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_64 = pipe9_io_pipe_phv_out_data_64; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_65 = pipe9_io_pipe_phv_out_data_65; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_66 = pipe9_io_pipe_phv_out_data_66; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_67 = pipe9_io_pipe_phv_out_data_67; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_68 = pipe9_io_pipe_phv_out_data_68; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_69 = pipe9_io_pipe_phv_out_data_69; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_70 = pipe9_io_pipe_phv_out_data_70; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_71 = pipe9_io_pipe_phv_out_data_71; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_72 = pipe9_io_pipe_phv_out_data_72; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_73 = pipe9_io_pipe_phv_out_data_73; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_74 = pipe9_io_pipe_phv_out_data_74; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_75 = pipe9_io_pipe_phv_out_data_75; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_76 = pipe9_io_pipe_phv_out_data_76; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_77 = pipe9_io_pipe_phv_out_data_77; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_78 = pipe9_io_pipe_phv_out_data_78; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_79 = pipe9_io_pipe_phv_out_data_79; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_80 = pipe9_io_pipe_phv_out_data_80; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_81 = pipe9_io_pipe_phv_out_data_81; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_82 = pipe9_io_pipe_phv_out_data_82; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_83 = pipe9_io_pipe_phv_out_data_83; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_84 = pipe9_io_pipe_phv_out_data_84; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_85 = pipe9_io_pipe_phv_out_data_85; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_86 = pipe9_io_pipe_phv_out_data_86; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_87 = pipe9_io_pipe_phv_out_data_87; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_88 = pipe9_io_pipe_phv_out_data_88; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_89 = pipe9_io_pipe_phv_out_data_89; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_90 = pipe9_io_pipe_phv_out_data_90; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_91 = pipe9_io_pipe_phv_out_data_91; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_92 = pipe9_io_pipe_phv_out_data_92; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_93 = pipe9_io_pipe_phv_out_data_93; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_94 = pipe9_io_pipe_phv_out_data_94; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_data_95 = pipe9_io_pipe_phv_out_data_95; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_header_0 = pipe9_io_pipe_phv_out_header_0; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_header_1 = pipe9_io_pipe_phv_out_header_1; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_header_2 = pipe9_io_pipe_phv_out_header_2; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_header_3 = pipe9_io_pipe_phv_out_header_3; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_header_4 = pipe9_io_pipe_phv_out_header_4; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_header_5 = pipe9_io_pipe_phv_out_header_5; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_header_6 = pipe9_io_pipe_phv_out_header_6; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_header_7 = pipe9_io_pipe_phv_out_header_7; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_header_8 = pipe9_io_pipe_phv_out_header_8; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_header_9 = pipe9_io_pipe_phv_out_header_9; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_header_10 = pipe9_io_pipe_phv_out_header_10; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_header_11 = pipe9_io_pipe_phv_out_header_11; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_header_12 = pipe9_io_pipe_phv_out_header_12; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_header_13 = pipe9_io_pipe_phv_out_header_13; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_header_14 = pipe9_io_pipe_phv_out_header_14; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_header_15 = pipe9_io_pipe_phv_out_header_15; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_parse_current_state = pipe9_io_pipe_phv_out_parse_current_state; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_parse_current_offset = pipe9_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_parse_transition_field = pipe9_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_next_processor_id = pipe9_io_pipe_phv_out_next_processor_id; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_next_config_id = pipe9_io_pipe_phv_out_next_config_id; // @[matcher.scala 290:27]
  assign pipe10_io_pipe_phv_in_is_valid_processor = pipe9_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 290:27]
  assign pipe10_io_key_in = pipe9_io_key_out; // @[matcher.scala 291:27]
  assign pipe10_io_cs_in = pipe9_io_cs_out; // @[matcher.scala 292:27]
  assign pipe10_io_addr_in = pipe9_io_addr_out; // @[matcher.scala 293:27]
  assign pipe10_io_cs_vec_in_0 = pipe9_io_cs_vec_out_0; // @[matcher.scala 294:27]
  assign pipe10_io_cs_vec_in_1 = pipe9_io_cs_vec_out_1; // @[matcher.scala 294:27]
  assign pipe10_io_cs_vec_in_2 = pipe9_io_cs_vec_out_2; // @[matcher.scala 294:27]
  assign pipe10_io_cs_vec_in_3 = pipe9_io_cs_vec_out_3; // @[matcher.scala 294:27]
  assign pipe10_io_cs_vec_in_4 = pipe9_io_cs_vec_out_4; // @[matcher.scala 294:27]
  assign pipe10_io_cs_vec_in_5 = pipe9_io_cs_vec_out_5; // @[matcher.scala 294:27]
  assign pipe10_io_cs_vec_in_6 = pipe9_io_cs_vec_out_6; // @[matcher.scala 294:27]
  assign pipe10_io_cs_vec_in_7 = pipe9_io_cs_vec_out_7; // @[matcher.scala 294:27]
  assign pipe10_io_mem_cluster_0_data = io_mem_cluster_0_data; // @[matcher.scala 295:27]
  assign pipe10_io_mem_cluster_1_data = io_mem_cluster_1_data; // @[matcher.scala 295:27]
  assign pipe10_io_mem_cluster_2_data = io_mem_cluster_2_data; // @[matcher.scala 295:27]
  assign pipe10_io_mem_cluster_3_data = io_mem_cluster_3_data; // @[matcher.scala 295:27]
  assign pipe10_io_mem_cluster_4_data = io_mem_cluster_4_data; // @[matcher.scala 295:27]
  assign pipe10_io_mem_cluster_5_data = io_mem_cluster_5_data; // @[matcher.scala 295:27]
  assign pipe10_io_mem_cluster_6_data = io_mem_cluster_6_data; // @[matcher.scala 295:27]
  assign pipe10_io_mem_cluster_7_data = io_mem_cluster_7_data; // @[matcher.scala 295:27]
  assign pipe11_clock = clock;
  assign pipe11_io_pipe_phv_in_data_0 = pipe10_io_pipe_phv_out_data_0; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_1 = pipe10_io_pipe_phv_out_data_1; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_2 = pipe10_io_pipe_phv_out_data_2; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_3 = pipe10_io_pipe_phv_out_data_3; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_4 = pipe10_io_pipe_phv_out_data_4; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_5 = pipe10_io_pipe_phv_out_data_5; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_6 = pipe10_io_pipe_phv_out_data_6; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_7 = pipe10_io_pipe_phv_out_data_7; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_8 = pipe10_io_pipe_phv_out_data_8; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_9 = pipe10_io_pipe_phv_out_data_9; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_10 = pipe10_io_pipe_phv_out_data_10; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_11 = pipe10_io_pipe_phv_out_data_11; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_12 = pipe10_io_pipe_phv_out_data_12; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_13 = pipe10_io_pipe_phv_out_data_13; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_14 = pipe10_io_pipe_phv_out_data_14; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_15 = pipe10_io_pipe_phv_out_data_15; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_16 = pipe10_io_pipe_phv_out_data_16; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_17 = pipe10_io_pipe_phv_out_data_17; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_18 = pipe10_io_pipe_phv_out_data_18; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_19 = pipe10_io_pipe_phv_out_data_19; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_20 = pipe10_io_pipe_phv_out_data_20; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_21 = pipe10_io_pipe_phv_out_data_21; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_22 = pipe10_io_pipe_phv_out_data_22; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_23 = pipe10_io_pipe_phv_out_data_23; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_24 = pipe10_io_pipe_phv_out_data_24; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_25 = pipe10_io_pipe_phv_out_data_25; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_26 = pipe10_io_pipe_phv_out_data_26; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_27 = pipe10_io_pipe_phv_out_data_27; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_28 = pipe10_io_pipe_phv_out_data_28; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_29 = pipe10_io_pipe_phv_out_data_29; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_30 = pipe10_io_pipe_phv_out_data_30; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_31 = pipe10_io_pipe_phv_out_data_31; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_32 = pipe10_io_pipe_phv_out_data_32; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_33 = pipe10_io_pipe_phv_out_data_33; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_34 = pipe10_io_pipe_phv_out_data_34; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_35 = pipe10_io_pipe_phv_out_data_35; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_36 = pipe10_io_pipe_phv_out_data_36; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_37 = pipe10_io_pipe_phv_out_data_37; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_38 = pipe10_io_pipe_phv_out_data_38; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_39 = pipe10_io_pipe_phv_out_data_39; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_40 = pipe10_io_pipe_phv_out_data_40; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_41 = pipe10_io_pipe_phv_out_data_41; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_42 = pipe10_io_pipe_phv_out_data_42; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_43 = pipe10_io_pipe_phv_out_data_43; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_44 = pipe10_io_pipe_phv_out_data_44; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_45 = pipe10_io_pipe_phv_out_data_45; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_46 = pipe10_io_pipe_phv_out_data_46; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_47 = pipe10_io_pipe_phv_out_data_47; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_48 = pipe10_io_pipe_phv_out_data_48; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_49 = pipe10_io_pipe_phv_out_data_49; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_50 = pipe10_io_pipe_phv_out_data_50; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_51 = pipe10_io_pipe_phv_out_data_51; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_52 = pipe10_io_pipe_phv_out_data_52; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_53 = pipe10_io_pipe_phv_out_data_53; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_54 = pipe10_io_pipe_phv_out_data_54; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_55 = pipe10_io_pipe_phv_out_data_55; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_56 = pipe10_io_pipe_phv_out_data_56; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_57 = pipe10_io_pipe_phv_out_data_57; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_58 = pipe10_io_pipe_phv_out_data_58; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_59 = pipe10_io_pipe_phv_out_data_59; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_60 = pipe10_io_pipe_phv_out_data_60; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_61 = pipe10_io_pipe_phv_out_data_61; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_62 = pipe10_io_pipe_phv_out_data_62; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_63 = pipe10_io_pipe_phv_out_data_63; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_64 = pipe10_io_pipe_phv_out_data_64; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_65 = pipe10_io_pipe_phv_out_data_65; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_66 = pipe10_io_pipe_phv_out_data_66; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_67 = pipe10_io_pipe_phv_out_data_67; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_68 = pipe10_io_pipe_phv_out_data_68; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_69 = pipe10_io_pipe_phv_out_data_69; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_70 = pipe10_io_pipe_phv_out_data_70; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_71 = pipe10_io_pipe_phv_out_data_71; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_72 = pipe10_io_pipe_phv_out_data_72; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_73 = pipe10_io_pipe_phv_out_data_73; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_74 = pipe10_io_pipe_phv_out_data_74; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_75 = pipe10_io_pipe_phv_out_data_75; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_76 = pipe10_io_pipe_phv_out_data_76; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_77 = pipe10_io_pipe_phv_out_data_77; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_78 = pipe10_io_pipe_phv_out_data_78; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_79 = pipe10_io_pipe_phv_out_data_79; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_80 = pipe10_io_pipe_phv_out_data_80; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_81 = pipe10_io_pipe_phv_out_data_81; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_82 = pipe10_io_pipe_phv_out_data_82; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_83 = pipe10_io_pipe_phv_out_data_83; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_84 = pipe10_io_pipe_phv_out_data_84; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_85 = pipe10_io_pipe_phv_out_data_85; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_86 = pipe10_io_pipe_phv_out_data_86; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_87 = pipe10_io_pipe_phv_out_data_87; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_88 = pipe10_io_pipe_phv_out_data_88; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_89 = pipe10_io_pipe_phv_out_data_89; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_90 = pipe10_io_pipe_phv_out_data_90; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_91 = pipe10_io_pipe_phv_out_data_91; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_92 = pipe10_io_pipe_phv_out_data_92; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_93 = pipe10_io_pipe_phv_out_data_93; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_94 = pipe10_io_pipe_phv_out_data_94; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_data_95 = pipe10_io_pipe_phv_out_data_95; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_header_0 = pipe10_io_pipe_phv_out_header_0; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_header_1 = pipe10_io_pipe_phv_out_header_1; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_header_2 = pipe10_io_pipe_phv_out_header_2; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_header_3 = pipe10_io_pipe_phv_out_header_3; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_header_4 = pipe10_io_pipe_phv_out_header_4; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_header_5 = pipe10_io_pipe_phv_out_header_5; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_header_6 = pipe10_io_pipe_phv_out_header_6; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_header_7 = pipe10_io_pipe_phv_out_header_7; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_header_8 = pipe10_io_pipe_phv_out_header_8; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_header_9 = pipe10_io_pipe_phv_out_header_9; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_header_10 = pipe10_io_pipe_phv_out_header_10; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_header_11 = pipe10_io_pipe_phv_out_header_11; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_header_12 = pipe10_io_pipe_phv_out_header_12; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_header_13 = pipe10_io_pipe_phv_out_header_13; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_header_14 = pipe10_io_pipe_phv_out_header_14; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_header_15 = pipe10_io_pipe_phv_out_header_15; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_parse_current_state = pipe10_io_pipe_phv_out_parse_current_state; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_parse_current_offset = pipe10_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_parse_transition_field = pipe10_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_next_processor_id = pipe10_io_pipe_phv_out_next_processor_id; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_next_config_id = pipe10_io_pipe_phv_out_next_config_id; // @[matcher.scala 297:27]
  assign pipe11_io_pipe_phv_in_is_valid_processor = pipe10_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 297:27]
  assign pipe11_io_table_config_0_table_width = table_config_0_table_width; // @[matcher.scala 301:28]
  assign pipe11_io_table_config_0_table_depth = table_config_0_table_depth; // @[matcher.scala 301:28]
  assign pipe11_io_table_config_1_table_width = table_config_1_table_width; // @[matcher.scala 301:28]
  assign pipe11_io_table_config_1_table_depth = table_config_1_table_depth; // @[matcher.scala 301:28]
  assign pipe11_io_key_in = pipe10_io_key_out; // @[matcher.scala 298:27]
  assign pipe11_io_cs_in = pipe10_io_cs_out; // @[matcher.scala 299:27]
  assign pipe11_io_data_in_0 = pipe10_io_data_out_0; // @[matcher.scala 300:27]
  assign pipe11_io_data_in_1 = pipe10_io_data_out_1; // @[matcher.scala 300:27]
  assign pipe11_io_data_in_2 = pipe10_io_data_out_2; // @[matcher.scala 300:27]
  assign pipe11_io_data_in_3 = pipe10_io_data_out_3; // @[matcher.scala 300:27]
  assign pipe11_io_data_in_4 = pipe10_io_data_out_4; // @[matcher.scala 300:27]
  assign pipe11_io_data_in_5 = pipe10_io_data_out_5; // @[matcher.scala 300:27]
  assign pipe11_io_data_in_6 = pipe10_io_data_out_6; // @[matcher.scala 300:27]
  assign pipe11_io_data_in_7 = pipe10_io_data_out_7; // @[matcher.scala 300:27]
  assign pipe12_clock = clock;
  assign pipe12_io_pipe_phv_in_data_0 = pipe11_io_pipe_phv_out_data_0; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_1 = pipe11_io_pipe_phv_out_data_1; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_2 = pipe11_io_pipe_phv_out_data_2; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_3 = pipe11_io_pipe_phv_out_data_3; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_4 = pipe11_io_pipe_phv_out_data_4; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_5 = pipe11_io_pipe_phv_out_data_5; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_6 = pipe11_io_pipe_phv_out_data_6; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_7 = pipe11_io_pipe_phv_out_data_7; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_8 = pipe11_io_pipe_phv_out_data_8; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_9 = pipe11_io_pipe_phv_out_data_9; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_10 = pipe11_io_pipe_phv_out_data_10; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_11 = pipe11_io_pipe_phv_out_data_11; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_12 = pipe11_io_pipe_phv_out_data_12; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_13 = pipe11_io_pipe_phv_out_data_13; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_14 = pipe11_io_pipe_phv_out_data_14; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_15 = pipe11_io_pipe_phv_out_data_15; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_16 = pipe11_io_pipe_phv_out_data_16; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_17 = pipe11_io_pipe_phv_out_data_17; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_18 = pipe11_io_pipe_phv_out_data_18; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_19 = pipe11_io_pipe_phv_out_data_19; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_20 = pipe11_io_pipe_phv_out_data_20; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_21 = pipe11_io_pipe_phv_out_data_21; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_22 = pipe11_io_pipe_phv_out_data_22; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_23 = pipe11_io_pipe_phv_out_data_23; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_24 = pipe11_io_pipe_phv_out_data_24; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_25 = pipe11_io_pipe_phv_out_data_25; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_26 = pipe11_io_pipe_phv_out_data_26; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_27 = pipe11_io_pipe_phv_out_data_27; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_28 = pipe11_io_pipe_phv_out_data_28; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_29 = pipe11_io_pipe_phv_out_data_29; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_30 = pipe11_io_pipe_phv_out_data_30; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_31 = pipe11_io_pipe_phv_out_data_31; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_32 = pipe11_io_pipe_phv_out_data_32; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_33 = pipe11_io_pipe_phv_out_data_33; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_34 = pipe11_io_pipe_phv_out_data_34; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_35 = pipe11_io_pipe_phv_out_data_35; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_36 = pipe11_io_pipe_phv_out_data_36; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_37 = pipe11_io_pipe_phv_out_data_37; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_38 = pipe11_io_pipe_phv_out_data_38; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_39 = pipe11_io_pipe_phv_out_data_39; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_40 = pipe11_io_pipe_phv_out_data_40; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_41 = pipe11_io_pipe_phv_out_data_41; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_42 = pipe11_io_pipe_phv_out_data_42; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_43 = pipe11_io_pipe_phv_out_data_43; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_44 = pipe11_io_pipe_phv_out_data_44; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_45 = pipe11_io_pipe_phv_out_data_45; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_46 = pipe11_io_pipe_phv_out_data_46; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_47 = pipe11_io_pipe_phv_out_data_47; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_48 = pipe11_io_pipe_phv_out_data_48; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_49 = pipe11_io_pipe_phv_out_data_49; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_50 = pipe11_io_pipe_phv_out_data_50; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_51 = pipe11_io_pipe_phv_out_data_51; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_52 = pipe11_io_pipe_phv_out_data_52; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_53 = pipe11_io_pipe_phv_out_data_53; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_54 = pipe11_io_pipe_phv_out_data_54; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_55 = pipe11_io_pipe_phv_out_data_55; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_56 = pipe11_io_pipe_phv_out_data_56; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_57 = pipe11_io_pipe_phv_out_data_57; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_58 = pipe11_io_pipe_phv_out_data_58; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_59 = pipe11_io_pipe_phv_out_data_59; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_60 = pipe11_io_pipe_phv_out_data_60; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_61 = pipe11_io_pipe_phv_out_data_61; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_62 = pipe11_io_pipe_phv_out_data_62; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_63 = pipe11_io_pipe_phv_out_data_63; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_64 = pipe11_io_pipe_phv_out_data_64; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_65 = pipe11_io_pipe_phv_out_data_65; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_66 = pipe11_io_pipe_phv_out_data_66; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_67 = pipe11_io_pipe_phv_out_data_67; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_68 = pipe11_io_pipe_phv_out_data_68; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_69 = pipe11_io_pipe_phv_out_data_69; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_70 = pipe11_io_pipe_phv_out_data_70; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_71 = pipe11_io_pipe_phv_out_data_71; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_72 = pipe11_io_pipe_phv_out_data_72; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_73 = pipe11_io_pipe_phv_out_data_73; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_74 = pipe11_io_pipe_phv_out_data_74; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_75 = pipe11_io_pipe_phv_out_data_75; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_76 = pipe11_io_pipe_phv_out_data_76; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_77 = pipe11_io_pipe_phv_out_data_77; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_78 = pipe11_io_pipe_phv_out_data_78; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_79 = pipe11_io_pipe_phv_out_data_79; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_80 = pipe11_io_pipe_phv_out_data_80; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_81 = pipe11_io_pipe_phv_out_data_81; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_82 = pipe11_io_pipe_phv_out_data_82; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_83 = pipe11_io_pipe_phv_out_data_83; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_84 = pipe11_io_pipe_phv_out_data_84; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_85 = pipe11_io_pipe_phv_out_data_85; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_86 = pipe11_io_pipe_phv_out_data_86; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_87 = pipe11_io_pipe_phv_out_data_87; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_88 = pipe11_io_pipe_phv_out_data_88; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_89 = pipe11_io_pipe_phv_out_data_89; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_90 = pipe11_io_pipe_phv_out_data_90; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_91 = pipe11_io_pipe_phv_out_data_91; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_92 = pipe11_io_pipe_phv_out_data_92; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_93 = pipe11_io_pipe_phv_out_data_93; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_94 = pipe11_io_pipe_phv_out_data_94; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_data_95 = pipe11_io_pipe_phv_out_data_95; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_header_0 = pipe11_io_pipe_phv_out_header_0; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_header_1 = pipe11_io_pipe_phv_out_header_1; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_header_2 = pipe11_io_pipe_phv_out_header_2; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_header_3 = pipe11_io_pipe_phv_out_header_3; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_header_4 = pipe11_io_pipe_phv_out_header_4; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_header_5 = pipe11_io_pipe_phv_out_header_5; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_header_6 = pipe11_io_pipe_phv_out_header_6; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_header_7 = pipe11_io_pipe_phv_out_header_7; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_header_8 = pipe11_io_pipe_phv_out_header_8; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_header_9 = pipe11_io_pipe_phv_out_header_9; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_header_10 = pipe11_io_pipe_phv_out_header_10; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_header_11 = pipe11_io_pipe_phv_out_header_11; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_header_12 = pipe11_io_pipe_phv_out_header_12; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_header_13 = pipe11_io_pipe_phv_out_header_13; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_header_14 = pipe11_io_pipe_phv_out_header_14; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_header_15 = pipe11_io_pipe_phv_out_header_15; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_parse_current_state = pipe11_io_pipe_phv_out_parse_current_state; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_parse_current_offset = pipe11_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_parse_transition_field = pipe11_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_next_processor_id = pipe11_io_pipe_phv_out_next_processor_id; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_next_config_id = pipe11_io_pipe_phv_out_next_config_id; // @[matcher.scala 303:27]
  assign pipe12_io_pipe_phv_in_is_valid_processor = pipe11_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 303:27]
  assign pipe12_io_key_config_0_key_length = key_config_0_key_length; // @[matcher.scala 306:27]
  assign pipe12_io_key_config_1_key_length = key_config_1_key_length; // @[matcher.scala 306:27]
  assign pipe12_io_key_in = pipe11_io_key_out; // @[matcher.scala 304:27]
  assign pipe12_io_data_in = pipe11_io_data_out; // @[matcher.scala 305:27]
  always @(posedge clock) begin
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_0_header_id <= io_mod_key_mod_header_id; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_0_internal_offset <= io_mod_key_mod_internal_offset; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_0_key_length <= io_mod_key_mod_key_length; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_1_header_id <= io_mod_key_mod_header_id; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_1_internal_offset <= io_mod_key_mod_internal_offset; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_1_key_length <= io_mod_key_mod_key_length; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_table_width <= io_mod_table_mod_table_width; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_table_depth <= io_mod_table_mod_table_depth; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_table_width <= io_mod_table_mod_table_width; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_table_depth <= io_mod_table_mod_table_depth; // @[matcher.scala 22:40]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  key_config_0_header_id = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  key_config_0_internal_offset = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  key_config_0_key_length = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  key_config_1_header_id = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  key_config_1_internal_offset = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  key_config_1_key_length = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  table_config_0_table_width = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  table_config_0_table_depth = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  table_config_1_table_width = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  table_config_1_table_depth = _RAND_9[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
