module Parser(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  input         io_pipe_phv_in_valid,
  input         io_pipe_phv_in_last,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  output        io_pipe_phv_out_valid,
  output        io_pipe_phv_out_last
);
  wire  mau_0_clock; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_159; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_parse_transition_field; // @[parser.scala 21:25]
  wire  mau_0_io_pipe_phv_in_next_config_id; // @[parser.scala 21:25]
  wire  mau_0_io_pipe_phv_in_is_valid_processor; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_159; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_parse_transition_field; // @[parser.scala 21:25]
  wire  mau_0_io_pipe_phv_out_next_config_id; // @[parser.scala 21:25]
  wire  mau_0_io_pipe_phv_out_is_valid_processor; // @[parser.scala 21:25]
  wire  mau_1_clock; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_159; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_parse_transition_field; // @[parser.scala 21:25]
  wire  mau_1_io_pipe_phv_in_next_config_id; // @[parser.scala 21:25]
  wire  mau_1_io_pipe_phv_in_is_valid_processor; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_159; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_parse_transition_field; // @[parser.scala 21:25]
  wire  mau_1_io_pipe_phv_out_next_config_id; // @[parser.scala 21:25]
  wire  mau_1_io_pipe_phv_out_is_valid_processor; // @[parser.scala 21:25]
  wire  mau_2_clock; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_159; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_parse_transition_field; // @[parser.scala 21:25]
  wire  mau_2_io_pipe_phv_in_next_config_id; // @[parser.scala 21:25]
  wire  mau_2_io_pipe_phv_in_is_valid_processor; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_159; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_parse_transition_field; // @[parser.scala 21:25]
  wire  mau_2_io_pipe_phv_out_next_config_id; // @[parser.scala 21:25]
  wire  mau_2_io_pipe_phv_out_is_valid_processor; // @[parser.scala 21:25]
  wire  mau_3_clock; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_159; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_parse_transition_field; // @[parser.scala 21:25]
  wire  mau_3_io_pipe_phv_in_next_config_id; // @[parser.scala 21:25]
  wire  mau_3_io_pipe_phv_in_is_valid_processor; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_159; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_parse_transition_field; // @[parser.scala 21:25]
  wire  mau_3_io_pipe_phv_out_next_config_id; // @[parser.scala 21:25]
  wire  mau_3_io_pipe_phv_out_is_valid_processor; // @[parser.scala 21:25]
  ParseModule mau_0 ( // @[parser.scala 21:25]
    .clock(mau_0_clock),
    .io_pipe_phv_in_data_0(mau_0_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_0_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_0_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_0_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_0_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_0_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_0_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_0_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_0_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_0_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_0_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_0_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_0_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_0_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_0_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_0_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_0_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_0_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_0_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_0_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_0_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_0_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_0_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_0_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_0_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_0_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_0_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_0_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_0_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_0_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_0_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_0_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_0_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_0_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_0_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_0_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_0_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_0_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_0_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_0_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_0_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_0_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_0_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_0_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_0_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_0_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_0_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_0_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_0_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_0_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_0_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_0_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_0_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_0_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_0_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_0_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_0_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_0_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_0_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_0_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_0_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_0_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_0_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_0_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_0_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_0_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_0_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_0_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_0_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_0_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_0_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_0_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_0_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_0_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_0_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_0_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_0_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_0_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_0_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_0_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_0_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_0_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_0_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_0_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_0_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_0_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_0_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_0_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_0_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_0_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_0_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_0_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_0_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_0_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_0_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_0_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_0_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_0_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_0_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_0_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_0_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_0_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_0_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_0_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_0_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_0_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_0_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_0_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_0_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_0_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_0_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_0_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_0_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_0_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_0_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_0_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_0_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_0_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_0_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_0_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_0_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_0_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_0_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_0_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_0_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_0_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_0_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_0_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_0_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_0_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_0_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_0_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_0_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_0_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_0_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_0_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_0_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_0_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_0_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_0_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_0_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_0_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_0_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_0_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_0_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_0_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_0_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_0_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_0_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_0_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_0_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_0_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_0_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_0_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_0_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_0_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_0_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_0_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_0_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_0_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(mau_0_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_0_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_0_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_0_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_0_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_0_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_0_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_0_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_0_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_0_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_0_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_0_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_0_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_0_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_0_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_0_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_0_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_0_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_0_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_config_id(mau_0_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_0_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_0_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_0_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_0_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_0_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_0_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_0_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_0_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_0_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_0_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_0_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_0_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_0_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_0_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_0_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_0_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_0_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_0_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_0_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_0_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_0_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_0_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_0_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_0_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_0_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_0_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_0_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_0_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_0_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_0_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_0_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_0_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_0_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_0_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_0_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_0_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_0_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_0_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_0_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_0_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_0_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_0_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_0_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_0_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_0_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_0_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_0_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_0_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_0_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_0_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_0_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_0_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_0_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_0_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_0_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_0_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_0_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_0_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_0_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_0_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_0_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_0_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_0_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_0_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_0_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_0_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_0_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_0_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_0_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_0_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_0_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_0_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_0_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_0_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_0_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_0_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_0_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_0_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_0_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_0_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_0_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_0_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_0_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_0_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_0_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_0_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_0_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_0_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_0_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_0_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_0_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_0_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_0_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_0_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_0_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_0_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_0_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_0_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_0_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_0_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_0_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_0_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_0_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_0_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_0_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_0_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_0_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_0_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_0_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_0_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_0_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_0_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_0_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_0_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_0_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_0_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_0_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_0_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_0_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_0_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_0_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_0_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_0_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_0_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_0_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_0_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_0_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_0_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_0_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_0_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_0_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_0_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_0_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_0_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_0_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_0_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_0_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_0_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_0_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_0_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_0_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_0_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_0_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_0_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_0_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_0_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_0_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_0_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_0_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_0_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_0_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_0_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_0_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_0_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_0_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_0_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_0_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_0_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_0_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_0_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_0_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(mau_0_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_0_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_0_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_0_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_0_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_0_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_0_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_0_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_0_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_0_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_0_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_0_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_0_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_0_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_0_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_0_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_0_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_0_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_0_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_config_id(mau_0_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_0_io_pipe_phv_out_is_valid_processor)
  );
  ParseModule mau_1 ( // @[parser.scala 21:25]
    .clock(mau_1_clock),
    .io_pipe_phv_in_data_0(mau_1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(mau_1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_config_id(mau_1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(mau_1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_config_id(mau_1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_1_io_pipe_phv_out_is_valid_processor)
  );
  ParseModule mau_2 ( // @[parser.scala 21:25]
    .clock(mau_2_clock),
    .io_pipe_phv_in_data_0(mau_2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(mau_2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_config_id(mau_2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(mau_2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_config_id(mau_2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_2_io_pipe_phv_out_is_valid_processor)
  );
  ParseModule mau_3 ( // @[parser.scala 21:25]
    .clock(mau_3_clock),
    .io_pipe_phv_in_data_0(mau_3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_3_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_3_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_3_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_3_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_3_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_3_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_3_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_3_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_3_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_3_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_3_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_3_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_3_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_3_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_3_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_3_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_3_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_3_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_3_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_3_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_3_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_3_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_3_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_3_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_3_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_3_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_3_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_3_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_3_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_3_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_3_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_3_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_3_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_3_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_3_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_3_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_3_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_3_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_3_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_3_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_3_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_3_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_3_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_3_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_3_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_3_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_3_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_3_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_3_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_3_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_3_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_3_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_3_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_3_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_3_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_3_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_3_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_3_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_3_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_3_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_3_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_3_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_3_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_3_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(mau_3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_config_id(mau_3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_3_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_3_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_3_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_3_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_3_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_3_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_3_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_3_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_3_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_3_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_3_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_3_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_3_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_3_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_3_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_3_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_3_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_3_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_3_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_3_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_3_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_3_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_3_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_3_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_3_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_3_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_3_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_3_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_3_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_3_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_3_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_3_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_3_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_3_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_3_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_3_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_3_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_3_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_3_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_3_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_3_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_3_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_3_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_3_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_3_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_3_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_3_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_3_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_3_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_3_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_3_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_3_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_3_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_3_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_3_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_3_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_3_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_3_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_3_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_3_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_3_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_3_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_3_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_3_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(mau_3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_config_id(mau_3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_3_io_pipe_phv_out_is_valid_processor)
  );
  assign io_pipe_phv_out_data_0 = io_pipe_phv_in_data_0; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_1 = io_pipe_phv_in_data_1; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_2 = io_pipe_phv_in_data_2; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_3 = io_pipe_phv_in_data_3; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_4 = io_pipe_phv_in_data_4; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_5 = io_pipe_phv_in_data_5; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_6 = io_pipe_phv_in_data_6; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_7 = io_pipe_phv_in_data_7; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_8 = io_pipe_phv_in_data_8; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_9 = io_pipe_phv_in_data_9; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_10 = io_pipe_phv_in_data_10; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_11 = io_pipe_phv_in_data_11; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_12 = io_pipe_phv_in_data_12; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_13 = io_pipe_phv_in_data_13; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_14 = io_pipe_phv_in_data_14; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_15 = io_pipe_phv_in_data_15; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_16 = io_pipe_phv_in_data_16; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_17 = io_pipe_phv_in_data_17; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_18 = io_pipe_phv_in_data_18; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_19 = io_pipe_phv_in_data_19; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_20 = io_pipe_phv_in_data_20; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_21 = io_pipe_phv_in_data_21; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_22 = io_pipe_phv_in_data_22; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_23 = io_pipe_phv_in_data_23; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_24 = io_pipe_phv_in_data_24; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_25 = io_pipe_phv_in_data_25; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_26 = io_pipe_phv_in_data_26; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_27 = io_pipe_phv_in_data_27; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_28 = io_pipe_phv_in_data_28; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_29 = io_pipe_phv_in_data_29; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_30 = io_pipe_phv_in_data_30; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_31 = io_pipe_phv_in_data_31; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_32 = io_pipe_phv_in_data_32; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_33 = io_pipe_phv_in_data_33; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_34 = io_pipe_phv_in_data_34; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_35 = io_pipe_phv_in_data_35; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_36 = io_pipe_phv_in_data_36; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_37 = io_pipe_phv_in_data_37; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_38 = io_pipe_phv_in_data_38; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_39 = io_pipe_phv_in_data_39; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_40 = io_pipe_phv_in_data_40; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_41 = io_pipe_phv_in_data_41; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_42 = io_pipe_phv_in_data_42; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_43 = io_pipe_phv_in_data_43; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_44 = io_pipe_phv_in_data_44; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_45 = io_pipe_phv_in_data_45; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_46 = io_pipe_phv_in_data_46; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_47 = io_pipe_phv_in_data_47; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_48 = io_pipe_phv_in_data_48; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_49 = io_pipe_phv_in_data_49; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_50 = io_pipe_phv_in_data_50; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_51 = io_pipe_phv_in_data_51; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_52 = io_pipe_phv_in_data_52; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_53 = io_pipe_phv_in_data_53; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_54 = io_pipe_phv_in_data_54; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_55 = io_pipe_phv_in_data_55; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_56 = io_pipe_phv_in_data_56; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_57 = io_pipe_phv_in_data_57; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_58 = io_pipe_phv_in_data_58; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_59 = io_pipe_phv_in_data_59; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_60 = io_pipe_phv_in_data_60; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_61 = io_pipe_phv_in_data_61; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_62 = io_pipe_phv_in_data_62; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_63 = io_pipe_phv_in_data_63; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_64 = io_pipe_phv_in_data_64; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_65 = io_pipe_phv_in_data_65; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_66 = io_pipe_phv_in_data_66; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_67 = io_pipe_phv_in_data_67; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_68 = io_pipe_phv_in_data_68; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_69 = io_pipe_phv_in_data_69; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_70 = io_pipe_phv_in_data_70; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_71 = io_pipe_phv_in_data_71; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_72 = io_pipe_phv_in_data_72; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_73 = io_pipe_phv_in_data_73; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_74 = io_pipe_phv_in_data_74; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_75 = io_pipe_phv_in_data_75; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_76 = io_pipe_phv_in_data_76; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_77 = io_pipe_phv_in_data_77; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_78 = io_pipe_phv_in_data_78; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_79 = io_pipe_phv_in_data_79; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_80 = io_pipe_phv_in_data_80; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_81 = io_pipe_phv_in_data_81; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_82 = io_pipe_phv_in_data_82; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_83 = io_pipe_phv_in_data_83; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_84 = io_pipe_phv_in_data_84; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_85 = io_pipe_phv_in_data_85; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_86 = io_pipe_phv_in_data_86; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_87 = io_pipe_phv_in_data_87; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_88 = io_pipe_phv_in_data_88; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_89 = io_pipe_phv_in_data_89; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_90 = io_pipe_phv_in_data_90; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_91 = io_pipe_phv_in_data_91; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_92 = io_pipe_phv_in_data_92; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_93 = io_pipe_phv_in_data_93; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_94 = io_pipe_phv_in_data_94; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_95 = io_pipe_phv_in_data_95; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_96 = io_pipe_phv_in_data_96; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_97 = io_pipe_phv_in_data_97; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_98 = io_pipe_phv_in_data_98; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_99 = io_pipe_phv_in_data_99; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_100 = io_pipe_phv_in_data_100; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_101 = io_pipe_phv_in_data_101; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_102 = io_pipe_phv_in_data_102; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_103 = io_pipe_phv_in_data_103; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_104 = io_pipe_phv_in_data_104; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_105 = io_pipe_phv_in_data_105; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_106 = io_pipe_phv_in_data_106; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_107 = io_pipe_phv_in_data_107; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_108 = io_pipe_phv_in_data_108; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_109 = io_pipe_phv_in_data_109; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_110 = io_pipe_phv_in_data_110; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_111 = io_pipe_phv_in_data_111; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_112 = io_pipe_phv_in_data_112; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_113 = io_pipe_phv_in_data_113; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_114 = io_pipe_phv_in_data_114; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_115 = io_pipe_phv_in_data_115; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_116 = io_pipe_phv_in_data_116; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_117 = io_pipe_phv_in_data_117; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_118 = io_pipe_phv_in_data_118; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_119 = io_pipe_phv_in_data_119; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_120 = io_pipe_phv_in_data_120; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_121 = io_pipe_phv_in_data_121; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_122 = io_pipe_phv_in_data_122; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_123 = io_pipe_phv_in_data_123; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_124 = io_pipe_phv_in_data_124; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_125 = io_pipe_phv_in_data_125; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_126 = io_pipe_phv_in_data_126; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_127 = io_pipe_phv_in_data_127; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_128 = io_pipe_phv_in_data_128; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_129 = io_pipe_phv_in_data_129; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_130 = io_pipe_phv_in_data_130; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_131 = io_pipe_phv_in_data_131; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_132 = io_pipe_phv_in_data_132; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_133 = io_pipe_phv_in_data_133; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_134 = io_pipe_phv_in_data_134; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_135 = io_pipe_phv_in_data_135; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_136 = io_pipe_phv_in_data_136; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_137 = io_pipe_phv_in_data_137; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_138 = io_pipe_phv_in_data_138; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_139 = io_pipe_phv_in_data_139; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_140 = io_pipe_phv_in_data_140; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_141 = io_pipe_phv_in_data_141; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_142 = io_pipe_phv_in_data_142; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_143 = io_pipe_phv_in_data_143; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_144 = io_pipe_phv_in_data_144; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_145 = io_pipe_phv_in_data_145; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_146 = io_pipe_phv_in_data_146; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_147 = io_pipe_phv_in_data_147; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_148 = io_pipe_phv_in_data_148; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_149 = io_pipe_phv_in_data_149; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_150 = io_pipe_phv_in_data_150; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_151 = io_pipe_phv_in_data_151; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_152 = io_pipe_phv_in_data_152; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_153 = io_pipe_phv_in_data_153; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_154 = io_pipe_phv_in_data_154; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_155 = io_pipe_phv_in_data_155; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_156 = io_pipe_phv_in_data_156; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_157 = io_pipe_phv_in_data_157; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_158 = io_pipe_phv_in_data_158; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_159 = io_pipe_phv_in_data_159; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_0 = io_pipe_phv_in_header_0; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_1 = io_pipe_phv_in_header_1; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_2 = io_pipe_phv_in_header_2; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_3 = io_pipe_phv_in_header_3; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_4 = io_pipe_phv_in_header_4; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_5 = io_pipe_phv_in_header_5; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_6 = io_pipe_phv_in_header_6; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_7 = io_pipe_phv_in_header_7; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_8 = io_pipe_phv_in_header_8; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_9 = io_pipe_phv_in_header_9; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_10 = io_pipe_phv_in_header_10; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_11 = io_pipe_phv_in_header_11; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_12 = io_pipe_phv_in_header_12; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_13 = io_pipe_phv_in_header_13; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_14 = io_pipe_phv_in_header_14; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_15 = io_pipe_phv_in_header_15; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_parse_current_state = io_pipe_phv_in_parse_current_state; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_next_processor_id = io_pipe_phv_in_next_processor_id; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_next_config_id = io_pipe_phv_in_next_config_id; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_valid = io_pipe_phv_in_valid; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_last = io_pipe_phv_in_last; // @[parser.scala 33:62 parser.scala 34:35]
  assign mau_0_clock = clock;
  assign mau_0_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[parser.scala 30:35]
  assign mau_1_clock = clock;
  assign mau_1_io_pipe_phv_in_data_0 = mau_0_io_pipe_phv_out_data_0; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_1 = mau_0_io_pipe_phv_out_data_1; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_2 = mau_0_io_pipe_phv_out_data_2; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_3 = mau_0_io_pipe_phv_out_data_3; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_4 = mau_0_io_pipe_phv_out_data_4; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_5 = mau_0_io_pipe_phv_out_data_5; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_6 = mau_0_io_pipe_phv_out_data_6; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_7 = mau_0_io_pipe_phv_out_data_7; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_8 = mau_0_io_pipe_phv_out_data_8; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_9 = mau_0_io_pipe_phv_out_data_9; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_10 = mau_0_io_pipe_phv_out_data_10; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_11 = mau_0_io_pipe_phv_out_data_11; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_12 = mau_0_io_pipe_phv_out_data_12; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_13 = mau_0_io_pipe_phv_out_data_13; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_14 = mau_0_io_pipe_phv_out_data_14; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_15 = mau_0_io_pipe_phv_out_data_15; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_16 = mau_0_io_pipe_phv_out_data_16; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_17 = mau_0_io_pipe_phv_out_data_17; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_18 = mau_0_io_pipe_phv_out_data_18; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_19 = mau_0_io_pipe_phv_out_data_19; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_20 = mau_0_io_pipe_phv_out_data_20; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_21 = mau_0_io_pipe_phv_out_data_21; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_22 = mau_0_io_pipe_phv_out_data_22; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_23 = mau_0_io_pipe_phv_out_data_23; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_24 = mau_0_io_pipe_phv_out_data_24; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_25 = mau_0_io_pipe_phv_out_data_25; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_26 = mau_0_io_pipe_phv_out_data_26; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_27 = mau_0_io_pipe_phv_out_data_27; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_28 = mau_0_io_pipe_phv_out_data_28; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_29 = mau_0_io_pipe_phv_out_data_29; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_30 = mau_0_io_pipe_phv_out_data_30; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_31 = mau_0_io_pipe_phv_out_data_31; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_32 = mau_0_io_pipe_phv_out_data_32; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_33 = mau_0_io_pipe_phv_out_data_33; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_34 = mau_0_io_pipe_phv_out_data_34; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_35 = mau_0_io_pipe_phv_out_data_35; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_36 = mau_0_io_pipe_phv_out_data_36; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_37 = mau_0_io_pipe_phv_out_data_37; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_38 = mau_0_io_pipe_phv_out_data_38; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_39 = mau_0_io_pipe_phv_out_data_39; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_40 = mau_0_io_pipe_phv_out_data_40; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_41 = mau_0_io_pipe_phv_out_data_41; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_42 = mau_0_io_pipe_phv_out_data_42; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_43 = mau_0_io_pipe_phv_out_data_43; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_44 = mau_0_io_pipe_phv_out_data_44; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_45 = mau_0_io_pipe_phv_out_data_45; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_46 = mau_0_io_pipe_phv_out_data_46; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_47 = mau_0_io_pipe_phv_out_data_47; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_48 = mau_0_io_pipe_phv_out_data_48; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_49 = mau_0_io_pipe_phv_out_data_49; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_50 = mau_0_io_pipe_phv_out_data_50; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_51 = mau_0_io_pipe_phv_out_data_51; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_52 = mau_0_io_pipe_phv_out_data_52; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_53 = mau_0_io_pipe_phv_out_data_53; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_54 = mau_0_io_pipe_phv_out_data_54; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_55 = mau_0_io_pipe_phv_out_data_55; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_56 = mau_0_io_pipe_phv_out_data_56; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_57 = mau_0_io_pipe_phv_out_data_57; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_58 = mau_0_io_pipe_phv_out_data_58; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_59 = mau_0_io_pipe_phv_out_data_59; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_60 = mau_0_io_pipe_phv_out_data_60; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_61 = mau_0_io_pipe_phv_out_data_61; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_62 = mau_0_io_pipe_phv_out_data_62; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_63 = mau_0_io_pipe_phv_out_data_63; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_64 = mau_0_io_pipe_phv_out_data_64; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_65 = mau_0_io_pipe_phv_out_data_65; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_66 = mau_0_io_pipe_phv_out_data_66; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_67 = mau_0_io_pipe_phv_out_data_67; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_68 = mau_0_io_pipe_phv_out_data_68; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_69 = mau_0_io_pipe_phv_out_data_69; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_70 = mau_0_io_pipe_phv_out_data_70; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_71 = mau_0_io_pipe_phv_out_data_71; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_72 = mau_0_io_pipe_phv_out_data_72; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_73 = mau_0_io_pipe_phv_out_data_73; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_74 = mau_0_io_pipe_phv_out_data_74; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_75 = mau_0_io_pipe_phv_out_data_75; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_76 = mau_0_io_pipe_phv_out_data_76; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_77 = mau_0_io_pipe_phv_out_data_77; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_78 = mau_0_io_pipe_phv_out_data_78; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_79 = mau_0_io_pipe_phv_out_data_79; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_80 = mau_0_io_pipe_phv_out_data_80; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_81 = mau_0_io_pipe_phv_out_data_81; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_82 = mau_0_io_pipe_phv_out_data_82; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_83 = mau_0_io_pipe_phv_out_data_83; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_84 = mau_0_io_pipe_phv_out_data_84; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_85 = mau_0_io_pipe_phv_out_data_85; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_86 = mau_0_io_pipe_phv_out_data_86; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_87 = mau_0_io_pipe_phv_out_data_87; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_88 = mau_0_io_pipe_phv_out_data_88; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_89 = mau_0_io_pipe_phv_out_data_89; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_90 = mau_0_io_pipe_phv_out_data_90; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_91 = mau_0_io_pipe_phv_out_data_91; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_92 = mau_0_io_pipe_phv_out_data_92; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_93 = mau_0_io_pipe_phv_out_data_93; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_94 = mau_0_io_pipe_phv_out_data_94; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_95 = mau_0_io_pipe_phv_out_data_95; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_96 = mau_0_io_pipe_phv_out_data_96; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_97 = mau_0_io_pipe_phv_out_data_97; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_98 = mau_0_io_pipe_phv_out_data_98; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_99 = mau_0_io_pipe_phv_out_data_99; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_100 = mau_0_io_pipe_phv_out_data_100; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_101 = mau_0_io_pipe_phv_out_data_101; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_102 = mau_0_io_pipe_phv_out_data_102; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_103 = mau_0_io_pipe_phv_out_data_103; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_104 = mau_0_io_pipe_phv_out_data_104; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_105 = mau_0_io_pipe_phv_out_data_105; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_106 = mau_0_io_pipe_phv_out_data_106; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_107 = mau_0_io_pipe_phv_out_data_107; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_108 = mau_0_io_pipe_phv_out_data_108; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_109 = mau_0_io_pipe_phv_out_data_109; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_110 = mau_0_io_pipe_phv_out_data_110; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_111 = mau_0_io_pipe_phv_out_data_111; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_112 = mau_0_io_pipe_phv_out_data_112; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_113 = mau_0_io_pipe_phv_out_data_113; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_114 = mau_0_io_pipe_phv_out_data_114; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_115 = mau_0_io_pipe_phv_out_data_115; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_116 = mau_0_io_pipe_phv_out_data_116; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_117 = mau_0_io_pipe_phv_out_data_117; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_118 = mau_0_io_pipe_phv_out_data_118; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_119 = mau_0_io_pipe_phv_out_data_119; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_120 = mau_0_io_pipe_phv_out_data_120; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_121 = mau_0_io_pipe_phv_out_data_121; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_122 = mau_0_io_pipe_phv_out_data_122; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_123 = mau_0_io_pipe_phv_out_data_123; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_124 = mau_0_io_pipe_phv_out_data_124; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_125 = mau_0_io_pipe_phv_out_data_125; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_126 = mau_0_io_pipe_phv_out_data_126; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_127 = mau_0_io_pipe_phv_out_data_127; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_128 = mau_0_io_pipe_phv_out_data_128; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_129 = mau_0_io_pipe_phv_out_data_129; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_130 = mau_0_io_pipe_phv_out_data_130; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_131 = mau_0_io_pipe_phv_out_data_131; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_132 = mau_0_io_pipe_phv_out_data_132; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_133 = mau_0_io_pipe_phv_out_data_133; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_134 = mau_0_io_pipe_phv_out_data_134; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_135 = mau_0_io_pipe_phv_out_data_135; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_136 = mau_0_io_pipe_phv_out_data_136; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_137 = mau_0_io_pipe_phv_out_data_137; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_138 = mau_0_io_pipe_phv_out_data_138; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_139 = mau_0_io_pipe_phv_out_data_139; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_140 = mau_0_io_pipe_phv_out_data_140; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_141 = mau_0_io_pipe_phv_out_data_141; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_142 = mau_0_io_pipe_phv_out_data_142; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_143 = mau_0_io_pipe_phv_out_data_143; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_144 = mau_0_io_pipe_phv_out_data_144; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_145 = mau_0_io_pipe_phv_out_data_145; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_146 = mau_0_io_pipe_phv_out_data_146; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_147 = mau_0_io_pipe_phv_out_data_147; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_148 = mau_0_io_pipe_phv_out_data_148; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_149 = mau_0_io_pipe_phv_out_data_149; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_150 = mau_0_io_pipe_phv_out_data_150; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_151 = mau_0_io_pipe_phv_out_data_151; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_152 = mau_0_io_pipe_phv_out_data_152; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_153 = mau_0_io_pipe_phv_out_data_153; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_154 = mau_0_io_pipe_phv_out_data_154; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_155 = mau_0_io_pipe_phv_out_data_155; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_156 = mau_0_io_pipe_phv_out_data_156; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_157 = mau_0_io_pipe_phv_out_data_157; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_158 = mau_0_io_pipe_phv_out_data_158; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_159 = mau_0_io_pipe_phv_out_data_159; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_0 = mau_0_io_pipe_phv_out_header_0; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_1 = mau_0_io_pipe_phv_out_header_1; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_2 = mau_0_io_pipe_phv_out_header_2; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_3 = mau_0_io_pipe_phv_out_header_3; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_4 = mau_0_io_pipe_phv_out_header_4; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_5 = mau_0_io_pipe_phv_out_header_5; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_6 = mau_0_io_pipe_phv_out_header_6; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_7 = mau_0_io_pipe_phv_out_header_7; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_8 = mau_0_io_pipe_phv_out_header_8; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_9 = mau_0_io_pipe_phv_out_header_9; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_10 = mau_0_io_pipe_phv_out_header_10; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_11 = mau_0_io_pipe_phv_out_header_11; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_12 = mau_0_io_pipe_phv_out_header_12; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_13 = mau_0_io_pipe_phv_out_header_13; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_14 = mau_0_io_pipe_phv_out_header_14; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_15 = mau_0_io_pipe_phv_out_header_15; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_parse_current_state = mau_0_io_pipe_phv_out_parse_current_state; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_parse_current_offset = mau_0_io_pipe_phv_out_parse_current_offset; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_parse_transition_field = mau_0_io_pipe_phv_out_parse_transition_field; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_next_config_id = mau_0_io_pipe_phv_out_next_config_id; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_is_valid_processor = mau_0_io_pipe_phv_out_is_valid_processor; // @[parser.scala 32:35]
  assign mau_2_clock = clock;
  assign mau_2_io_pipe_phv_in_data_0 = mau_1_io_pipe_phv_out_data_0; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_1 = mau_1_io_pipe_phv_out_data_1; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_2 = mau_1_io_pipe_phv_out_data_2; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_3 = mau_1_io_pipe_phv_out_data_3; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_4 = mau_1_io_pipe_phv_out_data_4; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_5 = mau_1_io_pipe_phv_out_data_5; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_6 = mau_1_io_pipe_phv_out_data_6; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_7 = mau_1_io_pipe_phv_out_data_7; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_8 = mau_1_io_pipe_phv_out_data_8; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_9 = mau_1_io_pipe_phv_out_data_9; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_10 = mau_1_io_pipe_phv_out_data_10; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_11 = mau_1_io_pipe_phv_out_data_11; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_12 = mau_1_io_pipe_phv_out_data_12; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_13 = mau_1_io_pipe_phv_out_data_13; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_14 = mau_1_io_pipe_phv_out_data_14; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_15 = mau_1_io_pipe_phv_out_data_15; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_16 = mau_1_io_pipe_phv_out_data_16; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_17 = mau_1_io_pipe_phv_out_data_17; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_18 = mau_1_io_pipe_phv_out_data_18; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_19 = mau_1_io_pipe_phv_out_data_19; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_20 = mau_1_io_pipe_phv_out_data_20; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_21 = mau_1_io_pipe_phv_out_data_21; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_22 = mau_1_io_pipe_phv_out_data_22; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_23 = mau_1_io_pipe_phv_out_data_23; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_24 = mau_1_io_pipe_phv_out_data_24; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_25 = mau_1_io_pipe_phv_out_data_25; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_26 = mau_1_io_pipe_phv_out_data_26; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_27 = mau_1_io_pipe_phv_out_data_27; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_28 = mau_1_io_pipe_phv_out_data_28; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_29 = mau_1_io_pipe_phv_out_data_29; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_30 = mau_1_io_pipe_phv_out_data_30; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_31 = mau_1_io_pipe_phv_out_data_31; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_32 = mau_1_io_pipe_phv_out_data_32; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_33 = mau_1_io_pipe_phv_out_data_33; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_34 = mau_1_io_pipe_phv_out_data_34; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_35 = mau_1_io_pipe_phv_out_data_35; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_36 = mau_1_io_pipe_phv_out_data_36; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_37 = mau_1_io_pipe_phv_out_data_37; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_38 = mau_1_io_pipe_phv_out_data_38; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_39 = mau_1_io_pipe_phv_out_data_39; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_40 = mau_1_io_pipe_phv_out_data_40; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_41 = mau_1_io_pipe_phv_out_data_41; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_42 = mau_1_io_pipe_phv_out_data_42; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_43 = mau_1_io_pipe_phv_out_data_43; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_44 = mau_1_io_pipe_phv_out_data_44; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_45 = mau_1_io_pipe_phv_out_data_45; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_46 = mau_1_io_pipe_phv_out_data_46; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_47 = mau_1_io_pipe_phv_out_data_47; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_48 = mau_1_io_pipe_phv_out_data_48; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_49 = mau_1_io_pipe_phv_out_data_49; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_50 = mau_1_io_pipe_phv_out_data_50; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_51 = mau_1_io_pipe_phv_out_data_51; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_52 = mau_1_io_pipe_phv_out_data_52; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_53 = mau_1_io_pipe_phv_out_data_53; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_54 = mau_1_io_pipe_phv_out_data_54; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_55 = mau_1_io_pipe_phv_out_data_55; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_56 = mau_1_io_pipe_phv_out_data_56; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_57 = mau_1_io_pipe_phv_out_data_57; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_58 = mau_1_io_pipe_phv_out_data_58; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_59 = mau_1_io_pipe_phv_out_data_59; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_60 = mau_1_io_pipe_phv_out_data_60; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_61 = mau_1_io_pipe_phv_out_data_61; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_62 = mau_1_io_pipe_phv_out_data_62; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_63 = mau_1_io_pipe_phv_out_data_63; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_64 = mau_1_io_pipe_phv_out_data_64; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_65 = mau_1_io_pipe_phv_out_data_65; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_66 = mau_1_io_pipe_phv_out_data_66; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_67 = mau_1_io_pipe_phv_out_data_67; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_68 = mau_1_io_pipe_phv_out_data_68; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_69 = mau_1_io_pipe_phv_out_data_69; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_70 = mau_1_io_pipe_phv_out_data_70; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_71 = mau_1_io_pipe_phv_out_data_71; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_72 = mau_1_io_pipe_phv_out_data_72; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_73 = mau_1_io_pipe_phv_out_data_73; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_74 = mau_1_io_pipe_phv_out_data_74; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_75 = mau_1_io_pipe_phv_out_data_75; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_76 = mau_1_io_pipe_phv_out_data_76; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_77 = mau_1_io_pipe_phv_out_data_77; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_78 = mau_1_io_pipe_phv_out_data_78; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_79 = mau_1_io_pipe_phv_out_data_79; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_80 = mau_1_io_pipe_phv_out_data_80; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_81 = mau_1_io_pipe_phv_out_data_81; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_82 = mau_1_io_pipe_phv_out_data_82; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_83 = mau_1_io_pipe_phv_out_data_83; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_84 = mau_1_io_pipe_phv_out_data_84; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_85 = mau_1_io_pipe_phv_out_data_85; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_86 = mau_1_io_pipe_phv_out_data_86; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_87 = mau_1_io_pipe_phv_out_data_87; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_88 = mau_1_io_pipe_phv_out_data_88; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_89 = mau_1_io_pipe_phv_out_data_89; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_90 = mau_1_io_pipe_phv_out_data_90; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_91 = mau_1_io_pipe_phv_out_data_91; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_92 = mau_1_io_pipe_phv_out_data_92; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_93 = mau_1_io_pipe_phv_out_data_93; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_94 = mau_1_io_pipe_phv_out_data_94; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_95 = mau_1_io_pipe_phv_out_data_95; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_96 = mau_1_io_pipe_phv_out_data_96; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_97 = mau_1_io_pipe_phv_out_data_97; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_98 = mau_1_io_pipe_phv_out_data_98; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_99 = mau_1_io_pipe_phv_out_data_99; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_100 = mau_1_io_pipe_phv_out_data_100; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_101 = mau_1_io_pipe_phv_out_data_101; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_102 = mau_1_io_pipe_phv_out_data_102; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_103 = mau_1_io_pipe_phv_out_data_103; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_104 = mau_1_io_pipe_phv_out_data_104; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_105 = mau_1_io_pipe_phv_out_data_105; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_106 = mau_1_io_pipe_phv_out_data_106; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_107 = mau_1_io_pipe_phv_out_data_107; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_108 = mau_1_io_pipe_phv_out_data_108; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_109 = mau_1_io_pipe_phv_out_data_109; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_110 = mau_1_io_pipe_phv_out_data_110; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_111 = mau_1_io_pipe_phv_out_data_111; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_112 = mau_1_io_pipe_phv_out_data_112; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_113 = mau_1_io_pipe_phv_out_data_113; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_114 = mau_1_io_pipe_phv_out_data_114; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_115 = mau_1_io_pipe_phv_out_data_115; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_116 = mau_1_io_pipe_phv_out_data_116; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_117 = mau_1_io_pipe_phv_out_data_117; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_118 = mau_1_io_pipe_phv_out_data_118; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_119 = mau_1_io_pipe_phv_out_data_119; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_120 = mau_1_io_pipe_phv_out_data_120; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_121 = mau_1_io_pipe_phv_out_data_121; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_122 = mau_1_io_pipe_phv_out_data_122; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_123 = mau_1_io_pipe_phv_out_data_123; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_124 = mau_1_io_pipe_phv_out_data_124; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_125 = mau_1_io_pipe_phv_out_data_125; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_126 = mau_1_io_pipe_phv_out_data_126; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_127 = mau_1_io_pipe_phv_out_data_127; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_128 = mau_1_io_pipe_phv_out_data_128; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_129 = mau_1_io_pipe_phv_out_data_129; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_130 = mau_1_io_pipe_phv_out_data_130; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_131 = mau_1_io_pipe_phv_out_data_131; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_132 = mau_1_io_pipe_phv_out_data_132; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_133 = mau_1_io_pipe_phv_out_data_133; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_134 = mau_1_io_pipe_phv_out_data_134; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_135 = mau_1_io_pipe_phv_out_data_135; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_136 = mau_1_io_pipe_phv_out_data_136; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_137 = mau_1_io_pipe_phv_out_data_137; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_138 = mau_1_io_pipe_phv_out_data_138; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_139 = mau_1_io_pipe_phv_out_data_139; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_140 = mau_1_io_pipe_phv_out_data_140; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_141 = mau_1_io_pipe_phv_out_data_141; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_142 = mau_1_io_pipe_phv_out_data_142; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_143 = mau_1_io_pipe_phv_out_data_143; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_144 = mau_1_io_pipe_phv_out_data_144; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_145 = mau_1_io_pipe_phv_out_data_145; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_146 = mau_1_io_pipe_phv_out_data_146; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_147 = mau_1_io_pipe_phv_out_data_147; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_148 = mau_1_io_pipe_phv_out_data_148; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_149 = mau_1_io_pipe_phv_out_data_149; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_150 = mau_1_io_pipe_phv_out_data_150; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_151 = mau_1_io_pipe_phv_out_data_151; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_152 = mau_1_io_pipe_phv_out_data_152; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_153 = mau_1_io_pipe_phv_out_data_153; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_154 = mau_1_io_pipe_phv_out_data_154; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_155 = mau_1_io_pipe_phv_out_data_155; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_156 = mau_1_io_pipe_phv_out_data_156; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_157 = mau_1_io_pipe_phv_out_data_157; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_158 = mau_1_io_pipe_phv_out_data_158; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_159 = mau_1_io_pipe_phv_out_data_159; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_0 = mau_1_io_pipe_phv_out_header_0; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_1 = mau_1_io_pipe_phv_out_header_1; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_2 = mau_1_io_pipe_phv_out_header_2; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_3 = mau_1_io_pipe_phv_out_header_3; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_4 = mau_1_io_pipe_phv_out_header_4; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_5 = mau_1_io_pipe_phv_out_header_5; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_6 = mau_1_io_pipe_phv_out_header_6; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_7 = mau_1_io_pipe_phv_out_header_7; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_8 = mau_1_io_pipe_phv_out_header_8; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_9 = mau_1_io_pipe_phv_out_header_9; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_10 = mau_1_io_pipe_phv_out_header_10; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_11 = mau_1_io_pipe_phv_out_header_11; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_12 = mau_1_io_pipe_phv_out_header_12; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_13 = mau_1_io_pipe_phv_out_header_13; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_14 = mau_1_io_pipe_phv_out_header_14; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_15 = mau_1_io_pipe_phv_out_header_15; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_parse_current_state = mau_1_io_pipe_phv_out_parse_current_state; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_parse_current_offset = mau_1_io_pipe_phv_out_parse_current_offset; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_parse_transition_field = mau_1_io_pipe_phv_out_parse_transition_field; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_next_config_id = mau_1_io_pipe_phv_out_next_config_id; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_is_valid_processor = mau_1_io_pipe_phv_out_is_valid_processor; // @[parser.scala 32:35]
  assign mau_3_clock = clock;
  assign mau_3_io_pipe_phv_in_data_0 = mau_2_io_pipe_phv_out_data_0; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_1 = mau_2_io_pipe_phv_out_data_1; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_2 = mau_2_io_pipe_phv_out_data_2; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_3 = mau_2_io_pipe_phv_out_data_3; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_4 = mau_2_io_pipe_phv_out_data_4; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_5 = mau_2_io_pipe_phv_out_data_5; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_6 = mau_2_io_pipe_phv_out_data_6; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_7 = mau_2_io_pipe_phv_out_data_7; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_8 = mau_2_io_pipe_phv_out_data_8; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_9 = mau_2_io_pipe_phv_out_data_9; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_10 = mau_2_io_pipe_phv_out_data_10; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_11 = mau_2_io_pipe_phv_out_data_11; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_12 = mau_2_io_pipe_phv_out_data_12; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_13 = mau_2_io_pipe_phv_out_data_13; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_14 = mau_2_io_pipe_phv_out_data_14; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_15 = mau_2_io_pipe_phv_out_data_15; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_16 = mau_2_io_pipe_phv_out_data_16; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_17 = mau_2_io_pipe_phv_out_data_17; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_18 = mau_2_io_pipe_phv_out_data_18; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_19 = mau_2_io_pipe_phv_out_data_19; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_20 = mau_2_io_pipe_phv_out_data_20; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_21 = mau_2_io_pipe_phv_out_data_21; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_22 = mau_2_io_pipe_phv_out_data_22; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_23 = mau_2_io_pipe_phv_out_data_23; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_24 = mau_2_io_pipe_phv_out_data_24; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_25 = mau_2_io_pipe_phv_out_data_25; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_26 = mau_2_io_pipe_phv_out_data_26; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_27 = mau_2_io_pipe_phv_out_data_27; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_28 = mau_2_io_pipe_phv_out_data_28; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_29 = mau_2_io_pipe_phv_out_data_29; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_30 = mau_2_io_pipe_phv_out_data_30; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_31 = mau_2_io_pipe_phv_out_data_31; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_32 = mau_2_io_pipe_phv_out_data_32; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_33 = mau_2_io_pipe_phv_out_data_33; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_34 = mau_2_io_pipe_phv_out_data_34; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_35 = mau_2_io_pipe_phv_out_data_35; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_36 = mau_2_io_pipe_phv_out_data_36; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_37 = mau_2_io_pipe_phv_out_data_37; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_38 = mau_2_io_pipe_phv_out_data_38; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_39 = mau_2_io_pipe_phv_out_data_39; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_40 = mau_2_io_pipe_phv_out_data_40; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_41 = mau_2_io_pipe_phv_out_data_41; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_42 = mau_2_io_pipe_phv_out_data_42; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_43 = mau_2_io_pipe_phv_out_data_43; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_44 = mau_2_io_pipe_phv_out_data_44; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_45 = mau_2_io_pipe_phv_out_data_45; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_46 = mau_2_io_pipe_phv_out_data_46; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_47 = mau_2_io_pipe_phv_out_data_47; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_48 = mau_2_io_pipe_phv_out_data_48; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_49 = mau_2_io_pipe_phv_out_data_49; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_50 = mau_2_io_pipe_phv_out_data_50; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_51 = mau_2_io_pipe_phv_out_data_51; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_52 = mau_2_io_pipe_phv_out_data_52; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_53 = mau_2_io_pipe_phv_out_data_53; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_54 = mau_2_io_pipe_phv_out_data_54; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_55 = mau_2_io_pipe_phv_out_data_55; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_56 = mau_2_io_pipe_phv_out_data_56; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_57 = mau_2_io_pipe_phv_out_data_57; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_58 = mau_2_io_pipe_phv_out_data_58; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_59 = mau_2_io_pipe_phv_out_data_59; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_60 = mau_2_io_pipe_phv_out_data_60; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_61 = mau_2_io_pipe_phv_out_data_61; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_62 = mau_2_io_pipe_phv_out_data_62; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_63 = mau_2_io_pipe_phv_out_data_63; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_64 = mau_2_io_pipe_phv_out_data_64; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_65 = mau_2_io_pipe_phv_out_data_65; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_66 = mau_2_io_pipe_phv_out_data_66; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_67 = mau_2_io_pipe_phv_out_data_67; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_68 = mau_2_io_pipe_phv_out_data_68; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_69 = mau_2_io_pipe_phv_out_data_69; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_70 = mau_2_io_pipe_phv_out_data_70; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_71 = mau_2_io_pipe_phv_out_data_71; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_72 = mau_2_io_pipe_phv_out_data_72; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_73 = mau_2_io_pipe_phv_out_data_73; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_74 = mau_2_io_pipe_phv_out_data_74; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_75 = mau_2_io_pipe_phv_out_data_75; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_76 = mau_2_io_pipe_phv_out_data_76; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_77 = mau_2_io_pipe_phv_out_data_77; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_78 = mau_2_io_pipe_phv_out_data_78; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_79 = mau_2_io_pipe_phv_out_data_79; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_80 = mau_2_io_pipe_phv_out_data_80; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_81 = mau_2_io_pipe_phv_out_data_81; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_82 = mau_2_io_pipe_phv_out_data_82; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_83 = mau_2_io_pipe_phv_out_data_83; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_84 = mau_2_io_pipe_phv_out_data_84; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_85 = mau_2_io_pipe_phv_out_data_85; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_86 = mau_2_io_pipe_phv_out_data_86; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_87 = mau_2_io_pipe_phv_out_data_87; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_88 = mau_2_io_pipe_phv_out_data_88; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_89 = mau_2_io_pipe_phv_out_data_89; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_90 = mau_2_io_pipe_phv_out_data_90; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_91 = mau_2_io_pipe_phv_out_data_91; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_92 = mau_2_io_pipe_phv_out_data_92; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_93 = mau_2_io_pipe_phv_out_data_93; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_94 = mau_2_io_pipe_phv_out_data_94; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_95 = mau_2_io_pipe_phv_out_data_95; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_96 = mau_2_io_pipe_phv_out_data_96; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_97 = mau_2_io_pipe_phv_out_data_97; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_98 = mau_2_io_pipe_phv_out_data_98; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_99 = mau_2_io_pipe_phv_out_data_99; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_100 = mau_2_io_pipe_phv_out_data_100; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_101 = mau_2_io_pipe_phv_out_data_101; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_102 = mau_2_io_pipe_phv_out_data_102; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_103 = mau_2_io_pipe_phv_out_data_103; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_104 = mau_2_io_pipe_phv_out_data_104; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_105 = mau_2_io_pipe_phv_out_data_105; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_106 = mau_2_io_pipe_phv_out_data_106; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_107 = mau_2_io_pipe_phv_out_data_107; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_108 = mau_2_io_pipe_phv_out_data_108; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_109 = mau_2_io_pipe_phv_out_data_109; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_110 = mau_2_io_pipe_phv_out_data_110; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_111 = mau_2_io_pipe_phv_out_data_111; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_112 = mau_2_io_pipe_phv_out_data_112; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_113 = mau_2_io_pipe_phv_out_data_113; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_114 = mau_2_io_pipe_phv_out_data_114; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_115 = mau_2_io_pipe_phv_out_data_115; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_116 = mau_2_io_pipe_phv_out_data_116; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_117 = mau_2_io_pipe_phv_out_data_117; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_118 = mau_2_io_pipe_phv_out_data_118; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_119 = mau_2_io_pipe_phv_out_data_119; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_120 = mau_2_io_pipe_phv_out_data_120; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_121 = mau_2_io_pipe_phv_out_data_121; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_122 = mau_2_io_pipe_phv_out_data_122; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_123 = mau_2_io_pipe_phv_out_data_123; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_124 = mau_2_io_pipe_phv_out_data_124; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_125 = mau_2_io_pipe_phv_out_data_125; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_126 = mau_2_io_pipe_phv_out_data_126; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_127 = mau_2_io_pipe_phv_out_data_127; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_128 = mau_2_io_pipe_phv_out_data_128; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_129 = mau_2_io_pipe_phv_out_data_129; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_130 = mau_2_io_pipe_phv_out_data_130; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_131 = mau_2_io_pipe_phv_out_data_131; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_132 = mau_2_io_pipe_phv_out_data_132; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_133 = mau_2_io_pipe_phv_out_data_133; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_134 = mau_2_io_pipe_phv_out_data_134; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_135 = mau_2_io_pipe_phv_out_data_135; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_136 = mau_2_io_pipe_phv_out_data_136; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_137 = mau_2_io_pipe_phv_out_data_137; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_138 = mau_2_io_pipe_phv_out_data_138; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_139 = mau_2_io_pipe_phv_out_data_139; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_140 = mau_2_io_pipe_phv_out_data_140; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_141 = mau_2_io_pipe_phv_out_data_141; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_142 = mau_2_io_pipe_phv_out_data_142; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_143 = mau_2_io_pipe_phv_out_data_143; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_144 = mau_2_io_pipe_phv_out_data_144; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_145 = mau_2_io_pipe_phv_out_data_145; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_146 = mau_2_io_pipe_phv_out_data_146; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_147 = mau_2_io_pipe_phv_out_data_147; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_148 = mau_2_io_pipe_phv_out_data_148; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_149 = mau_2_io_pipe_phv_out_data_149; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_150 = mau_2_io_pipe_phv_out_data_150; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_151 = mau_2_io_pipe_phv_out_data_151; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_152 = mau_2_io_pipe_phv_out_data_152; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_153 = mau_2_io_pipe_phv_out_data_153; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_154 = mau_2_io_pipe_phv_out_data_154; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_155 = mau_2_io_pipe_phv_out_data_155; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_156 = mau_2_io_pipe_phv_out_data_156; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_157 = mau_2_io_pipe_phv_out_data_157; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_158 = mau_2_io_pipe_phv_out_data_158; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_159 = mau_2_io_pipe_phv_out_data_159; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_0 = mau_2_io_pipe_phv_out_header_0; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_1 = mau_2_io_pipe_phv_out_header_1; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_2 = mau_2_io_pipe_phv_out_header_2; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_3 = mau_2_io_pipe_phv_out_header_3; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_4 = mau_2_io_pipe_phv_out_header_4; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_5 = mau_2_io_pipe_phv_out_header_5; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_6 = mau_2_io_pipe_phv_out_header_6; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_7 = mau_2_io_pipe_phv_out_header_7; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_8 = mau_2_io_pipe_phv_out_header_8; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_9 = mau_2_io_pipe_phv_out_header_9; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_10 = mau_2_io_pipe_phv_out_header_10; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_11 = mau_2_io_pipe_phv_out_header_11; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_12 = mau_2_io_pipe_phv_out_header_12; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_13 = mau_2_io_pipe_phv_out_header_13; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_14 = mau_2_io_pipe_phv_out_header_14; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_15 = mau_2_io_pipe_phv_out_header_15; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_parse_current_state = mau_2_io_pipe_phv_out_parse_current_state; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_parse_current_offset = mau_2_io_pipe_phv_out_parse_current_offset; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_parse_transition_field = mau_2_io_pipe_phv_out_parse_transition_field; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_next_config_id = mau_2_io_pipe_phv_out_next_config_id; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_is_valid_processor = mau_2_io_pipe_phv_out_is_valid_processor; // @[parser.scala 32:35]
endmodule
