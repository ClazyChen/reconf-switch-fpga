module PrimitiveGetSourcePISA(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  input  [7:0]  io_args_in_0,
  input  [7:0]  io_args_in_1,
  input  [7:0]  io_args_in_2,
  input  [7:0]  io_args_in_3,
  input  [7:0]  io_args_in_4,
  input  [7:0]  io_args_in_5,
  input  [7:0]  io_args_in_6,
  input  [17:0] io_vliw_in_0,
  input  [17:0] io_vliw_in_1,
  input  [17:0] io_vliw_in_2,
  input  [17:0] io_vliw_in_3,
  input  [17:0] io_vliw_in_4,
  input  [17:0] io_vliw_in_5,
  input  [17:0] io_vliw_in_6,
  input  [17:0] io_vliw_in_7,
  input  [17:0] io_vliw_in_8,
  input  [17:0] io_vliw_in_9,
  input  [17:0] io_vliw_in_10,
  input  [17:0] io_vliw_in_11,
  input  [17:0] io_vliw_in_12,
  input  [17:0] io_vliw_in_13,
  input  [17:0] io_vliw_in_14,
  input  [17:0] io_vliw_in_15,
  input  [17:0] io_vliw_in_16,
  input  [17:0] io_vliw_in_17,
  input  [17:0] io_vliw_in_18,
  input  [17:0] io_vliw_in_19,
  input  [17:0] io_vliw_in_20,
  input  [17:0] io_vliw_in_21,
  input  [17:0] io_vliw_in_22,
  input  [17:0] io_vliw_in_23,
  input  [17:0] io_vliw_in_24,
  input  [17:0] io_vliw_in_25,
  input  [17:0] io_vliw_in_26,
  input  [17:0] io_vliw_in_27,
  input  [17:0] io_vliw_in_28,
  input  [17:0] io_vliw_in_29,
  input  [17:0] io_vliw_in_30,
  input  [17:0] io_vliw_in_31,
  input  [17:0] io_vliw_in_32,
  input  [17:0] io_vliw_in_33,
  input  [17:0] io_vliw_in_34,
  input  [17:0] io_vliw_in_35,
  input  [17:0] io_vliw_in_36,
  input  [17:0] io_vliw_in_37,
  input  [17:0] io_vliw_in_38,
  input  [17:0] io_vliw_in_39,
  input  [17:0] io_vliw_in_40,
  input  [17:0] io_vliw_in_41,
  input  [17:0] io_vliw_in_42,
  input  [17:0] io_vliw_in_43,
  input  [17:0] io_vliw_in_44,
  input  [17:0] io_vliw_in_45,
  input  [17:0] io_vliw_in_46,
  input  [17:0] io_vliw_in_47,
  input  [17:0] io_vliw_in_48,
  input  [17:0] io_vliw_in_49,
  input  [17:0] io_vliw_in_50,
  input  [17:0] io_vliw_in_51,
  input  [17:0] io_vliw_in_52,
  input  [17:0] io_vliw_in_53,
  input  [17:0] io_vliw_in_54,
  input  [17:0] io_vliw_in_55,
  input  [17:0] io_vliw_in_56,
  input  [17:0] io_vliw_in_57,
  input  [17:0] io_vliw_in_58,
  input  [17:0] io_vliw_in_59,
  input  [17:0] io_vliw_in_60,
  input  [17:0] io_vliw_in_61,
  input  [17:0] io_vliw_in_62,
  input  [17:0] io_vliw_in_63,
  input  [17:0] io_vliw_in_64,
  input  [17:0] io_vliw_in_65,
  input  [17:0] io_vliw_in_66,
  input  [17:0] io_vliw_in_67,
  input  [17:0] io_vliw_in_68,
  input  [17:0] io_vliw_in_69,
  input  [14:0] io_nid_in,
  output [14:0] io_nid_out,
  output [1:0]  io_tag_out_0,
  output [1:0]  io_tag_out_1,
  output [1:0]  io_tag_out_2,
  output [1:0]  io_tag_out_3,
  output [1:0]  io_tag_out_4,
  output [1:0]  io_tag_out_5,
  output [1:0]  io_tag_out_6,
  output [1:0]  io_tag_out_7,
  output [1:0]  io_tag_out_8,
  output [1:0]  io_tag_out_9,
  output [1:0]  io_tag_out_10,
  output [1:0]  io_tag_out_11,
  output [1:0]  io_tag_out_12,
  output [1:0]  io_tag_out_13,
  output [1:0]  io_tag_out_14,
  output [1:0]  io_tag_out_15,
  output [1:0]  io_tag_out_16,
  output [1:0]  io_tag_out_17,
  output [1:0]  io_tag_out_18,
  output [1:0]  io_tag_out_19,
  output [1:0]  io_tag_out_20,
  output [1:0]  io_tag_out_21,
  output [1:0]  io_tag_out_22,
  output [1:0]  io_tag_out_23,
  output [1:0]  io_tag_out_24,
  output [1:0]  io_tag_out_25,
  output [1:0]  io_tag_out_26,
  output [1:0]  io_tag_out_27,
  output [1:0]  io_tag_out_28,
  output [1:0]  io_tag_out_29,
  output [1:0]  io_tag_out_30,
  output [1:0]  io_tag_out_31,
  output [1:0]  io_tag_out_32,
  output [1:0]  io_tag_out_33,
  output [1:0]  io_tag_out_34,
  output [1:0]  io_tag_out_35,
  output [1:0]  io_tag_out_36,
  output [1:0]  io_tag_out_37,
  output [1:0]  io_tag_out_38,
  output [1:0]  io_tag_out_39,
  output [1:0]  io_tag_out_40,
  output [1:0]  io_tag_out_41,
  output [1:0]  io_tag_out_42,
  output [1:0]  io_tag_out_43,
  output [1:0]  io_tag_out_44,
  output [1:0]  io_tag_out_45,
  output [1:0]  io_tag_out_46,
  output [1:0]  io_tag_out_47,
  output [1:0]  io_tag_out_48,
  output [1:0]  io_tag_out_49,
  output [1:0]  io_tag_out_50,
  output [1:0]  io_tag_out_51,
  output [1:0]  io_tag_out_52,
  output [1:0]  io_tag_out_53,
  output [1:0]  io_tag_out_54,
  output [1:0]  io_tag_out_55,
  output [1:0]  io_tag_out_56,
  output [1:0]  io_tag_out_57,
  output [1:0]  io_tag_out_58,
  output [1:0]  io_tag_out_59,
  output [1:0]  io_tag_out_60,
  output [1:0]  io_tag_out_61,
  output [1:0]  io_tag_out_62,
  output [1:0]  io_tag_out_63,
  output [1:0]  io_tag_out_64,
  output [1:0]  io_tag_out_65,
  output [1:0]  io_tag_out_66,
  output [1:0]  io_tag_out_67,
  output [1:0]  io_tag_out_68,
  output [1:0]  io_tag_out_69,
  output [7:0]  io_field_set_field8_0,
  output [7:0]  io_field_set_field8_1,
  output [7:0]  io_field_set_field8_2,
  output [7:0]  io_field_set_field8_3,
  output [7:0]  io_field_set_field8_4,
  output [7:0]  io_field_set_field8_5,
  output [7:0]  io_field_set_field8_6,
  output [7:0]  io_field_set_field8_7,
  output [7:0]  io_field_set_field8_8,
  output [7:0]  io_field_set_field8_9,
  output [7:0]  io_field_set_field8_10,
  output [7:0]  io_field_set_field8_11,
  output [7:0]  io_field_set_field8_12,
  output [7:0]  io_field_set_field8_13,
  output [7:0]  io_field_set_field8_14,
  output [7:0]  io_field_set_field8_15,
  output [7:0]  io_field_set_field8_16,
  output [7:0]  io_field_set_field8_17,
  output [7:0]  io_field_set_field8_18,
  output [7:0]  io_field_set_field8_19,
  output [7:0]  io_field_set_field8_20,
  output [7:0]  io_field_set_field8_21,
  output [7:0]  io_field_set_field8_22,
  output [7:0]  io_field_set_field8_23,
  output [7:0]  io_field_set_field8_24,
  output [7:0]  io_field_set_field8_25,
  output [7:0]  io_field_set_field8_26,
  output [7:0]  io_field_set_field8_27,
  output [7:0]  io_field_set_field8_28,
  output [7:0]  io_field_set_field8_29,
  output [7:0]  io_field_set_field8_30,
  output [7:0]  io_field_set_field8_31,
  output [15:0] io_field_set_field16_0,
  output [15:0] io_field_set_field16_1,
  output [15:0] io_field_set_field16_2,
  output [15:0] io_field_set_field16_3,
  output [15:0] io_field_set_field16_4,
  output [15:0] io_field_set_field16_5,
  output [15:0] io_field_set_field16_6,
  output [15:0] io_field_set_field16_7,
  output [15:0] io_field_set_field16_8,
  output [15:0] io_field_set_field16_9,
  output [15:0] io_field_set_field16_10,
  output [15:0] io_field_set_field16_11,
  output [15:0] io_field_set_field16_12,
  output [15:0] io_field_set_field16_13,
  output [15:0] io_field_set_field16_14,
  output [15:0] io_field_set_field16_15,
  output [15:0] io_field_set_field16_16,
  output [15:0] io_field_set_field16_17,
  output [15:0] io_field_set_field16_18,
  output [15:0] io_field_set_field16_19,
  output [15:0] io_field_set_field16_20,
  output [15:0] io_field_set_field16_21,
  output [15:0] io_field_set_field16_22,
  output [15:0] io_field_set_field16_23,
  output [15:0] io_field_set_field16_24,
  output [15:0] io_field_set_field16_25,
  output [15:0] io_field_set_field16_26,
  output [15:0] io_field_set_field16_27,
  output [15:0] io_field_set_field16_28,
  output [15:0] io_field_set_field16_29,
  output [15:0] io_field_set_field16_30,
  output [15:0] io_field_set_field16_31,
  output [15:0] io_field_set_field16_32,
  output [15:0] io_field_set_field16_33,
  output [15:0] io_field_set_field16_34,
  output [15:0] io_field_set_field16_35,
  output [15:0] io_field_set_field16_36,
  output [15:0] io_field_set_field16_37
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_1; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_2; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_3; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_4; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_5; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_6; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_7; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_8; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_9; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_10; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_11; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_12; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_13; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_14; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_15; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_16; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_17; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_18; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_19; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_20; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_21; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_22; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_23; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_24; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_25; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_26; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_27; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_28; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_29; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_30; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_31; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_32; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_33; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_34; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_35; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_36; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_37; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_38; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_39; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_40; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_41; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_42; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_43; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_44; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_45; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_46; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_47; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_48; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_49; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_50; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_51; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_52; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_53; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_54; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_55; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_56; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_57; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_58; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_59; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_60; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_61; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_62; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_63; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_64; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_65; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_66; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_67; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_68; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_69; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_70; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_71; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_72; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_73; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_74; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_75; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_76; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_77; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_78; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_79; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_80; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_81; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_82; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_83; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_84; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_85; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_86; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_87; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_88; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_89; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_90; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_91; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_92; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_93; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_94; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_95; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_96; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_97; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_98; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_99; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_100; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_101; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_102; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_103; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_104; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_105; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_106; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_107; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_108; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_109; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_110; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_111; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_112; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_113; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_114; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_115; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_116; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_117; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_118; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_119; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_120; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_121; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_122; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_123; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_124; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_125; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_126; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_127; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_128; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_129; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_130; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_131; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_132; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_133; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_134; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_135; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_136; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_137; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_138; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_139; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_140; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_141; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_142; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_143; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_144; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_145; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_146; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_147; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_148; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_149; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_150; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_151; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_152; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_153; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_154; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_155; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_156; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_157; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_158; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_159; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_160; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_161; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_162; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_163; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_164; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_165; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_166; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_167; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_168; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_169; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_170; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_171; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_172; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_173; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_174; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_175; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_176; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_177; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_178; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_179; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_180; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_181; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_182; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_183; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_184; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_185; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_186; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_187; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_188; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_189; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_190; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_191; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_192; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_193; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_194; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_195; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_196; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_197; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_198; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_199; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_200; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_201; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_202; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_203; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_204; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_205; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_206; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_207; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_208; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_209; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_210; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_211; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_212; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_213; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_214; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_215; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_216; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_217; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_218; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_219; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_220; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_221; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_222; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_223; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_224; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_225; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_226; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_227; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_228; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_229; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_230; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_231; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_232; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_233; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_234; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_235; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_236; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_237; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_238; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_239; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_240; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_241; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_242; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_243; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_244; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_245; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_246; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_247; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_248; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_249; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_250; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_251; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_252; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_253; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_254; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_255; // @[executor_pisa.scala 161:22]
  reg [3:0] phv_next_processor_id; // @[executor_pisa.scala 161:22]
  reg  phv_next_config_id; // @[executor_pisa.scala 161:22]
  reg [7:0] args_0; // @[executor_pisa.scala 165:23]
  reg [7:0] args_1; // @[executor_pisa.scala 165:23]
  reg [7:0] args_2; // @[executor_pisa.scala 165:23]
  reg [7:0] args_3; // @[executor_pisa.scala 165:23]
  reg [7:0] args_4; // @[executor_pisa.scala 165:23]
  reg [7:0] args_5; // @[executor_pisa.scala 165:23]
  reg [7:0] args_6; // @[executor_pisa.scala 165:23]
  reg [17:0] vliw_0; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_1; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_2; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_3; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_4; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_5; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_6; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_7; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_8; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_9; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_10; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_11; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_12; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_13; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_14; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_15; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_16; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_17; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_18; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_19; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_20; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_21; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_22; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_23; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_24; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_25; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_26; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_27; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_28; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_29; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_30; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_31; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_32; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_33; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_34; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_35; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_36; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_37; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_38; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_39; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_40; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_41; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_42; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_43; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_44; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_45; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_46; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_47; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_48; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_49; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_50; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_51; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_52; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_53; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_54; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_55; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_56; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_57; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_58; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_59; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_60; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_61; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_62; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_63; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_64; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_65; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_66; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_67; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_68; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_69; // @[executor_pisa.scala 168:23]
  reg [14:0] nid; // @[executor_pisa.scala 171:23]
  wire [3:0] opcode = vliw_0[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2 = vliw_0[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset = parameter_2[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length = parameter_2[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T = {{1'd0}, args_offset}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset = _total_offset_T[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1 = 3'h1 == total_offset ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2 = 3'h2 == total_offset ? args_2 : _GEN_1; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3 = 3'h3 == total_offset ? args_3 : _GEN_2; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4 = 3'h4 == total_offset ? args_4 : _GEN_3; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5 = 3'h5 == total_offset ? args_5 : _GEN_4; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_6 = 3'h6 == total_offset ? args_6 : _GEN_5; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_7 = total_offset < 3'h7 ? _GEN_6 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_0 = 3'h0 < args_length ? _GEN_7 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_9 = opcode == 4'ha ? field_bytes_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_10 = opcode == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3 = opcode == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_1 = _T_3 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_11 = opcode == 4'h8 | opcode == 4'hb ? parameter_2[7:0] : _GEN_9; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_12 = opcode == 4'h8 | opcode == 4'hb ? _field_tag_T_1 : _GEN_10; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_13 = 14'h0 == parameter_2 ? phv_data_0 : _GEN_11; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_14 = 14'h1 == parameter_2 ? phv_data_1 : _GEN_13; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_15 = 14'h2 == parameter_2 ? phv_data_2 : _GEN_14; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_16 = 14'h3 == parameter_2 ? phv_data_3 : _GEN_15; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_17 = 14'h4 == parameter_2 ? phv_data_4 : _GEN_16; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_18 = 14'h5 == parameter_2 ? phv_data_5 : _GEN_17; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_19 = 14'h6 == parameter_2 ? phv_data_6 : _GEN_18; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_20 = 14'h7 == parameter_2 ? phv_data_7 : _GEN_19; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_21 = 14'h8 == parameter_2 ? phv_data_8 : _GEN_20; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_22 = 14'h9 == parameter_2 ? phv_data_9 : _GEN_21; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_23 = 14'ha == parameter_2 ? phv_data_10 : _GEN_22; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_24 = 14'hb == parameter_2 ? phv_data_11 : _GEN_23; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_25 = 14'hc == parameter_2 ? phv_data_12 : _GEN_24; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_26 = 14'hd == parameter_2 ? phv_data_13 : _GEN_25; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_27 = 14'he == parameter_2 ? phv_data_14 : _GEN_26; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_28 = 14'hf == parameter_2 ? phv_data_15 : _GEN_27; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_29 = 14'h10 == parameter_2 ? phv_data_16 : _GEN_28; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_30 = 14'h11 == parameter_2 ? phv_data_17 : _GEN_29; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_31 = 14'h12 == parameter_2 ? phv_data_18 : _GEN_30; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_32 = 14'h13 == parameter_2 ? phv_data_19 : _GEN_31; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_33 = 14'h14 == parameter_2 ? phv_data_20 : _GEN_32; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_34 = 14'h15 == parameter_2 ? phv_data_21 : _GEN_33; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_35 = 14'h16 == parameter_2 ? phv_data_22 : _GEN_34; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_36 = 14'h17 == parameter_2 ? phv_data_23 : _GEN_35; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_37 = 14'h18 == parameter_2 ? phv_data_24 : _GEN_36; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_38 = 14'h19 == parameter_2 ? phv_data_25 : _GEN_37; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_39 = 14'h1a == parameter_2 ? phv_data_26 : _GEN_38; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_40 = 14'h1b == parameter_2 ? phv_data_27 : _GEN_39; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_41 = 14'h1c == parameter_2 ? phv_data_28 : _GEN_40; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_42 = 14'h1d == parameter_2 ? phv_data_29 : _GEN_41; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_43 = 14'h1e == parameter_2 ? phv_data_30 : _GEN_42; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_44 = 14'h1f == parameter_2 ? phv_data_31 : _GEN_43; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_1 = vliw_1[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_1 = vliw_1[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_1 = parameter_2_1[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_1 = parameter_2_1[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_1 = {{1'd0}, args_offset_1}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_1 = _total_offset_T_1[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_48 = 3'h1 == total_offset_1 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_49 = 3'h2 == total_offset_1 ? args_2 : _GEN_48; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_50 = 3'h3 == total_offset_1 ? args_3 : _GEN_49; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_51 = 3'h4 == total_offset_1 ? args_4 : _GEN_50; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_52 = 3'h5 == total_offset_1 ? args_5 : _GEN_51; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_53 = 3'h6 == total_offset_1 ? args_6 : _GEN_52; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_54 = total_offset_1 < 3'h7 ? _GEN_53 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_1_0 = 3'h0 < args_length_1 ? _GEN_54 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_56 = opcode_1 == 4'ha ? field_bytes_1_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_57 = opcode_1 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_42 = opcode_1 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_3 = _T_42 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_58 = opcode_1 == 4'h8 | opcode_1 == 4'hb ? parameter_2_1[7:0] : _GEN_56; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_59 = opcode_1 == 4'h8 | opcode_1 == 4'hb ? _field_tag_T_3 : _GEN_57; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_60 = 14'h0 == parameter_2_1 ? phv_data_0 : _GEN_58; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_61 = 14'h1 == parameter_2_1 ? phv_data_1 : _GEN_60; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_62 = 14'h2 == parameter_2_1 ? phv_data_2 : _GEN_61; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_63 = 14'h3 == parameter_2_1 ? phv_data_3 : _GEN_62; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_64 = 14'h4 == parameter_2_1 ? phv_data_4 : _GEN_63; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_65 = 14'h5 == parameter_2_1 ? phv_data_5 : _GEN_64; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_66 = 14'h6 == parameter_2_1 ? phv_data_6 : _GEN_65; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_67 = 14'h7 == parameter_2_1 ? phv_data_7 : _GEN_66; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_68 = 14'h8 == parameter_2_1 ? phv_data_8 : _GEN_67; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_69 = 14'h9 == parameter_2_1 ? phv_data_9 : _GEN_68; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_70 = 14'ha == parameter_2_1 ? phv_data_10 : _GEN_69; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_71 = 14'hb == parameter_2_1 ? phv_data_11 : _GEN_70; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_72 = 14'hc == parameter_2_1 ? phv_data_12 : _GEN_71; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_73 = 14'hd == parameter_2_1 ? phv_data_13 : _GEN_72; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_74 = 14'he == parameter_2_1 ? phv_data_14 : _GEN_73; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_75 = 14'hf == parameter_2_1 ? phv_data_15 : _GEN_74; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_76 = 14'h10 == parameter_2_1 ? phv_data_16 : _GEN_75; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_77 = 14'h11 == parameter_2_1 ? phv_data_17 : _GEN_76; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_78 = 14'h12 == parameter_2_1 ? phv_data_18 : _GEN_77; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_79 = 14'h13 == parameter_2_1 ? phv_data_19 : _GEN_78; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_80 = 14'h14 == parameter_2_1 ? phv_data_20 : _GEN_79; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_81 = 14'h15 == parameter_2_1 ? phv_data_21 : _GEN_80; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_82 = 14'h16 == parameter_2_1 ? phv_data_22 : _GEN_81; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_83 = 14'h17 == parameter_2_1 ? phv_data_23 : _GEN_82; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_84 = 14'h18 == parameter_2_1 ? phv_data_24 : _GEN_83; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_85 = 14'h19 == parameter_2_1 ? phv_data_25 : _GEN_84; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_86 = 14'h1a == parameter_2_1 ? phv_data_26 : _GEN_85; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_87 = 14'h1b == parameter_2_1 ? phv_data_27 : _GEN_86; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_88 = 14'h1c == parameter_2_1 ? phv_data_28 : _GEN_87; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_89 = 14'h1d == parameter_2_1 ? phv_data_29 : _GEN_88; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_90 = 14'h1e == parameter_2_1 ? phv_data_30 : _GEN_89; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_91 = 14'h1f == parameter_2_1 ? phv_data_31 : _GEN_90; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_2 = vliw_2[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_2 = vliw_2[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_2 = parameter_2_2[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_2 = parameter_2_2[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_2 = {{1'd0}, args_offset_2}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_2 = _total_offset_T_2[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_95 = 3'h1 == total_offset_2 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_96 = 3'h2 == total_offset_2 ? args_2 : _GEN_95; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_97 = 3'h3 == total_offset_2 ? args_3 : _GEN_96; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_98 = 3'h4 == total_offset_2 ? args_4 : _GEN_97; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_99 = 3'h5 == total_offset_2 ? args_5 : _GEN_98; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_100 = 3'h6 == total_offset_2 ? args_6 : _GEN_99; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_101 = total_offset_2 < 3'h7 ? _GEN_100 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_2_0 = 3'h0 < args_length_2 ? _GEN_101 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_103 = opcode_2 == 4'ha ? field_bytes_2_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_104 = opcode_2 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_81 = opcode_2 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_5 = _T_81 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_105 = opcode_2 == 4'h8 | opcode_2 == 4'hb ? parameter_2_2[7:0] : _GEN_103; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_106 = opcode_2 == 4'h8 | opcode_2 == 4'hb ? _field_tag_T_5 : _GEN_104; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_107 = 14'h0 == parameter_2_2 ? phv_data_0 : _GEN_105; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_108 = 14'h1 == parameter_2_2 ? phv_data_1 : _GEN_107; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_109 = 14'h2 == parameter_2_2 ? phv_data_2 : _GEN_108; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_110 = 14'h3 == parameter_2_2 ? phv_data_3 : _GEN_109; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_111 = 14'h4 == parameter_2_2 ? phv_data_4 : _GEN_110; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_112 = 14'h5 == parameter_2_2 ? phv_data_5 : _GEN_111; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_113 = 14'h6 == parameter_2_2 ? phv_data_6 : _GEN_112; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_114 = 14'h7 == parameter_2_2 ? phv_data_7 : _GEN_113; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_115 = 14'h8 == parameter_2_2 ? phv_data_8 : _GEN_114; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_116 = 14'h9 == parameter_2_2 ? phv_data_9 : _GEN_115; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_117 = 14'ha == parameter_2_2 ? phv_data_10 : _GEN_116; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_118 = 14'hb == parameter_2_2 ? phv_data_11 : _GEN_117; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_119 = 14'hc == parameter_2_2 ? phv_data_12 : _GEN_118; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_120 = 14'hd == parameter_2_2 ? phv_data_13 : _GEN_119; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_121 = 14'he == parameter_2_2 ? phv_data_14 : _GEN_120; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_122 = 14'hf == parameter_2_2 ? phv_data_15 : _GEN_121; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_123 = 14'h10 == parameter_2_2 ? phv_data_16 : _GEN_122; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_124 = 14'h11 == parameter_2_2 ? phv_data_17 : _GEN_123; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_125 = 14'h12 == parameter_2_2 ? phv_data_18 : _GEN_124; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_126 = 14'h13 == parameter_2_2 ? phv_data_19 : _GEN_125; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_127 = 14'h14 == parameter_2_2 ? phv_data_20 : _GEN_126; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_128 = 14'h15 == parameter_2_2 ? phv_data_21 : _GEN_127; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_129 = 14'h16 == parameter_2_2 ? phv_data_22 : _GEN_128; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_130 = 14'h17 == parameter_2_2 ? phv_data_23 : _GEN_129; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_131 = 14'h18 == parameter_2_2 ? phv_data_24 : _GEN_130; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_132 = 14'h19 == parameter_2_2 ? phv_data_25 : _GEN_131; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_133 = 14'h1a == parameter_2_2 ? phv_data_26 : _GEN_132; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_134 = 14'h1b == parameter_2_2 ? phv_data_27 : _GEN_133; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_135 = 14'h1c == parameter_2_2 ? phv_data_28 : _GEN_134; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_136 = 14'h1d == parameter_2_2 ? phv_data_29 : _GEN_135; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_137 = 14'h1e == parameter_2_2 ? phv_data_30 : _GEN_136; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_138 = 14'h1f == parameter_2_2 ? phv_data_31 : _GEN_137; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_3 = vliw_3[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_3 = vliw_3[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_3 = parameter_2_3[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_3 = parameter_2_3[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_3 = {{1'd0}, args_offset_3}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_3 = _total_offset_T_3[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_142 = 3'h1 == total_offset_3 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_143 = 3'h2 == total_offset_3 ? args_2 : _GEN_142; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_144 = 3'h3 == total_offset_3 ? args_3 : _GEN_143; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_145 = 3'h4 == total_offset_3 ? args_4 : _GEN_144; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_146 = 3'h5 == total_offset_3 ? args_5 : _GEN_145; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_147 = 3'h6 == total_offset_3 ? args_6 : _GEN_146; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_148 = total_offset_3 < 3'h7 ? _GEN_147 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_3_0 = 3'h0 < args_length_3 ? _GEN_148 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_150 = opcode_3 == 4'ha ? field_bytes_3_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_151 = opcode_3 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_120 = opcode_3 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_7 = _T_120 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_152 = opcode_3 == 4'h8 | opcode_3 == 4'hb ? parameter_2_3[7:0] : _GEN_150; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_153 = opcode_3 == 4'h8 | opcode_3 == 4'hb ? _field_tag_T_7 : _GEN_151; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_154 = 14'h0 == parameter_2_3 ? phv_data_0 : _GEN_152; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_155 = 14'h1 == parameter_2_3 ? phv_data_1 : _GEN_154; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_156 = 14'h2 == parameter_2_3 ? phv_data_2 : _GEN_155; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_157 = 14'h3 == parameter_2_3 ? phv_data_3 : _GEN_156; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_158 = 14'h4 == parameter_2_3 ? phv_data_4 : _GEN_157; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_159 = 14'h5 == parameter_2_3 ? phv_data_5 : _GEN_158; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_160 = 14'h6 == parameter_2_3 ? phv_data_6 : _GEN_159; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_161 = 14'h7 == parameter_2_3 ? phv_data_7 : _GEN_160; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_162 = 14'h8 == parameter_2_3 ? phv_data_8 : _GEN_161; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_163 = 14'h9 == parameter_2_3 ? phv_data_9 : _GEN_162; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_164 = 14'ha == parameter_2_3 ? phv_data_10 : _GEN_163; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_165 = 14'hb == parameter_2_3 ? phv_data_11 : _GEN_164; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_166 = 14'hc == parameter_2_3 ? phv_data_12 : _GEN_165; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_167 = 14'hd == parameter_2_3 ? phv_data_13 : _GEN_166; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_168 = 14'he == parameter_2_3 ? phv_data_14 : _GEN_167; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_169 = 14'hf == parameter_2_3 ? phv_data_15 : _GEN_168; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_170 = 14'h10 == parameter_2_3 ? phv_data_16 : _GEN_169; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_171 = 14'h11 == parameter_2_3 ? phv_data_17 : _GEN_170; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_172 = 14'h12 == parameter_2_3 ? phv_data_18 : _GEN_171; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_173 = 14'h13 == parameter_2_3 ? phv_data_19 : _GEN_172; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_174 = 14'h14 == parameter_2_3 ? phv_data_20 : _GEN_173; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_175 = 14'h15 == parameter_2_3 ? phv_data_21 : _GEN_174; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_176 = 14'h16 == parameter_2_3 ? phv_data_22 : _GEN_175; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_177 = 14'h17 == parameter_2_3 ? phv_data_23 : _GEN_176; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_178 = 14'h18 == parameter_2_3 ? phv_data_24 : _GEN_177; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_179 = 14'h19 == parameter_2_3 ? phv_data_25 : _GEN_178; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_180 = 14'h1a == parameter_2_3 ? phv_data_26 : _GEN_179; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_181 = 14'h1b == parameter_2_3 ? phv_data_27 : _GEN_180; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_182 = 14'h1c == parameter_2_3 ? phv_data_28 : _GEN_181; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_183 = 14'h1d == parameter_2_3 ? phv_data_29 : _GEN_182; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_184 = 14'h1e == parameter_2_3 ? phv_data_30 : _GEN_183; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_185 = 14'h1f == parameter_2_3 ? phv_data_31 : _GEN_184; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_4 = vliw_4[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_4 = vliw_4[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_4 = parameter_2_4[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_4 = parameter_2_4[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_4 = {{1'd0}, args_offset_4}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_4 = _total_offset_T_4[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_189 = 3'h1 == total_offset_4 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_190 = 3'h2 == total_offset_4 ? args_2 : _GEN_189; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_191 = 3'h3 == total_offset_4 ? args_3 : _GEN_190; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_192 = 3'h4 == total_offset_4 ? args_4 : _GEN_191; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_193 = 3'h5 == total_offset_4 ? args_5 : _GEN_192; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_194 = 3'h6 == total_offset_4 ? args_6 : _GEN_193; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_195 = total_offset_4 < 3'h7 ? _GEN_194 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_4_0 = 3'h0 < args_length_4 ? _GEN_195 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_197 = opcode_4 == 4'ha ? field_bytes_4_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_198 = opcode_4 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_159 = opcode_4 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_9 = _T_159 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_199 = opcode_4 == 4'h8 | opcode_4 == 4'hb ? parameter_2_4[7:0] : _GEN_197; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_200 = opcode_4 == 4'h8 | opcode_4 == 4'hb ? _field_tag_T_9 : _GEN_198; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_201 = 14'h0 == parameter_2_4 ? phv_data_0 : _GEN_199; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_202 = 14'h1 == parameter_2_4 ? phv_data_1 : _GEN_201; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_203 = 14'h2 == parameter_2_4 ? phv_data_2 : _GEN_202; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_204 = 14'h3 == parameter_2_4 ? phv_data_3 : _GEN_203; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_205 = 14'h4 == parameter_2_4 ? phv_data_4 : _GEN_204; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_206 = 14'h5 == parameter_2_4 ? phv_data_5 : _GEN_205; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_207 = 14'h6 == parameter_2_4 ? phv_data_6 : _GEN_206; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_208 = 14'h7 == parameter_2_4 ? phv_data_7 : _GEN_207; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_209 = 14'h8 == parameter_2_4 ? phv_data_8 : _GEN_208; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_210 = 14'h9 == parameter_2_4 ? phv_data_9 : _GEN_209; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_211 = 14'ha == parameter_2_4 ? phv_data_10 : _GEN_210; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_212 = 14'hb == parameter_2_4 ? phv_data_11 : _GEN_211; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_213 = 14'hc == parameter_2_4 ? phv_data_12 : _GEN_212; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_214 = 14'hd == parameter_2_4 ? phv_data_13 : _GEN_213; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_215 = 14'he == parameter_2_4 ? phv_data_14 : _GEN_214; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_216 = 14'hf == parameter_2_4 ? phv_data_15 : _GEN_215; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_217 = 14'h10 == parameter_2_4 ? phv_data_16 : _GEN_216; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_218 = 14'h11 == parameter_2_4 ? phv_data_17 : _GEN_217; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_219 = 14'h12 == parameter_2_4 ? phv_data_18 : _GEN_218; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_220 = 14'h13 == parameter_2_4 ? phv_data_19 : _GEN_219; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_221 = 14'h14 == parameter_2_4 ? phv_data_20 : _GEN_220; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_222 = 14'h15 == parameter_2_4 ? phv_data_21 : _GEN_221; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_223 = 14'h16 == parameter_2_4 ? phv_data_22 : _GEN_222; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_224 = 14'h17 == parameter_2_4 ? phv_data_23 : _GEN_223; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_225 = 14'h18 == parameter_2_4 ? phv_data_24 : _GEN_224; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_226 = 14'h19 == parameter_2_4 ? phv_data_25 : _GEN_225; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_227 = 14'h1a == parameter_2_4 ? phv_data_26 : _GEN_226; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_228 = 14'h1b == parameter_2_4 ? phv_data_27 : _GEN_227; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_229 = 14'h1c == parameter_2_4 ? phv_data_28 : _GEN_228; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_230 = 14'h1d == parameter_2_4 ? phv_data_29 : _GEN_229; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_231 = 14'h1e == parameter_2_4 ? phv_data_30 : _GEN_230; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_232 = 14'h1f == parameter_2_4 ? phv_data_31 : _GEN_231; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_5 = vliw_5[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_5 = vliw_5[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_5 = parameter_2_5[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_5 = parameter_2_5[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_5 = {{1'd0}, args_offset_5}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_5 = _total_offset_T_5[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_236 = 3'h1 == total_offset_5 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_237 = 3'h2 == total_offset_5 ? args_2 : _GEN_236; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_238 = 3'h3 == total_offset_5 ? args_3 : _GEN_237; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_239 = 3'h4 == total_offset_5 ? args_4 : _GEN_238; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_240 = 3'h5 == total_offset_5 ? args_5 : _GEN_239; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_241 = 3'h6 == total_offset_5 ? args_6 : _GEN_240; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_242 = total_offset_5 < 3'h7 ? _GEN_241 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_5_0 = 3'h0 < args_length_5 ? _GEN_242 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_244 = opcode_5 == 4'ha ? field_bytes_5_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_245 = opcode_5 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_198 = opcode_5 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_11 = _T_198 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_246 = opcode_5 == 4'h8 | opcode_5 == 4'hb ? parameter_2_5[7:0] : _GEN_244; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_247 = opcode_5 == 4'h8 | opcode_5 == 4'hb ? _field_tag_T_11 : _GEN_245; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_248 = 14'h0 == parameter_2_5 ? phv_data_0 : _GEN_246; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_249 = 14'h1 == parameter_2_5 ? phv_data_1 : _GEN_248; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_250 = 14'h2 == parameter_2_5 ? phv_data_2 : _GEN_249; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_251 = 14'h3 == parameter_2_5 ? phv_data_3 : _GEN_250; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_252 = 14'h4 == parameter_2_5 ? phv_data_4 : _GEN_251; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_253 = 14'h5 == parameter_2_5 ? phv_data_5 : _GEN_252; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_254 = 14'h6 == parameter_2_5 ? phv_data_6 : _GEN_253; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_255 = 14'h7 == parameter_2_5 ? phv_data_7 : _GEN_254; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_256 = 14'h8 == parameter_2_5 ? phv_data_8 : _GEN_255; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_257 = 14'h9 == parameter_2_5 ? phv_data_9 : _GEN_256; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_258 = 14'ha == parameter_2_5 ? phv_data_10 : _GEN_257; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_259 = 14'hb == parameter_2_5 ? phv_data_11 : _GEN_258; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_260 = 14'hc == parameter_2_5 ? phv_data_12 : _GEN_259; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_261 = 14'hd == parameter_2_5 ? phv_data_13 : _GEN_260; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_262 = 14'he == parameter_2_5 ? phv_data_14 : _GEN_261; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_263 = 14'hf == parameter_2_5 ? phv_data_15 : _GEN_262; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_264 = 14'h10 == parameter_2_5 ? phv_data_16 : _GEN_263; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_265 = 14'h11 == parameter_2_5 ? phv_data_17 : _GEN_264; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_266 = 14'h12 == parameter_2_5 ? phv_data_18 : _GEN_265; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_267 = 14'h13 == parameter_2_5 ? phv_data_19 : _GEN_266; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_268 = 14'h14 == parameter_2_5 ? phv_data_20 : _GEN_267; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_269 = 14'h15 == parameter_2_5 ? phv_data_21 : _GEN_268; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_270 = 14'h16 == parameter_2_5 ? phv_data_22 : _GEN_269; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_271 = 14'h17 == parameter_2_5 ? phv_data_23 : _GEN_270; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_272 = 14'h18 == parameter_2_5 ? phv_data_24 : _GEN_271; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_273 = 14'h19 == parameter_2_5 ? phv_data_25 : _GEN_272; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_274 = 14'h1a == parameter_2_5 ? phv_data_26 : _GEN_273; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_275 = 14'h1b == parameter_2_5 ? phv_data_27 : _GEN_274; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_276 = 14'h1c == parameter_2_5 ? phv_data_28 : _GEN_275; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_277 = 14'h1d == parameter_2_5 ? phv_data_29 : _GEN_276; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_278 = 14'h1e == parameter_2_5 ? phv_data_30 : _GEN_277; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_279 = 14'h1f == parameter_2_5 ? phv_data_31 : _GEN_278; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_6 = vliw_6[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_6 = vliw_6[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_6 = parameter_2_6[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_6 = parameter_2_6[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_6 = {{1'd0}, args_offset_6}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_6 = _total_offset_T_6[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_283 = 3'h1 == total_offset_6 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_284 = 3'h2 == total_offset_6 ? args_2 : _GEN_283; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_285 = 3'h3 == total_offset_6 ? args_3 : _GEN_284; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_286 = 3'h4 == total_offset_6 ? args_4 : _GEN_285; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_287 = 3'h5 == total_offset_6 ? args_5 : _GEN_286; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_288 = 3'h6 == total_offset_6 ? args_6 : _GEN_287; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_289 = total_offset_6 < 3'h7 ? _GEN_288 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_6_0 = 3'h0 < args_length_6 ? _GEN_289 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_291 = opcode_6 == 4'ha ? field_bytes_6_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_292 = opcode_6 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_237 = opcode_6 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_13 = _T_237 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_293 = opcode_6 == 4'h8 | opcode_6 == 4'hb ? parameter_2_6[7:0] : _GEN_291; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_294 = opcode_6 == 4'h8 | opcode_6 == 4'hb ? _field_tag_T_13 : _GEN_292; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_295 = 14'h0 == parameter_2_6 ? phv_data_0 : _GEN_293; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_296 = 14'h1 == parameter_2_6 ? phv_data_1 : _GEN_295; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_297 = 14'h2 == parameter_2_6 ? phv_data_2 : _GEN_296; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_298 = 14'h3 == parameter_2_6 ? phv_data_3 : _GEN_297; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_299 = 14'h4 == parameter_2_6 ? phv_data_4 : _GEN_298; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_300 = 14'h5 == parameter_2_6 ? phv_data_5 : _GEN_299; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_301 = 14'h6 == parameter_2_6 ? phv_data_6 : _GEN_300; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_302 = 14'h7 == parameter_2_6 ? phv_data_7 : _GEN_301; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_303 = 14'h8 == parameter_2_6 ? phv_data_8 : _GEN_302; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_304 = 14'h9 == parameter_2_6 ? phv_data_9 : _GEN_303; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_305 = 14'ha == parameter_2_6 ? phv_data_10 : _GEN_304; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_306 = 14'hb == parameter_2_6 ? phv_data_11 : _GEN_305; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_307 = 14'hc == parameter_2_6 ? phv_data_12 : _GEN_306; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_308 = 14'hd == parameter_2_6 ? phv_data_13 : _GEN_307; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_309 = 14'he == parameter_2_6 ? phv_data_14 : _GEN_308; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_310 = 14'hf == parameter_2_6 ? phv_data_15 : _GEN_309; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_311 = 14'h10 == parameter_2_6 ? phv_data_16 : _GEN_310; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_312 = 14'h11 == parameter_2_6 ? phv_data_17 : _GEN_311; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_313 = 14'h12 == parameter_2_6 ? phv_data_18 : _GEN_312; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_314 = 14'h13 == parameter_2_6 ? phv_data_19 : _GEN_313; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_315 = 14'h14 == parameter_2_6 ? phv_data_20 : _GEN_314; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_316 = 14'h15 == parameter_2_6 ? phv_data_21 : _GEN_315; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_317 = 14'h16 == parameter_2_6 ? phv_data_22 : _GEN_316; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_318 = 14'h17 == parameter_2_6 ? phv_data_23 : _GEN_317; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_319 = 14'h18 == parameter_2_6 ? phv_data_24 : _GEN_318; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_320 = 14'h19 == parameter_2_6 ? phv_data_25 : _GEN_319; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_321 = 14'h1a == parameter_2_6 ? phv_data_26 : _GEN_320; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_322 = 14'h1b == parameter_2_6 ? phv_data_27 : _GEN_321; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_323 = 14'h1c == parameter_2_6 ? phv_data_28 : _GEN_322; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_324 = 14'h1d == parameter_2_6 ? phv_data_29 : _GEN_323; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_325 = 14'h1e == parameter_2_6 ? phv_data_30 : _GEN_324; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_326 = 14'h1f == parameter_2_6 ? phv_data_31 : _GEN_325; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_7 = vliw_7[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_7 = vliw_7[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_7 = parameter_2_7[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_7 = parameter_2_7[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_7 = {{1'd0}, args_offset_7}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_7 = _total_offset_T_7[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_330 = 3'h1 == total_offset_7 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_331 = 3'h2 == total_offset_7 ? args_2 : _GEN_330; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_332 = 3'h3 == total_offset_7 ? args_3 : _GEN_331; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_333 = 3'h4 == total_offset_7 ? args_4 : _GEN_332; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_334 = 3'h5 == total_offset_7 ? args_5 : _GEN_333; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_335 = 3'h6 == total_offset_7 ? args_6 : _GEN_334; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_336 = total_offset_7 < 3'h7 ? _GEN_335 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_7_0 = 3'h0 < args_length_7 ? _GEN_336 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_338 = opcode_7 == 4'ha ? field_bytes_7_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_339 = opcode_7 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_276 = opcode_7 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_15 = _T_276 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_340 = opcode_7 == 4'h8 | opcode_7 == 4'hb ? parameter_2_7[7:0] : _GEN_338; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_341 = opcode_7 == 4'h8 | opcode_7 == 4'hb ? _field_tag_T_15 : _GEN_339; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_342 = 14'h0 == parameter_2_7 ? phv_data_0 : _GEN_340; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_343 = 14'h1 == parameter_2_7 ? phv_data_1 : _GEN_342; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_344 = 14'h2 == parameter_2_7 ? phv_data_2 : _GEN_343; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_345 = 14'h3 == parameter_2_7 ? phv_data_3 : _GEN_344; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_346 = 14'h4 == parameter_2_7 ? phv_data_4 : _GEN_345; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_347 = 14'h5 == parameter_2_7 ? phv_data_5 : _GEN_346; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_348 = 14'h6 == parameter_2_7 ? phv_data_6 : _GEN_347; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_349 = 14'h7 == parameter_2_7 ? phv_data_7 : _GEN_348; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_350 = 14'h8 == parameter_2_7 ? phv_data_8 : _GEN_349; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_351 = 14'h9 == parameter_2_7 ? phv_data_9 : _GEN_350; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_352 = 14'ha == parameter_2_7 ? phv_data_10 : _GEN_351; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_353 = 14'hb == parameter_2_7 ? phv_data_11 : _GEN_352; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_354 = 14'hc == parameter_2_7 ? phv_data_12 : _GEN_353; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_355 = 14'hd == parameter_2_7 ? phv_data_13 : _GEN_354; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_356 = 14'he == parameter_2_7 ? phv_data_14 : _GEN_355; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_357 = 14'hf == parameter_2_7 ? phv_data_15 : _GEN_356; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_358 = 14'h10 == parameter_2_7 ? phv_data_16 : _GEN_357; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_359 = 14'h11 == parameter_2_7 ? phv_data_17 : _GEN_358; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_360 = 14'h12 == parameter_2_7 ? phv_data_18 : _GEN_359; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_361 = 14'h13 == parameter_2_7 ? phv_data_19 : _GEN_360; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_362 = 14'h14 == parameter_2_7 ? phv_data_20 : _GEN_361; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_363 = 14'h15 == parameter_2_7 ? phv_data_21 : _GEN_362; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_364 = 14'h16 == parameter_2_7 ? phv_data_22 : _GEN_363; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_365 = 14'h17 == parameter_2_7 ? phv_data_23 : _GEN_364; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_366 = 14'h18 == parameter_2_7 ? phv_data_24 : _GEN_365; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_367 = 14'h19 == parameter_2_7 ? phv_data_25 : _GEN_366; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_368 = 14'h1a == parameter_2_7 ? phv_data_26 : _GEN_367; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_369 = 14'h1b == parameter_2_7 ? phv_data_27 : _GEN_368; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_370 = 14'h1c == parameter_2_7 ? phv_data_28 : _GEN_369; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_371 = 14'h1d == parameter_2_7 ? phv_data_29 : _GEN_370; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_372 = 14'h1e == parameter_2_7 ? phv_data_30 : _GEN_371; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_373 = 14'h1f == parameter_2_7 ? phv_data_31 : _GEN_372; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_8 = vliw_8[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_8 = vliw_8[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_8 = parameter_2_8[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_8 = parameter_2_8[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_8 = {{1'd0}, args_offset_8}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_8 = _total_offset_T_8[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_377 = 3'h1 == total_offset_8 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_378 = 3'h2 == total_offset_8 ? args_2 : _GEN_377; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_379 = 3'h3 == total_offset_8 ? args_3 : _GEN_378; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_380 = 3'h4 == total_offset_8 ? args_4 : _GEN_379; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_381 = 3'h5 == total_offset_8 ? args_5 : _GEN_380; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_382 = 3'h6 == total_offset_8 ? args_6 : _GEN_381; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_383 = total_offset_8 < 3'h7 ? _GEN_382 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_8_0 = 3'h0 < args_length_8 ? _GEN_383 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_385 = opcode_8 == 4'ha ? field_bytes_8_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_386 = opcode_8 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_315 = opcode_8 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_17 = _T_315 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_387 = opcode_8 == 4'h8 | opcode_8 == 4'hb ? parameter_2_8[7:0] : _GEN_385; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_388 = opcode_8 == 4'h8 | opcode_8 == 4'hb ? _field_tag_T_17 : _GEN_386; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_389 = 14'h0 == parameter_2_8 ? phv_data_0 : _GEN_387; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_390 = 14'h1 == parameter_2_8 ? phv_data_1 : _GEN_389; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_391 = 14'h2 == parameter_2_8 ? phv_data_2 : _GEN_390; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_392 = 14'h3 == parameter_2_8 ? phv_data_3 : _GEN_391; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_393 = 14'h4 == parameter_2_8 ? phv_data_4 : _GEN_392; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_394 = 14'h5 == parameter_2_8 ? phv_data_5 : _GEN_393; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_395 = 14'h6 == parameter_2_8 ? phv_data_6 : _GEN_394; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_396 = 14'h7 == parameter_2_8 ? phv_data_7 : _GEN_395; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_397 = 14'h8 == parameter_2_8 ? phv_data_8 : _GEN_396; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_398 = 14'h9 == parameter_2_8 ? phv_data_9 : _GEN_397; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_399 = 14'ha == parameter_2_8 ? phv_data_10 : _GEN_398; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_400 = 14'hb == parameter_2_8 ? phv_data_11 : _GEN_399; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_401 = 14'hc == parameter_2_8 ? phv_data_12 : _GEN_400; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_402 = 14'hd == parameter_2_8 ? phv_data_13 : _GEN_401; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_403 = 14'he == parameter_2_8 ? phv_data_14 : _GEN_402; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_404 = 14'hf == parameter_2_8 ? phv_data_15 : _GEN_403; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_405 = 14'h10 == parameter_2_8 ? phv_data_16 : _GEN_404; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_406 = 14'h11 == parameter_2_8 ? phv_data_17 : _GEN_405; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_407 = 14'h12 == parameter_2_8 ? phv_data_18 : _GEN_406; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_408 = 14'h13 == parameter_2_8 ? phv_data_19 : _GEN_407; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_409 = 14'h14 == parameter_2_8 ? phv_data_20 : _GEN_408; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_410 = 14'h15 == parameter_2_8 ? phv_data_21 : _GEN_409; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_411 = 14'h16 == parameter_2_8 ? phv_data_22 : _GEN_410; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_412 = 14'h17 == parameter_2_8 ? phv_data_23 : _GEN_411; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_413 = 14'h18 == parameter_2_8 ? phv_data_24 : _GEN_412; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_414 = 14'h19 == parameter_2_8 ? phv_data_25 : _GEN_413; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_415 = 14'h1a == parameter_2_8 ? phv_data_26 : _GEN_414; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_416 = 14'h1b == parameter_2_8 ? phv_data_27 : _GEN_415; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_417 = 14'h1c == parameter_2_8 ? phv_data_28 : _GEN_416; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_418 = 14'h1d == parameter_2_8 ? phv_data_29 : _GEN_417; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_419 = 14'h1e == parameter_2_8 ? phv_data_30 : _GEN_418; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_420 = 14'h1f == parameter_2_8 ? phv_data_31 : _GEN_419; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_9 = vliw_9[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_9 = vliw_9[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_9 = parameter_2_9[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_9 = parameter_2_9[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_9 = {{1'd0}, args_offset_9}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_9 = _total_offset_T_9[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_424 = 3'h1 == total_offset_9 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_425 = 3'h2 == total_offset_9 ? args_2 : _GEN_424; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_426 = 3'h3 == total_offset_9 ? args_3 : _GEN_425; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_427 = 3'h4 == total_offset_9 ? args_4 : _GEN_426; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_428 = 3'h5 == total_offset_9 ? args_5 : _GEN_427; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_429 = 3'h6 == total_offset_9 ? args_6 : _GEN_428; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_430 = total_offset_9 < 3'h7 ? _GEN_429 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_9_0 = 3'h0 < args_length_9 ? _GEN_430 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_432 = opcode_9 == 4'ha ? field_bytes_9_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_433 = opcode_9 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_354 = opcode_9 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_19 = _T_354 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_434 = opcode_9 == 4'h8 | opcode_9 == 4'hb ? parameter_2_9[7:0] : _GEN_432; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_435 = opcode_9 == 4'h8 | opcode_9 == 4'hb ? _field_tag_T_19 : _GEN_433; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_436 = 14'h0 == parameter_2_9 ? phv_data_0 : _GEN_434; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_437 = 14'h1 == parameter_2_9 ? phv_data_1 : _GEN_436; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_438 = 14'h2 == parameter_2_9 ? phv_data_2 : _GEN_437; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_439 = 14'h3 == parameter_2_9 ? phv_data_3 : _GEN_438; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_440 = 14'h4 == parameter_2_9 ? phv_data_4 : _GEN_439; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_441 = 14'h5 == parameter_2_9 ? phv_data_5 : _GEN_440; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_442 = 14'h6 == parameter_2_9 ? phv_data_6 : _GEN_441; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_443 = 14'h7 == parameter_2_9 ? phv_data_7 : _GEN_442; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_444 = 14'h8 == parameter_2_9 ? phv_data_8 : _GEN_443; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_445 = 14'h9 == parameter_2_9 ? phv_data_9 : _GEN_444; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_446 = 14'ha == parameter_2_9 ? phv_data_10 : _GEN_445; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_447 = 14'hb == parameter_2_9 ? phv_data_11 : _GEN_446; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_448 = 14'hc == parameter_2_9 ? phv_data_12 : _GEN_447; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_449 = 14'hd == parameter_2_9 ? phv_data_13 : _GEN_448; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_450 = 14'he == parameter_2_9 ? phv_data_14 : _GEN_449; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_451 = 14'hf == parameter_2_9 ? phv_data_15 : _GEN_450; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_452 = 14'h10 == parameter_2_9 ? phv_data_16 : _GEN_451; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_453 = 14'h11 == parameter_2_9 ? phv_data_17 : _GEN_452; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_454 = 14'h12 == parameter_2_9 ? phv_data_18 : _GEN_453; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_455 = 14'h13 == parameter_2_9 ? phv_data_19 : _GEN_454; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_456 = 14'h14 == parameter_2_9 ? phv_data_20 : _GEN_455; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_457 = 14'h15 == parameter_2_9 ? phv_data_21 : _GEN_456; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_458 = 14'h16 == parameter_2_9 ? phv_data_22 : _GEN_457; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_459 = 14'h17 == parameter_2_9 ? phv_data_23 : _GEN_458; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_460 = 14'h18 == parameter_2_9 ? phv_data_24 : _GEN_459; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_461 = 14'h19 == parameter_2_9 ? phv_data_25 : _GEN_460; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_462 = 14'h1a == parameter_2_9 ? phv_data_26 : _GEN_461; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_463 = 14'h1b == parameter_2_9 ? phv_data_27 : _GEN_462; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_464 = 14'h1c == parameter_2_9 ? phv_data_28 : _GEN_463; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_465 = 14'h1d == parameter_2_9 ? phv_data_29 : _GEN_464; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_466 = 14'h1e == parameter_2_9 ? phv_data_30 : _GEN_465; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_467 = 14'h1f == parameter_2_9 ? phv_data_31 : _GEN_466; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_10 = vliw_10[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_10 = vliw_10[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_10 = parameter_2_10[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_10 = parameter_2_10[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_10 = {{1'd0}, args_offset_10}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_10 = _total_offset_T_10[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_471 = 3'h1 == total_offset_10 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_472 = 3'h2 == total_offset_10 ? args_2 : _GEN_471; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_473 = 3'h3 == total_offset_10 ? args_3 : _GEN_472; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_474 = 3'h4 == total_offset_10 ? args_4 : _GEN_473; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_475 = 3'h5 == total_offset_10 ? args_5 : _GEN_474; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_476 = 3'h6 == total_offset_10 ? args_6 : _GEN_475; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_477 = total_offset_10 < 3'h7 ? _GEN_476 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_10_0 = 3'h0 < args_length_10 ? _GEN_477 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_479 = opcode_10 == 4'ha ? field_bytes_10_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_480 = opcode_10 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_393 = opcode_10 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_21 = _T_393 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_481 = opcode_10 == 4'h8 | opcode_10 == 4'hb ? parameter_2_10[7:0] : _GEN_479; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_482 = opcode_10 == 4'h8 | opcode_10 == 4'hb ? _field_tag_T_21 : _GEN_480; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_483 = 14'h0 == parameter_2_10 ? phv_data_0 : _GEN_481; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_484 = 14'h1 == parameter_2_10 ? phv_data_1 : _GEN_483; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_485 = 14'h2 == parameter_2_10 ? phv_data_2 : _GEN_484; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_486 = 14'h3 == parameter_2_10 ? phv_data_3 : _GEN_485; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_487 = 14'h4 == parameter_2_10 ? phv_data_4 : _GEN_486; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_488 = 14'h5 == parameter_2_10 ? phv_data_5 : _GEN_487; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_489 = 14'h6 == parameter_2_10 ? phv_data_6 : _GEN_488; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_490 = 14'h7 == parameter_2_10 ? phv_data_7 : _GEN_489; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_491 = 14'h8 == parameter_2_10 ? phv_data_8 : _GEN_490; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_492 = 14'h9 == parameter_2_10 ? phv_data_9 : _GEN_491; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_493 = 14'ha == parameter_2_10 ? phv_data_10 : _GEN_492; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_494 = 14'hb == parameter_2_10 ? phv_data_11 : _GEN_493; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_495 = 14'hc == parameter_2_10 ? phv_data_12 : _GEN_494; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_496 = 14'hd == parameter_2_10 ? phv_data_13 : _GEN_495; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_497 = 14'he == parameter_2_10 ? phv_data_14 : _GEN_496; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_498 = 14'hf == parameter_2_10 ? phv_data_15 : _GEN_497; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_499 = 14'h10 == parameter_2_10 ? phv_data_16 : _GEN_498; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_500 = 14'h11 == parameter_2_10 ? phv_data_17 : _GEN_499; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_501 = 14'h12 == parameter_2_10 ? phv_data_18 : _GEN_500; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_502 = 14'h13 == parameter_2_10 ? phv_data_19 : _GEN_501; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_503 = 14'h14 == parameter_2_10 ? phv_data_20 : _GEN_502; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_504 = 14'h15 == parameter_2_10 ? phv_data_21 : _GEN_503; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_505 = 14'h16 == parameter_2_10 ? phv_data_22 : _GEN_504; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_506 = 14'h17 == parameter_2_10 ? phv_data_23 : _GEN_505; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_507 = 14'h18 == parameter_2_10 ? phv_data_24 : _GEN_506; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_508 = 14'h19 == parameter_2_10 ? phv_data_25 : _GEN_507; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_509 = 14'h1a == parameter_2_10 ? phv_data_26 : _GEN_508; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_510 = 14'h1b == parameter_2_10 ? phv_data_27 : _GEN_509; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_511 = 14'h1c == parameter_2_10 ? phv_data_28 : _GEN_510; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_512 = 14'h1d == parameter_2_10 ? phv_data_29 : _GEN_511; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_513 = 14'h1e == parameter_2_10 ? phv_data_30 : _GEN_512; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_514 = 14'h1f == parameter_2_10 ? phv_data_31 : _GEN_513; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_11 = vliw_11[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_11 = vliw_11[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_11 = parameter_2_11[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_11 = parameter_2_11[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_11 = {{1'd0}, args_offset_11}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_11 = _total_offset_T_11[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_518 = 3'h1 == total_offset_11 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_519 = 3'h2 == total_offset_11 ? args_2 : _GEN_518; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_520 = 3'h3 == total_offset_11 ? args_3 : _GEN_519; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_521 = 3'h4 == total_offset_11 ? args_4 : _GEN_520; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_522 = 3'h5 == total_offset_11 ? args_5 : _GEN_521; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_523 = 3'h6 == total_offset_11 ? args_6 : _GEN_522; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_524 = total_offset_11 < 3'h7 ? _GEN_523 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_11_0 = 3'h0 < args_length_11 ? _GEN_524 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_526 = opcode_11 == 4'ha ? field_bytes_11_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_527 = opcode_11 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_432 = opcode_11 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_23 = _T_432 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_528 = opcode_11 == 4'h8 | opcode_11 == 4'hb ? parameter_2_11[7:0] : _GEN_526; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_529 = opcode_11 == 4'h8 | opcode_11 == 4'hb ? _field_tag_T_23 : _GEN_527; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_530 = 14'h0 == parameter_2_11 ? phv_data_0 : _GEN_528; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_531 = 14'h1 == parameter_2_11 ? phv_data_1 : _GEN_530; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_532 = 14'h2 == parameter_2_11 ? phv_data_2 : _GEN_531; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_533 = 14'h3 == parameter_2_11 ? phv_data_3 : _GEN_532; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_534 = 14'h4 == parameter_2_11 ? phv_data_4 : _GEN_533; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_535 = 14'h5 == parameter_2_11 ? phv_data_5 : _GEN_534; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_536 = 14'h6 == parameter_2_11 ? phv_data_6 : _GEN_535; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_537 = 14'h7 == parameter_2_11 ? phv_data_7 : _GEN_536; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_538 = 14'h8 == parameter_2_11 ? phv_data_8 : _GEN_537; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_539 = 14'h9 == parameter_2_11 ? phv_data_9 : _GEN_538; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_540 = 14'ha == parameter_2_11 ? phv_data_10 : _GEN_539; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_541 = 14'hb == parameter_2_11 ? phv_data_11 : _GEN_540; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_542 = 14'hc == parameter_2_11 ? phv_data_12 : _GEN_541; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_543 = 14'hd == parameter_2_11 ? phv_data_13 : _GEN_542; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_544 = 14'he == parameter_2_11 ? phv_data_14 : _GEN_543; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_545 = 14'hf == parameter_2_11 ? phv_data_15 : _GEN_544; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_546 = 14'h10 == parameter_2_11 ? phv_data_16 : _GEN_545; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_547 = 14'h11 == parameter_2_11 ? phv_data_17 : _GEN_546; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_548 = 14'h12 == parameter_2_11 ? phv_data_18 : _GEN_547; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_549 = 14'h13 == parameter_2_11 ? phv_data_19 : _GEN_548; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_550 = 14'h14 == parameter_2_11 ? phv_data_20 : _GEN_549; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_551 = 14'h15 == parameter_2_11 ? phv_data_21 : _GEN_550; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_552 = 14'h16 == parameter_2_11 ? phv_data_22 : _GEN_551; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_553 = 14'h17 == parameter_2_11 ? phv_data_23 : _GEN_552; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_554 = 14'h18 == parameter_2_11 ? phv_data_24 : _GEN_553; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_555 = 14'h19 == parameter_2_11 ? phv_data_25 : _GEN_554; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_556 = 14'h1a == parameter_2_11 ? phv_data_26 : _GEN_555; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_557 = 14'h1b == parameter_2_11 ? phv_data_27 : _GEN_556; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_558 = 14'h1c == parameter_2_11 ? phv_data_28 : _GEN_557; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_559 = 14'h1d == parameter_2_11 ? phv_data_29 : _GEN_558; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_560 = 14'h1e == parameter_2_11 ? phv_data_30 : _GEN_559; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_561 = 14'h1f == parameter_2_11 ? phv_data_31 : _GEN_560; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_12 = vliw_12[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_12 = vliw_12[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_12 = parameter_2_12[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_12 = parameter_2_12[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_12 = {{1'd0}, args_offset_12}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_12 = _total_offset_T_12[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_565 = 3'h1 == total_offset_12 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_566 = 3'h2 == total_offset_12 ? args_2 : _GEN_565; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_567 = 3'h3 == total_offset_12 ? args_3 : _GEN_566; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_568 = 3'h4 == total_offset_12 ? args_4 : _GEN_567; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_569 = 3'h5 == total_offset_12 ? args_5 : _GEN_568; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_570 = 3'h6 == total_offset_12 ? args_6 : _GEN_569; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_571 = total_offset_12 < 3'h7 ? _GEN_570 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_12_0 = 3'h0 < args_length_12 ? _GEN_571 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_573 = opcode_12 == 4'ha ? field_bytes_12_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_574 = opcode_12 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_471 = opcode_12 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_25 = _T_471 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_575 = opcode_12 == 4'h8 | opcode_12 == 4'hb ? parameter_2_12[7:0] : _GEN_573; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_576 = opcode_12 == 4'h8 | opcode_12 == 4'hb ? _field_tag_T_25 : _GEN_574; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_577 = 14'h0 == parameter_2_12 ? phv_data_0 : _GEN_575; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_578 = 14'h1 == parameter_2_12 ? phv_data_1 : _GEN_577; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_579 = 14'h2 == parameter_2_12 ? phv_data_2 : _GEN_578; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_580 = 14'h3 == parameter_2_12 ? phv_data_3 : _GEN_579; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_581 = 14'h4 == parameter_2_12 ? phv_data_4 : _GEN_580; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_582 = 14'h5 == parameter_2_12 ? phv_data_5 : _GEN_581; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_583 = 14'h6 == parameter_2_12 ? phv_data_6 : _GEN_582; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_584 = 14'h7 == parameter_2_12 ? phv_data_7 : _GEN_583; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_585 = 14'h8 == parameter_2_12 ? phv_data_8 : _GEN_584; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_586 = 14'h9 == parameter_2_12 ? phv_data_9 : _GEN_585; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_587 = 14'ha == parameter_2_12 ? phv_data_10 : _GEN_586; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_588 = 14'hb == parameter_2_12 ? phv_data_11 : _GEN_587; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_589 = 14'hc == parameter_2_12 ? phv_data_12 : _GEN_588; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_590 = 14'hd == parameter_2_12 ? phv_data_13 : _GEN_589; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_591 = 14'he == parameter_2_12 ? phv_data_14 : _GEN_590; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_592 = 14'hf == parameter_2_12 ? phv_data_15 : _GEN_591; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_593 = 14'h10 == parameter_2_12 ? phv_data_16 : _GEN_592; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_594 = 14'h11 == parameter_2_12 ? phv_data_17 : _GEN_593; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_595 = 14'h12 == parameter_2_12 ? phv_data_18 : _GEN_594; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_596 = 14'h13 == parameter_2_12 ? phv_data_19 : _GEN_595; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_597 = 14'h14 == parameter_2_12 ? phv_data_20 : _GEN_596; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_598 = 14'h15 == parameter_2_12 ? phv_data_21 : _GEN_597; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_599 = 14'h16 == parameter_2_12 ? phv_data_22 : _GEN_598; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_600 = 14'h17 == parameter_2_12 ? phv_data_23 : _GEN_599; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_601 = 14'h18 == parameter_2_12 ? phv_data_24 : _GEN_600; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_602 = 14'h19 == parameter_2_12 ? phv_data_25 : _GEN_601; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_603 = 14'h1a == parameter_2_12 ? phv_data_26 : _GEN_602; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_604 = 14'h1b == parameter_2_12 ? phv_data_27 : _GEN_603; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_605 = 14'h1c == parameter_2_12 ? phv_data_28 : _GEN_604; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_606 = 14'h1d == parameter_2_12 ? phv_data_29 : _GEN_605; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_607 = 14'h1e == parameter_2_12 ? phv_data_30 : _GEN_606; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_608 = 14'h1f == parameter_2_12 ? phv_data_31 : _GEN_607; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_13 = vliw_13[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_13 = vliw_13[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_13 = parameter_2_13[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_13 = parameter_2_13[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_13 = {{1'd0}, args_offset_13}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_13 = _total_offset_T_13[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_612 = 3'h1 == total_offset_13 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_613 = 3'h2 == total_offset_13 ? args_2 : _GEN_612; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_614 = 3'h3 == total_offset_13 ? args_3 : _GEN_613; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_615 = 3'h4 == total_offset_13 ? args_4 : _GEN_614; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_616 = 3'h5 == total_offset_13 ? args_5 : _GEN_615; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_617 = 3'h6 == total_offset_13 ? args_6 : _GEN_616; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_618 = total_offset_13 < 3'h7 ? _GEN_617 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_13_0 = 3'h0 < args_length_13 ? _GEN_618 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_620 = opcode_13 == 4'ha ? field_bytes_13_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_621 = opcode_13 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_510 = opcode_13 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_27 = _T_510 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_622 = opcode_13 == 4'h8 | opcode_13 == 4'hb ? parameter_2_13[7:0] : _GEN_620; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_623 = opcode_13 == 4'h8 | opcode_13 == 4'hb ? _field_tag_T_27 : _GEN_621; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_624 = 14'h0 == parameter_2_13 ? phv_data_0 : _GEN_622; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_625 = 14'h1 == parameter_2_13 ? phv_data_1 : _GEN_624; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_626 = 14'h2 == parameter_2_13 ? phv_data_2 : _GEN_625; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_627 = 14'h3 == parameter_2_13 ? phv_data_3 : _GEN_626; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_628 = 14'h4 == parameter_2_13 ? phv_data_4 : _GEN_627; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_629 = 14'h5 == parameter_2_13 ? phv_data_5 : _GEN_628; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_630 = 14'h6 == parameter_2_13 ? phv_data_6 : _GEN_629; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_631 = 14'h7 == parameter_2_13 ? phv_data_7 : _GEN_630; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_632 = 14'h8 == parameter_2_13 ? phv_data_8 : _GEN_631; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_633 = 14'h9 == parameter_2_13 ? phv_data_9 : _GEN_632; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_634 = 14'ha == parameter_2_13 ? phv_data_10 : _GEN_633; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_635 = 14'hb == parameter_2_13 ? phv_data_11 : _GEN_634; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_636 = 14'hc == parameter_2_13 ? phv_data_12 : _GEN_635; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_637 = 14'hd == parameter_2_13 ? phv_data_13 : _GEN_636; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_638 = 14'he == parameter_2_13 ? phv_data_14 : _GEN_637; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_639 = 14'hf == parameter_2_13 ? phv_data_15 : _GEN_638; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_640 = 14'h10 == parameter_2_13 ? phv_data_16 : _GEN_639; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_641 = 14'h11 == parameter_2_13 ? phv_data_17 : _GEN_640; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_642 = 14'h12 == parameter_2_13 ? phv_data_18 : _GEN_641; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_643 = 14'h13 == parameter_2_13 ? phv_data_19 : _GEN_642; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_644 = 14'h14 == parameter_2_13 ? phv_data_20 : _GEN_643; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_645 = 14'h15 == parameter_2_13 ? phv_data_21 : _GEN_644; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_646 = 14'h16 == parameter_2_13 ? phv_data_22 : _GEN_645; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_647 = 14'h17 == parameter_2_13 ? phv_data_23 : _GEN_646; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_648 = 14'h18 == parameter_2_13 ? phv_data_24 : _GEN_647; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_649 = 14'h19 == parameter_2_13 ? phv_data_25 : _GEN_648; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_650 = 14'h1a == parameter_2_13 ? phv_data_26 : _GEN_649; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_651 = 14'h1b == parameter_2_13 ? phv_data_27 : _GEN_650; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_652 = 14'h1c == parameter_2_13 ? phv_data_28 : _GEN_651; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_653 = 14'h1d == parameter_2_13 ? phv_data_29 : _GEN_652; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_654 = 14'h1e == parameter_2_13 ? phv_data_30 : _GEN_653; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_655 = 14'h1f == parameter_2_13 ? phv_data_31 : _GEN_654; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_14 = vliw_14[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_14 = vliw_14[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_14 = parameter_2_14[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_14 = parameter_2_14[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_14 = {{1'd0}, args_offset_14}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_14 = _total_offset_T_14[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_659 = 3'h1 == total_offset_14 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_660 = 3'h2 == total_offset_14 ? args_2 : _GEN_659; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_661 = 3'h3 == total_offset_14 ? args_3 : _GEN_660; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_662 = 3'h4 == total_offset_14 ? args_4 : _GEN_661; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_663 = 3'h5 == total_offset_14 ? args_5 : _GEN_662; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_664 = 3'h6 == total_offset_14 ? args_6 : _GEN_663; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_665 = total_offset_14 < 3'h7 ? _GEN_664 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_14_0 = 3'h0 < args_length_14 ? _GEN_665 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_667 = opcode_14 == 4'ha ? field_bytes_14_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_668 = opcode_14 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_549 = opcode_14 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_29 = _T_549 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_669 = opcode_14 == 4'h8 | opcode_14 == 4'hb ? parameter_2_14[7:0] : _GEN_667; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_670 = opcode_14 == 4'h8 | opcode_14 == 4'hb ? _field_tag_T_29 : _GEN_668; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_671 = 14'h0 == parameter_2_14 ? phv_data_0 : _GEN_669; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_672 = 14'h1 == parameter_2_14 ? phv_data_1 : _GEN_671; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_673 = 14'h2 == parameter_2_14 ? phv_data_2 : _GEN_672; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_674 = 14'h3 == parameter_2_14 ? phv_data_3 : _GEN_673; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_675 = 14'h4 == parameter_2_14 ? phv_data_4 : _GEN_674; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_676 = 14'h5 == parameter_2_14 ? phv_data_5 : _GEN_675; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_677 = 14'h6 == parameter_2_14 ? phv_data_6 : _GEN_676; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_678 = 14'h7 == parameter_2_14 ? phv_data_7 : _GEN_677; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_679 = 14'h8 == parameter_2_14 ? phv_data_8 : _GEN_678; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_680 = 14'h9 == parameter_2_14 ? phv_data_9 : _GEN_679; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_681 = 14'ha == parameter_2_14 ? phv_data_10 : _GEN_680; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_682 = 14'hb == parameter_2_14 ? phv_data_11 : _GEN_681; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_683 = 14'hc == parameter_2_14 ? phv_data_12 : _GEN_682; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_684 = 14'hd == parameter_2_14 ? phv_data_13 : _GEN_683; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_685 = 14'he == parameter_2_14 ? phv_data_14 : _GEN_684; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_686 = 14'hf == parameter_2_14 ? phv_data_15 : _GEN_685; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_687 = 14'h10 == parameter_2_14 ? phv_data_16 : _GEN_686; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_688 = 14'h11 == parameter_2_14 ? phv_data_17 : _GEN_687; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_689 = 14'h12 == parameter_2_14 ? phv_data_18 : _GEN_688; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_690 = 14'h13 == parameter_2_14 ? phv_data_19 : _GEN_689; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_691 = 14'h14 == parameter_2_14 ? phv_data_20 : _GEN_690; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_692 = 14'h15 == parameter_2_14 ? phv_data_21 : _GEN_691; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_693 = 14'h16 == parameter_2_14 ? phv_data_22 : _GEN_692; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_694 = 14'h17 == parameter_2_14 ? phv_data_23 : _GEN_693; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_695 = 14'h18 == parameter_2_14 ? phv_data_24 : _GEN_694; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_696 = 14'h19 == parameter_2_14 ? phv_data_25 : _GEN_695; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_697 = 14'h1a == parameter_2_14 ? phv_data_26 : _GEN_696; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_698 = 14'h1b == parameter_2_14 ? phv_data_27 : _GEN_697; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_699 = 14'h1c == parameter_2_14 ? phv_data_28 : _GEN_698; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_700 = 14'h1d == parameter_2_14 ? phv_data_29 : _GEN_699; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_701 = 14'h1e == parameter_2_14 ? phv_data_30 : _GEN_700; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_702 = 14'h1f == parameter_2_14 ? phv_data_31 : _GEN_701; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_15 = vliw_15[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_15 = vliw_15[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_15 = parameter_2_15[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_15 = parameter_2_15[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_15 = {{1'd0}, args_offset_15}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_15 = _total_offset_T_15[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_706 = 3'h1 == total_offset_15 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_707 = 3'h2 == total_offset_15 ? args_2 : _GEN_706; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_708 = 3'h3 == total_offset_15 ? args_3 : _GEN_707; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_709 = 3'h4 == total_offset_15 ? args_4 : _GEN_708; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_710 = 3'h5 == total_offset_15 ? args_5 : _GEN_709; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_711 = 3'h6 == total_offset_15 ? args_6 : _GEN_710; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_712 = total_offset_15 < 3'h7 ? _GEN_711 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_15_0 = 3'h0 < args_length_15 ? _GEN_712 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_714 = opcode_15 == 4'ha ? field_bytes_15_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_715 = opcode_15 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_588 = opcode_15 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_31 = _T_588 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_716 = opcode_15 == 4'h8 | opcode_15 == 4'hb ? parameter_2_15[7:0] : _GEN_714; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_717 = opcode_15 == 4'h8 | opcode_15 == 4'hb ? _field_tag_T_31 : _GEN_715; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_718 = 14'h0 == parameter_2_15 ? phv_data_0 : _GEN_716; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_719 = 14'h1 == parameter_2_15 ? phv_data_1 : _GEN_718; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_720 = 14'h2 == parameter_2_15 ? phv_data_2 : _GEN_719; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_721 = 14'h3 == parameter_2_15 ? phv_data_3 : _GEN_720; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_722 = 14'h4 == parameter_2_15 ? phv_data_4 : _GEN_721; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_723 = 14'h5 == parameter_2_15 ? phv_data_5 : _GEN_722; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_724 = 14'h6 == parameter_2_15 ? phv_data_6 : _GEN_723; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_725 = 14'h7 == parameter_2_15 ? phv_data_7 : _GEN_724; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_726 = 14'h8 == parameter_2_15 ? phv_data_8 : _GEN_725; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_727 = 14'h9 == parameter_2_15 ? phv_data_9 : _GEN_726; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_728 = 14'ha == parameter_2_15 ? phv_data_10 : _GEN_727; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_729 = 14'hb == parameter_2_15 ? phv_data_11 : _GEN_728; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_730 = 14'hc == parameter_2_15 ? phv_data_12 : _GEN_729; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_731 = 14'hd == parameter_2_15 ? phv_data_13 : _GEN_730; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_732 = 14'he == parameter_2_15 ? phv_data_14 : _GEN_731; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_733 = 14'hf == parameter_2_15 ? phv_data_15 : _GEN_732; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_734 = 14'h10 == parameter_2_15 ? phv_data_16 : _GEN_733; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_735 = 14'h11 == parameter_2_15 ? phv_data_17 : _GEN_734; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_736 = 14'h12 == parameter_2_15 ? phv_data_18 : _GEN_735; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_737 = 14'h13 == parameter_2_15 ? phv_data_19 : _GEN_736; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_738 = 14'h14 == parameter_2_15 ? phv_data_20 : _GEN_737; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_739 = 14'h15 == parameter_2_15 ? phv_data_21 : _GEN_738; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_740 = 14'h16 == parameter_2_15 ? phv_data_22 : _GEN_739; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_741 = 14'h17 == parameter_2_15 ? phv_data_23 : _GEN_740; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_742 = 14'h18 == parameter_2_15 ? phv_data_24 : _GEN_741; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_743 = 14'h19 == parameter_2_15 ? phv_data_25 : _GEN_742; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_744 = 14'h1a == parameter_2_15 ? phv_data_26 : _GEN_743; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_745 = 14'h1b == parameter_2_15 ? phv_data_27 : _GEN_744; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_746 = 14'h1c == parameter_2_15 ? phv_data_28 : _GEN_745; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_747 = 14'h1d == parameter_2_15 ? phv_data_29 : _GEN_746; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_748 = 14'h1e == parameter_2_15 ? phv_data_30 : _GEN_747; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_749 = 14'h1f == parameter_2_15 ? phv_data_31 : _GEN_748; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_16 = vliw_16[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_16 = vliw_16[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_16 = parameter_2_16[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_16 = parameter_2_16[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_16 = {{1'd0}, args_offset_16}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_16 = _total_offset_T_16[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_753 = 3'h1 == total_offset_16 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_754 = 3'h2 == total_offset_16 ? args_2 : _GEN_753; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_755 = 3'h3 == total_offset_16 ? args_3 : _GEN_754; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_756 = 3'h4 == total_offset_16 ? args_4 : _GEN_755; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_757 = 3'h5 == total_offset_16 ? args_5 : _GEN_756; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_758 = 3'h6 == total_offset_16 ? args_6 : _GEN_757; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_759 = total_offset_16 < 3'h7 ? _GEN_758 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_16_0 = 3'h0 < args_length_16 ? _GEN_759 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_761 = opcode_16 == 4'ha ? field_bytes_16_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_762 = opcode_16 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_627 = opcode_16 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_33 = _T_627 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_763 = opcode_16 == 4'h8 | opcode_16 == 4'hb ? parameter_2_16[7:0] : _GEN_761; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_764 = opcode_16 == 4'h8 | opcode_16 == 4'hb ? _field_tag_T_33 : _GEN_762; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_765 = 14'h0 == parameter_2_16 ? phv_data_0 : _GEN_763; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_766 = 14'h1 == parameter_2_16 ? phv_data_1 : _GEN_765; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_767 = 14'h2 == parameter_2_16 ? phv_data_2 : _GEN_766; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_768 = 14'h3 == parameter_2_16 ? phv_data_3 : _GEN_767; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_769 = 14'h4 == parameter_2_16 ? phv_data_4 : _GEN_768; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_770 = 14'h5 == parameter_2_16 ? phv_data_5 : _GEN_769; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_771 = 14'h6 == parameter_2_16 ? phv_data_6 : _GEN_770; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_772 = 14'h7 == parameter_2_16 ? phv_data_7 : _GEN_771; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_773 = 14'h8 == parameter_2_16 ? phv_data_8 : _GEN_772; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_774 = 14'h9 == parameter_2_16 ? phv_data_9 : _GEN_773; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_775 = 14'ha == parameter_2_16 ? phv_data_10 : _GEN_774; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_776 = 14'hb == parameter_2_16 ? phv_data_11 : _GEN_775; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_777 = 14'hc == parameter_2_16 ? phv_data_12 : _GEN_776; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_778 = 14'hd == parameter_2_16 ? phv_data_13 : _GEN_777; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_779 = 14'he == parameter_2_16 ? phv_data_14 : _GEN_778; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_780 = 14'hf == parameter_2_16 ? phv_data_15 : _GEN_779; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_781 = 14'h10 == parameter_2_16 ? phv_data_16 : _GEN_780; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_782 = 14'h11 == parameter_2_16 ? phv_data_17 : _GEN_781; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_783 = 14'h12 == parameter_2_16 ? phv_data_18 : _GEN_782; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_784 = 14'h13 == parameter_2_16 ? phv_data_19 : _GEN_783; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_785 = 14'h14 == parameter_2_16 ? phv_data_20 : _GEN_784; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_786 = 14'h15 == parameter_2_16 ? phv_data_21 : _GEN_785; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_787 = 14'h16 == parameter_2_16 ? phv_data_22 : _GEN_786; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_788 = 14'h17 == parameter_2_16 ? phv_data_23 : _GEN_787; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_789 = 14'h18 == parameter_2_16 ? phv_data_24 : _GEN_788; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_790 = 14'h19 == parameter_2_16 ? phv_data_25 : _GEN_789; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_791 = 14'h1a == parameter_2_16 ? phv_data_26 : _GEN_790; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_792 = 14'h1b == parameter_2_16 ? phv_data_27 : _GEN_791; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_793 = 14'h1c == parameter_2_16 ? phv_data_28 : _GEN_792; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_794 = 14'h1d == parameter_2_16 ? phv_data_29 : _GEN_793; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_795 = 14'h1e == parameter_2_16 ? phv_data_30 : _GEN_794; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_796 = 14'h1f == parameter_2_16 ? phv_data_31 : _GEN_795; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_17 = vliw_17[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_17 = vliw_17[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_17 = parameter_2_17[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_17 = parameter_2_17[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_17 = {{1'd0}, args_offset_17}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_17 = _total_offset_T_17[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_800 = 3'h1 == total_offset_17 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_801 = 3'h2 == total_offset_17 ? args_2 : _GEN_800; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_802 = 3'h3 == total_offset_17 ? args_3 : _GEN_801; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_803 = 3'h4 == total_offset_17 ? args_4 : _GEN_802; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_804 = 3'h5 == total_offset_17 ? args_5 : _GEN_803; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_805 = 3'h6 == total_offset_17 ? args_6 : _GEN_804; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_806 = total_offset_17 < 3'h7 ? _GEN_805 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_17_0 = 3'h0 < args_length_17 ? _GEN_806 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_808 = opcode_17 == 4'ha ? field_bytes_17_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_809 = opcode_17 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_666 = opcode_17 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_35 = _T_666 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_810 = opcode_17 == 4'h8 | opcode_17 == 4'hb ? parameter_2_17[7:0] : _GEN_808; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_811 = opcode_17 == 4'h8 | opcode_17 == 4'hb ? _field_tag_T_35 : _GEN_809; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_812 = 14'h0 == parameter_2_17 ? phv_data_0 : _GEN_810; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_813 = 14'h1 == parameter_2_17 ? phv_data_1 : _GEN_812; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_814 = 14'h2 == parameter_2_17 ? phv_data_2 : _GEN_813; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_815 = 14'h3 == parameter_2_17 ? phv_data_3 : _GEN_814; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_816 = 14'h4 == parameter_2_17 ? phv_data_4 : _GEN_815; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_817 = 14'h5 == parameter_2_17 ? phv_data_5 : _GEN_816; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_818 = 14'h6 == parameter_2_17 ? phv_data_6 : _GEN_817; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_819 = 14'h7 == parameter_2_17 ? phv_data_7 : _GEN_818; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_820 = 14'h8 == parameter_2_17 ? phv_data_8 : _GEN_819; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_821 = 14'h9 == parameter_2_17 ? phv_data_9 : _GEN_820; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_822 = 14'ha == parameter_2_17 ? phv_data_10 : _GEN_821; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_823 = 14'hb == parameter_2_17 ? phv_data_11 : _GEN_822; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_824 = 14'hc == parameter_2_17 ? phv_data_12 : _GEN_823; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_825 = 14'hd == parameter_2_17 ? phv_data_13 : _GEN_824; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_826 = 14'he == parameter_2_17 ? phv_data_14 : _GEN_825; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_827 = 14'hf == parameter_2_17 ? phv_data_15 : _GEN_826; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_828 = 14'h10 == parameter_2_17 ? phv_data_16 : _GEN_827; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_829 = 14'h11 == parameter_2_17 ? phv_data_17 : _GEN_828; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_830 = 14'h12 == parameter_2_17 ? phv_data_18 : _GEN_829; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_831 = 14'h13 == parameter_2_17 ? phv_data_19 : _GEN_830; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_832 = 14'h14 == parameter_2_17 ? phv_data_20 : _GEN_831; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_833 = 14'h15 == parameter_2_17 ? phv_data_21 : _GEN_832; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_834 = 14'h16 == parameter_2_17 ? phv_data_22 : _GEN_833; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_835 = 14'h17 == parameter_2_17 ? phv_data_23 : _GEN_834; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_836 = 14'h18 == parameter_2_17 ? phv_data_24 : _GEN_835; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_837 = 14'h19 == parameter_2_17 ? phv_data_25 : _GEN_836; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_838 = 14'h1a == parameter_2_17 ? phv_data_26 : _GEN_837; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_839 = 14'h1b == parameter_2_17 ? phv_data_27 : _GEN_838; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_840 = 14'h1c == parameter_2_17 ? phv_data_28 : _GEN_839; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_841 = 14'h1d == parameter_2_17 ? phv_data_29 : _GEN_840; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_842 = 14'h1e == parameter_2_17 ? phv_data_30 : _GEN_841; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_843 = 14'h1f == parameter_2_17 ? phv_data_31 : _GEN_842; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_18 = vliw_18[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_18 = vliw_18[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_18 = parameter_2_18[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_18 = parameter_2_18[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_18 = {{1'd0}, args_offset_18}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_18 = _total_offset_T_18[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_847 = 3'h1 == total_offset_18 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_848 = 3'h2 == total_offset_18 ? args_2 : _GEN_847; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_849 = 3'h3 == total_offset_18 ? args_3 : _GEN_848; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_850 = 3'h4 == total_offset_18 ? args_4 : _GEN_849; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_851 = 3'h5 == total_offset_18 ? args_5 : _GEN_850; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_852 = 3'h6 == total_offset_18 ? args_6 : _GEN_851; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_853 = total_offset_18 < 3'h7 ? _GEN_852 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_18_0 = 3'h0 < args_length_18 ? _GEN_853 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_855 = opcode_18 == 4'ha ? field_bytes_18_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_856 = opcode_18 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_705 = opcode_18 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_37 = _T_705 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_857 = opcode_18 == 4'h8 | opcode_18 == 4'hb ? parameter_2_18[7:0] : _GEN_855; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_858 = opcode_18 == 4'h8 | opcode_18 == 4'hb ? _field_tag_T_37 : _GEN_856; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_859 = 14'h0 == parameter_2_18 ? phv_data_0 : _GEN_857; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_860 = 14'h1 == parameter_2_18 ? phv_data_1 : _GEN_859; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_861 = 14'h2 == parameter_2_18 ? phv_data_2 : _GEN_860; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_862 = 14'h3 == parameter_2_18 ? phv_data_3 : _GEN_861; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_863 = 14'h4 == parameter_2_18 ? phv_data_4 : _GEN_862; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_864 = 14'h5 == parameter_2_18 ? phv_data_5 : _GEN_863; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_865 = 14'h6 == parameter_2_18 ? phv_data_6 : _GEN_864; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_866 = 14'h7 == parameter_2_18 ? phv_data_7 : _GEN_865; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_867 = 14'h8 == parameter_2_18 ? phv_data_8 : _GEN_866; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_868 = 14'h9 == parameter_2_18 ? phv_data_9 : _GEN_867; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_869 = 14'ha == parameter_2_18 ? phv_data_10 : _GEN_868; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_870 = 14'hb == parameter_2_18 ? phv_data_11 : _GEN_869; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_871 = 14'hc == parameter_2_18 ? phv_data_12 : _GEN_870; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_872 = 14'hd == parameter_2_18 ? phv_data_13 : _GEN_871; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_873 = 14'he == parameter_2_18 ? phv_data_14 : _GEN_872; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_874 = 14'hf == parameter_2_18 ? phv_data_15 : _GEN_873; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_875 = 14'h10 == parameter_2_18 ? phv_data_16 : _GEN_874; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_876 = 14'h11 == parameter_2_18 ? phv_data_17 : _GEN_875; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_877 = 14'h12 == parameter_2_18 ? phv_data_18 : _GEN_876; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_878 = 14'h13 == parameter_2_18 ? phv_data_19 : _GEN_877; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_879 = 14'h14 == parameter_2_18 ? phv_data_20 : _GEN_878; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_880 = 14'h15 == parameter_2_18 ? phv_data_21 : _GEN_879; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_881 = 14'h16 == parameter_2_18 ? phv_data_22 : _GEN_880; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_882 = 14'h17 == parameter_2_18 ? phv_data_23 : _GEN_881; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_883 = 14'h18 == parameter_2_18 ? phv_data_24 : _GEN_882; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_884 = 14'h19 == parameter_2_18 ? phv_data_25 : _GEN_883; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_885 = 14'h1a == parameter_2_18 ? phv_data_26 : _GEN_884; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_886 = 14'h1b == parameter_2_18 ? phv_data_27 : _GEN_885; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_887 = 14'h1c == parameter_2_18 ? phv_data_28 : _GEN_886; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_888 = 14'h1d == parameter_2_18 ? phv_data_29 : _GEN_887; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_889 = 14'h1e == parameter_2_18 ? phv_data_30 : _GEN_888; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_890 = 14'h1f == parameter_2_18 ? phv_data_31 : _GEN_889; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_19 = vliw_19[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_19 = vliw_19[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_19 = parameter_2_19[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_19 = parameter_2_19[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_19 = {{1'd0}, args_offset_19}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_19 = _total_offset_T_19[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_894 = 3'h1 == total_offset_19 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_895 = 3'h2 == total_offset_19 ? args_2 : _GEN_894; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_896 = 3'h3 == total_offset_19 ? args_3 : _GEN_895; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_897 = 3'h4 == total_offset_19 ? args_4 : _GEN_896; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_898 = 3'h5 == total_offset_19 ? args_5 : _GEN_897; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_899 = 3'h6 == total_offset_19 ? args_6 : _GEN_898; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_900 = total_offset_19 < 3'h7 ? _GEN_899 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_19_0 = 3'h0 < args_length_19 ? _GEN_900 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_902 = opcode_19 == 4'ha ? field_bytes_19_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_903 = opcode_19 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_744 = opcode_19 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_39 = _T_744 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_904 = opcode_19 == 4'h8 | opcode_19 == 4'hb ? parameter_2_19[7:0] : _GEN_902; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_905 = opcode_19 == 4'h8 | opcode_19 == 4'hb ? _field_tag_T_39 : _GEN_903; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_906 = 14'h0 == parameter_2_19 ? phv_data_0 : _GEN_904; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_907 = 14'h1 == parameter_2_19 ? phv_data_1 : _GEN_906; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_908 = 14'h2 == parameter_2_19 ? phv_data_2 : _GEN_907; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_909 = 14'h3 == parameter_2_19 ? phv_data_3 : _GEN_908; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_910 = 14'h4 == parameter_2_19 ? phv_data_4 : _GEN_909; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_911 = 14'h5 == parameter_2_19 ? phv_data_5 : _GEN_910; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_912 = 14'h6 == parameter_2_19 ? phv_data_6 : _GEN_911; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_913 = 14'h7 == parameter_2_19 ? phv_data_7 : _GEN_912; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_914 = 14'h8 == parameter_2_19 ? phv_data_8 : _GEN_913; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_915 = 14'h9 == parameter_2_19 ? phv_data_9 : _GEN_914; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_916 = 14'ha == parameter_2_19 ? phv_data_10 : _GEN_915; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_917 = 14'hb == parameter_2_19 ? phv_data_11 : _GEN_916; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_918 = 14'hc == parameter_2_19 ? phv_data_12 : _GEN_917; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_919 = 14'hd == parameter_2_19 ? phv_data_13 : _GEN_918; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_920 = 14'he == parameter_2_19 ? phv_data_14 : _GEN_919; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_921 = 14'hf == parameter_2_19 ? phv_data_15 : _GEN_920; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_922 = 14'h10 == parameter_2_19 ? phv_data_16 : _GEN_921; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_923 = 14'h11 == parameter_2_19 ? phv_data_17 : _GEN_922; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_924 = 14'h12 == parameter_2_19 ? phv_data_18 : _GEN_923; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_925 = 14'h13 == parameter_2_19 ? phv_data_19 : _GEN_924; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_926 = 14'h14 == parameter_2_19 ? phv_data_20 : _GEN_925; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_927 = 14'h15 == parameter_2_19 ? phv_data_21 : _GEN_926; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_928 = 14'h16 == parameter_2_19 ? phv_data_22 : _GEN_927; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_929 = 14'h17 == parameter_2_19 ? phv_data_23 : _GEN_928; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_930 = 14'h18 == parameter_2_19 ? phv_data_24 : _GEN_929; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_931 = 14'h19 == parameter_2_19 ? phv_data_25 : _GEN_930; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_932 = 14'h1a == parameter_2_19 ? phv_data_26 : _GEN_931; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_933 = 14'h1b == parameter_2_19 ? phv_data_27 : _GEN_932; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_934 = 14'h1c == parameter_2_19 ? phv_data_28 : _GEN_933; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_935 = 14'h1d == parameter_2_19 ? phv_data_29 : _GEN_934; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_936 = 14'h1e == parameter_2_19 ? phv_data_30 : _GEN_935; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_937 = 14'h1f == parameter_2_19 ? phv_data_31 : _GEN_936; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_20 = vliw_20[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_20 = vliw_20[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_20 = parameter_2_20[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_20 = parameter_2_20[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_20 = {{1'd0}, args_offset_20}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_20 = _total_offset_T_20[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_941 = 3'h1 == total_offset_20 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_942 = 3'h2 == total_offset_20 ? args_2 : _GEN_941; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_943 = 3'h3 == total_offset_20 ? args_3 : _GEN_942; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_944 = 3'h4 == total_offset_20 ? args_4 : _GEN_943; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_945 = 3'h5 == total_offset_20 ? args_5 : _GEN_944; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_946 = 3'h6 == total_offset_20 ? args_6 : _GEN_945; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_947 = total_offset_20 < 3'h7 ? _GEN_946 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_20_0 = 3'h0 < args_length_20 ? _GEN_947 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_949 = opcode_20 == 4'ha ? field_bytes_20_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_950 = opcode_20 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_783 = opcode_20 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_41 = _T_783 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_951 = opcode_20 == 4'h8 | opcode_20 == 4'hb ? parameter_2_20[7:0] : _GEN_949; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_952 = opcode_20 == 4'h8 | opcode_20 == 4'hb ? _field_tag_T_41 : _GEN_950; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_953 = 14'h0 == parameter_2_20 ? phv_data_0 : _GEN_951; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_954 = 14'h1 == parameter_2_20 ? phv_data_1 : _GEN_953; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_955 = 14'h2 == parameter_2_20 ? phv_data_2 : _GEN_954; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_956 = 14'h3 == parameter_2_20 ? phv_data_3 : _GEN_955; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_957 = 14'h4 == parameter_2_20 ? phv_data_4 : _GEN_956; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_958 = 14'h5 == parameter_2_20 ? phv_data_5 : _GEN_957; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_959 = 14'h6 == parameter_2_20 ? phv_data_6 : _GEN_958; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_960 = 14'h7 == parameter_2_20 ? phv_data_7 : _GEN_959; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_961 = 14'h8 == parameter_2_20 ? phv_data_8 : _GEN_960; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_962 = 14'h9 == parameter_2_20 ? phv_data_9 : _GEN_961; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_963 = 14'ha == parameter_2_20 ? phv_data_10 : _GEN_962; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_964 = 14'hb == parameter_2_20 ? phv_data_11 : _GEN_963; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_965 = 14'hc == parameter_2_20 ? phv_data_12 : _GEN_964; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_966 = 14'hd == parameter_2_20 ? phv_data_13 : _GEN_965; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_967 = 14'he == parameter_2_20 ? phv_data_14 : _GEN_966; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_968 = 14'hf == parameter_2_20 ? phv_data_15 : _GEN_967; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_969 = 14'h10 == parameter_2_20 ? phv_data_16 : _GEN_968; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_970 = 14'h11 == parameter_2_20 ? phv_data_17 : _GEN_969; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_971 = 14'h12 == parameter_2_20 ? phv_data_18 : _GEN_970; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_972 = 14'h13 == parameter_2_20 ? phv_data_19 : _GEN_971; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_973 = 14'h14 == parameter_2_20 ? phv_data_20 : _GEN_972; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_974 = 14'h15 == parameter_2_20 ? phv_data_21 : _GEN_973; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_975 = 14'h16 == parameter_2_20 ? phv_data_22 : _GEN_974; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_976 = 14'h17 == parameter_2_20 ? phv_data_23 : _GEN_975; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_977 = 14'h18 == parameter_2_20 ? phv_data_24 : _GEN_976; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_978 = 14'h19 == parameter_2_20 ? phv_data_25 : _GEN_977; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_979 = 14'h1a == parameter_2_20 ? phv_data_26 : _GEN_978; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_980 = 14'h1b == parameter_2_20 ? phv_data_27 : _GEN_979; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_981 = 14'h1c == parameter_2_20 ? phv_data_28 : _GEN_980; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_982 = 14'h1d == parameter_2_20 ? phv_data_29 : _GEN_981; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_983 = 14'h1e == parameter_2_20 ? phv_data_30 : _GEN_982; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_984 = 14'h1f == parameter_2_20 ? phv_data_31 : _GEN_983; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_21 = vliw_21[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_21 = vliw_21[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_21 = parameter_2_21[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_21 = parameter_2_21[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_21 = {{1'd0}, args_offset_21}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_21 = _total_offset_T_21[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_988 = 3'h1 == total_offset_21 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_989 = 3'h2 == total_offset_21 ? args_2 : _GEN_988; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_990 = 3'h3 == total_offset_21 ? args_3 : _GEN_989; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_991 = 3'h4 == total_offset_21 ? args_4 : _GEN_990; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_992 = 3'h5 == total_offset_21 ? args_5 : _GEN_991; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_993 = 3'h6 == total_offset_21 ? args_6 : _GEN_992; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_994 = total_offset_21 < 3'h7 ? _GEN_993 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_21_0 = 3'h0 < args_length_21 ? _GEN_994 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_996 = opcode_21 == 4'ha ? field_bytes_21_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_997 = opcode_21 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_822 = opcode_21 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_43 = _T_822 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_998 = opcode_21 == 4'h8 | opcode_21 == 4'hb ? parameter_2_21[7:0] : _GEN_996; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_999 = opcode_21 == 4'h8 | opcode_21 == 4'hb ? _field_tag_T_43 : _GEN_997; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1000 = 14'h0 == parameter_2_21 ? phv_data_0 : _GEN_998; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1001 = 14'h1 == parameter_2_21 ? phv_data_1 : _GEN_1000; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1002 = 14'h2 == parameter_2_21 ? phv_data_2 : _GEN_1001; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1003 = 14'h3 == parameter_2_21 ? phv_data_3 : _GEN_1002; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1004 = 14'h4 == parameter_2_21 ? phv_data_4 : _GEN_1003; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1005 = 14'h5 == parameter_2_21 ? phv_data_5 : _GEN_1004; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1006 = 14'h6 == parameter_2_21 ? phv_data_6 : _GEN_1005; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1007 = 14'h7 == parameter_2_21 ? phv_data_7 : _GEN_1006; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1008 = 14'h8 == parameter_2_21 ? phv_data_8 : _GEN_1007; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1009 = 14'h9 == parameter_2_21 ? phv_data_9 : _GEN_1008; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1010 = 14'ha == parameter_2_21 ? phv_data_10 : _GEN_1009; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1011 = 14'hb == parameter_2_21 ? phv_data_11 : _GEN_1010; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1012 = 14'hc == parameter_2_21 ? phv_data_12 : _GEN_1011; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1013 = 14'hd == parameter_2_21 ? phv_data_13 : _GEN_1012; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1014 = 14'he == parameter_2_21 ? phv_data_14 : _GEN_1013; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1015 = 14'hf == parameter_2_21 ? phv_data_15 : _GEN_1014; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1016 = 14'h10 == parameter_2_21 ? phv_data_16 : _GEN_1015; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1017 = 14'h11 == parameter_2_21 ? phv_data_17 : _GEN_1016; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1018 = 14'h12 == parameter_2_21 ? phv_data_18 : _GEN_1017; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1019 = 14'h13 == parameter_2_21 ? phv_data_19 : _GEN_1018; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1020 = 14'h14 == parameter_2_21 ? phv_data_20 : _GEN_1019; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1021 = 14'h15 == parameter_2_21 ? phv_data_21 : _GEN_1020; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1022 = 14'h16 == parameter_2_21 ? phv_data_22 : _GEN_1021; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1023 = 14'h17 == parameter_2_21 ? phv_data_23 : _GEN_1022; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1024 = 14'h18 == parameter_2_21 ? phv_data_24 : _GEN_1023; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1025 = 14'h19 == parameter_2_21 ? phv_data_25 : _GEN_1024; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1026 = 14'h1a == parameter_2_21 ? phv_data_26 : _GEN_1025; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1027 = 14'h1b == parameter_2_21 ? phv_data_27 : _GEN_1026; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1028 = 14'h1c == parameter_2_21 ? phv_data_28 : _GEN_1027; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1029 = 14'h1d == parameter_2_21 ? phv_data_29 : _GEN_1028; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1030 = 14'h1e == parameter_2_21 ? phv_data_30 : _GEN_1029; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1031 = 14'h1f == parameter_2_21 ? phv_data_31 : _GEN_1030; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_22 = vliw_22[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_22 = vliw_22[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_22 = parameter_2_22[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_22 = parameter_2_22[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_22 = {{1'd0}, args_offset_22}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_22 = _total_offset_T_22[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1035 = 3'h1 == total_offset_22 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1036 = 3'h2 == total_offset_22 ? args_2 : _GEN_1035; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1037 = 3'h3 == total_offset_22 ? args_3 : _GEN_1036; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1038 = 3'h4 == total_offset_22 ? args_4 : _GEN_1037; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1039 = 3'h5 == total_offset_22 ? args_5 : _GEN_1038; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1040 = 3'h6 == total_offset_22 ? args_6 : _GEN_1039; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1041 = total_offset_22 < 3'h7 ? _GEN_1040 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_22_0 = 3'h0 < args_length_22 ? _GEN_1041 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1043 = opcode_22 == 4'ha ? field_bytes_22_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1044 = opcode_22 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_861 = opcode_22 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_45 = _T_861 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1045 = opcode_22 == 4'h8 | opcode_22 == 4'hb ? parameter_2_22[7:0] : _GEN_1043; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1046 = opcode_22 == 4'h8 | opcode_22 == 4'hb ? _field_tag_T_45 : _GEN_1044; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1047 = 14'h0 == parameter_2_22 ? phv_data_0 : _GEN_1045; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1048 = 14'h1 == parameter_2_22 ? phv_data_1 : _GEN_1047; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1049 = 14'h2 == parameter_2_22 ? phv_data_2 : _GEN_1048; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1050 = 14'h3 == parameter_2_22 ? phv_data_3 : _GEN_1049; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1051 = 14'h4 == parameter_2_22 ? phv_data_4 : _GEN_1050; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1052 = 14'h5 == parameter_2_22 ? phv_data_5 : _GEN_1051; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1053 = 14'h6 == parameter_2_22 ? phv_data_6 : _GEN_1052; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1054 = 14'h7 == parameter_2_22 ? phv_data_7 : _GEN_1053; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1055 = 14'h8 == parameter_2_22 ? phv_data_8 : _GEN_1054; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1056 = 14'h9 == parameter_2_22 ? phv_data_9 : _GEN_1055; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1057 = 14'ha == parameter_2_22 ? phv_data_10 : _GEN_1056; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1058 = 14'hb == parameter_2_22 ? phv_data_11 : _GEN_1057; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1059 = 14'hc == parameter_2_22 ? phv_data_12 : _GEN_1058; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1060 = 14'hd == parameter_2_22 ? phv_data_13 : _GEN_1059; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1061 = 14'he == parameter_2_22 ? phv_data_14 : _GEN_1060; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1062 = 14'hf == parameter_2_22 ? phv_data_15 : _GEN_1061; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1063 = 14'h10 == parameter_2_22 ? phv_data_16 : _GEN_1062; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1064 = 14'h11 == parameter_2_22 ? phv_data_17 : _GEN_1063; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1065 = 14'h12 == parameter_2_22 ? phv_data_18 : _GEN_1064; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1066 = 14'h13 == parameter_2_22 ? phv_data_19 : _GEN_1065; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1067 = 14'h14 == parameter_2_22 ? phv_data_20 : _GEN_1066; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1068 = 14'h15 == parameter_2_22 ? phv_data_21 : _GEN_1067; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1069 = 14'h16 == parameter_2_22 ? phv_data_22 : _GEN_1068; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1070 = 14'h17 == parameter_2_22 ? phv_data_23 : _GEN_1069; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1071 = 14'h18 == parameter_2_22 ? phv_data_24 : _GEN_1070; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1072 = 14'h19 == parameter_2_22 ? phv_data_25 : _GEN_1071; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1073 = 14'h1a == parameter_2_22 ? phv_data_26 : _GEN_1072; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1074 = 14'h1b == parameter_2_22 ? phv_data_27 : _GEN_1073; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1075 = 14'h1c == parameter_2_22 ? phv_data_28 : _GEN_1074; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1076 = 14'h1d == parameter_2_22 ? phv_data_29 : _GEN_1075; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1077 = 14'h1e == parameter_2_22 ? phv_data_30 : _GEN_1076; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1078 = 14'h1f == parameter_2_22 ? phv_data_31 : _GEN_1077; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_23 = vliw_23[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_23 = vliw_23[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_23 = parameter_2_23[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_23 = parameter_2_23[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_23 = {{1'd0}, args_offset_23}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_23 = _total_offset_T_23[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1082 = 3'h1 == total_offset_23 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1083 = 3'h2 == total_offset_23 ? args_2 : _GEN_1082; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1084 = 3'h3 == total_offset_23 ? args_3 : _GEN_1083; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1085 = 3'h4 == total_offset_23 ? args_4 : _GEN_1084; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1086 = 3'h5 == total_offset_23 ? args_5 : _GEN_1085; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1087 = 3'h6 == total_offset_23 ? args_6 : _GEN_1086; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1088 = total_offset_23 < 3'h7 ? _GEN_1087 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_23_0 = 3'h0 < args_length_23 ? _GEN_1088 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1090 = opcode_23 == 4'ha ? field_bytes_23_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1091 = opcode_23 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_900 = opcode_23 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_47 = _T_900 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1092 = opcode_23 == 4'h8 | opcode_23 == 4'hb ? parameter_2_23[7:0] : _GEN_1090; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1093 = opcode_23 == 4'h8 | opcode_23 == 4'hb ? _field_tag_T_47 : _GEN_1091; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1094 = 14'h0 == parameter_2_23 ? phv_data_0 : _GEN_1092; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1095 = 14'h1 == parameter_2_23 ? phv_data_1 : _GEN_1094; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1096 = 14'h2 == parameter_2_23 ? phv_data_2 : _GEN_1095; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1097 = 14'h3 == parameter_2_23 ? phv_data_3 : _GEN_1096; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1098 = 14'h4 == parameter_2_23 ? phv_data_4 : _GEN_1097; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1099 = 14'h5 == parameter_2_23 ? phv_data_5 : _GEN_1098; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1100 = 14'h6 == parameter_2_23 ? phv_data_6 : _GEN_1099; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1101 = 14'h7 == parameter_2_23 ? phv_data_7 : _GEN_1100; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1102 = 14'h8 == parameter_2_23 ? phv_data_8 : _GEN_1101; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1103 = 14'h9 == parameter_2_23 ? phv_data_9 : _GEN_1102; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1104 = 14'ha == parameter_2_23 ? phv_data_10 : _GEN_1103; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1105 = 14'hb == parameter_2_23 ? phv_data_11 : _GEN_1104; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1106 = 14'hc == parameter_2_23 ? phv_data_12 : _GEN_1105; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1107 = 14'hd == parameter_2_23 ? phv_data_13 : _GEN_1106; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1108 = 14'he == parameter_2_23 ? phv_data_14 : _GEN_1107; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1109 = 14'hf == parameter_2_23 ? phv_data_15 : _GEN_1108; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1110 = 14'h10 == parameter_2_23 ? phv_data_16 : _GEN_1109; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1111 = 14'h11 == parameter_2_23 ? phv_data_17 : _GEN_1110; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1112 = 14'h12 == parameter_2_23 ? phv_data_18 : _GEN_1111; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1113 = 14'h13 == parameter_2_23 ? phv_data_19 : _GEN_1112; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1114 = 14'h14 == parameter_2_23 ? phv_data_20 : _GEN_1113; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1115 = 14'h15 == parameter_2_23 ? phv_data_21 : _GEN_1114; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1116 = 14'h16 == parameter_2_23 ? phv_data_22 : _GEN_1115; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1117 = 14'h17 == parameter_2_23 ? phv_data_23 : _GEN_1116; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1118 = 14'h18 == parameter_2_23 ? phv_data_24 : _GEN_1117; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1119 = 14'h19 == parameter_2_23 ? phv_data_25 : _GEN_1118; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1120 = 14'h1a == parameter_2_23 ? phv_data_26 : _GEN_1119; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1121 = 14'h1b == parameter_2_23 ? phv_data_27 : _GEN_1120; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1122 = 14'h1c == parameter_2_23 ? phv_data_28 : _GEN_1121; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1123 = 14'h1d == parameter_2_23 ? phv_data_29 : _GEN_1122; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1124 = 14'h1e == parameter_2_23 ? phv_data_30 : _GEN_1123; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1125 = 14'h1f == parameter_2_23 ? phv_data_31 : _GEN_1124; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_24 = vliw_24[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_24 = vliw_24[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_24 = parameter_2_24[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_24 = parameter_2_24[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_24 = {{1'd0}, args_offset_24}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_24 = _total_offset_T_24[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1129 = 3'h1 == total_offset_24 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1130 = 3'h2 == total_offset_24 ? args_2 : _GEN_1129; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1131 = 3'h3 == total_offset_24 ? args_3 : _GEN_1130; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1132 = 3'h4 == total_offset_24 ? args_4 : _GEN_1131; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1133 = 3'h5 == total_offset_24 ? args_5 : _GEN_1132; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1134 = 3'h6 == total_offset_24 ? args_6 : _GEN_1133; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1135 = total_offset_24 < 3'h7 ? _GEN_1134 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_24_0 = 3'h0 < args_length_24 ? _GEN_1135 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1137 = opcode_24 == 4'ha ? field_bytes_24_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1138 = opcode_24 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_939 = opcode_24 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_49 = _T_939 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1139 = opcode_24 == 4'h8 | opcode_24 == 4'hb ? parameter_2_24[7:0] : _GEN_1137; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1140 = opcode_24 == 4'h8 | opcode_24 == 4'hb ? _field_tag_T_49 : _GEN_1138; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1141 = 14'h0 == parameter_2_24 ? phv_data_0 : _GEN_1139; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1142 = 14'h1 == parameter_2_24 ? phv_data_1 : _GEN_1141; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1143 = 14'h2 == parameter_2_24 ? phv_data_2 : _GEN_1142; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1144 = 14'h3 == parameter_2_24 ? phv_data_3 : _GEN_1143; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1145 = 14'h4 == parameter_2_24 ? phv_data_4 : _GEN_1144; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1146 = 14'h5 == parameter_2_24 ? phv_data_5 : _GEN_1145; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1147 = 14'h6 == parameter_2_24 ? phv_data_6 : _GEN_1146; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1148 = 14'h7 == parameter_2_24 ? phv_data_7 : _GEN_1147; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1149 = 14'h8 == parameter_2_24 ? phv_data_8 : _GEN_1148; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1150 = 14'h9 == parameter_2_24 ? phv_data_9 : _GEN_1149; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1151 = 14'ha == parameter_2_24 ? phv_data_10 : _GEN_1150; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1152 = 14'hb == parameter_2_24 ? phv_data_11 : _GEN_1151; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1153 = 14'hc == parameter_2_24 ? phv_data_12 : _GEN_1152; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1154 = 14'hd == parameter_2_24 ? phv_data_13 : _GEN_1153; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1155 = 14'he == parameter_2_24 ? phv_data_14 : _GEN_1154; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1156 = 14'hf == parameter_2_24 ? phv_data_15 : _GEN_1155; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1157 = 14'h10 == parameter_2_24 ? phv_data_16 : _GEN_1156; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1158 = 14'h11 == parameter_2_24 ? phv_data_17 : _GEN_1157; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1159 = 14'h12 == parameter_2_24 ? phv_data_18 : _GEN_1158; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1160 = 14'h13 == parameter_2_24 ? phv_data_19 : _GEN_1159; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1161 = 14'h14 == parameter_2_24 ? phv_data_20 : _GEN_1160; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1162 = 14'h15 == parameter_2_24 ? phv_data_21 : _GEN_1161; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1163 = 14'h16 == parameter_2_24 ? phv_data_22 : _GEN_1162; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1164 = 14'h17 == parameter_2_24 ? phv_data_23 : _GEN_1163; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1165 = 14'h18 == parameter_2_24 ? phv_data_24 : _GEN_1164; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1166 = 14'h19 == parameter_2_24 ? phv_data_25 : _GEN_1165; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1167 = 14'h1a == parameter_2_24 ? phv_data_26 : _GEN_1166; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1168 = 14'h1b == parameter_2_24 ? phv_data_27 : _GEN_1167; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1169 = 14'h1c == parameter_2_24 ? phv_data_28 : _GEN_1168; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1170 = 14'h1d == parameter_2_24 ? phv_data_29 : _GEN_1169; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1171 = 14'h1e == parameter_2_24 ? phv_data_30 : _GEN_1170; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1172 = 14'h1f == parameter_2_24 ? phv_data_31 : _GEN_1171; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_25 = vliw_25[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_25 = vliw_25[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_25 = parameter_2_25[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_25 = parameter_2_25[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_25 = {{1'd0}, args_offset_25}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_25 = _total_offset_T_25[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1176 = 3'h1 == total_offset_25 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1177 = 3'h2 == total_offset_25 ? args_2 : _GEN_1176; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1178 = 3'h3 == total_offset_25 ? args_3 : _GEN_1177; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1179 = 3'h4 == total_offset_25 ? args_4 : _GEN_1178; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1180 = 3'h5 == total_offset_25 ? args_5 : _GEN_1179; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1181 = 3'h6 == total_offset_25 ? args_6 : _GEN_1180; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1182 = total_offset_25 < 3'h7 ? _GEN_1181 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_25_0 = 3'h0 < args_length_25 ? _GEN_1182 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1184 = opcode_25 == 4'ha ? field_bytes_25_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1185 = opcode_25 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_978 = opcode_25 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_51 = _T_978 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1186 = opcode_25 == 4'h8 | opcode_25 == 4'hb ? parameter_2_25[7:0] : _GEN_1184; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1187 = opcode_25 == 4'h8 | opcode_25 == 4'hb ? _field_tag_T_51 : _GEN_1185; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1188 = 14'h0 == parameter_2_25 ? phv_data_0 : _GEN_1186; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1189 = 14'h1 == parameter_2_25 ? phv_data_1 : _GEN_1188; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1190 = 14'h2 == parameter_2_25 ? phv_data_2 : _GEN_1189; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1191 = 14'h3 == parameter_2_25 ? phv_data_3 : _GEN_1190; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1192 = 14'h4 == parameter_2_25 ? phv_data_4 : _GEN_1191; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1193 = 14'h5 == parameter_2_25 ? phv_data_5 : _GEN_1192; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1194 = 14'h6 == parameter_2_25 ? phv_data_6 : _GEN_1193; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1195 = 14'h7 == parameter_2_25 ? phv_data_7 : _GEN_1194; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1196 = 14'h8 == parameter_2_25 ? phv_data_8 : _GEN_1195; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1197 = 14'h9 == parameter_2_25 ? phv_data_9 : _GEN_1196; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1198 = 14'ha == parameter_2_25 ? phv_data_10 : _GEN_1197; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1199 = 14'hb == parameter_2_25 ? phv_data_11 : _GEN_1198; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1200 = 14'hc == parameter_2_25 ? phv_data_12 : _GEN_1199; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1201 = 14'hd == parameter_2_25 ? phv_data_13 : _GEN_1200; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1202 = 14'he == parameter_2_25 ? phv_data_14 : _GEN_1201; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1203 = 14'hf == parameter_2_25 ? phv_data_15 : _GEN_1202; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1204 = 14'h10 == parameter_2_25 ? phv_data_16 : _GEN_1203; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1205 = 14'h11 == parameter_2_25 ? phv_data_17 : _GEN_1204; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1206 = 14'h12 == parameter_2_25 ? phv_data_18 : _GEN_1205; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1207 = 14'h13 == parameter_2_25 ? phv_data_19 : _GEN_1206; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1208 = 14'h14 == parameter_2_25 ? phv_data_20 : _GEN_1207; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1209 = 14'h15 == parameter_2_25 ? phv_data_21 : _GEN_1208; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1210 = 14'h16 == parameter_2_25 ? phv_data_22 : _GEN_1209; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1211 = 14'h17 == parameter_2_25 ? phv_data_23 : _GEN_1210; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1212 = 14'h18 == parameter_2_25 ? phv_data_24 : _GEN_1211; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1213 = 14'h19 == parameter_2_25 ? phv_data_25 : _GEN_1212; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1214 = 14'h1a == parameter_2_25 ? phv_data_26 : _GEN_1213; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1215 = 14'h1b == parameter_2_25 ? phv_data_27 : _GEN_1214; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1216 = 14'h1c == parameter_2_25 ? phv_data_28 : _GEN_1215; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1217 = 14'h1d == parameter_2_25 ? phv_data_29 : _GEN_1216; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1218 = 14'h1e == parameter_2_25 ? phv_data_30 : _GEN_1217; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1219 = 14'h1f == parameter_2_25 ? phv_data_31 : _GEN_1218; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_26 = vliw_26[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_26 = vliw_26[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_26 = parameter_2_26[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_26 = parameter_2_26[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_26 = {{1'd0}, args_offset_26}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_26 = _total_offset_T_26[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1223 = 3'h1 == total_offset_26 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1224 = 3'h2 == total_offset_26 ? args_2 : _GEN_1223; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1225 = 3'h3 == total_offset_26 ? args_3 : _GEN_1224; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1226 = 3'h4 == total_offset_26 ? args_4 : _GEN_1225; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1227 = 3'h5 == total_offset_26 ? args_5 : _GEN_1226; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1228 = 3'h6 == total_offset_26 ? args_6 : _GEN_1227; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1229 = total_offset_26 < 3'h7 ? _GEN_1228 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_26_0 = 3'h0 < args_length_26 ? _GEN_1229 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1231 = opcode_26 == 4'ha ? field_bytes_26_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1232 = opcode_26 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1017 = opcode_26 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_53 = _T_1017 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1233 = opcode_26 == 4'h8 | opcode_26 == 4'hb ? parameter_2_26[7:0] : _GEN_1231; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1234 = opcode_26 == 4'h8 | opcode_26 == 4'hb ? _field_tag_T_53 : _GEN_1232; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1235 = 14'h0 == parameter_2_26 ? phv_data_0 : _GEN_1233; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1236 = 14'h1 == parameter_2_26 ? phv_data_1 : _GEN_1235; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1237 = 14'h2 == parameter_2_26 ? phv_data_2 : _GEN_1236; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1238 = 14'h3 == parameter_2_26 ? phv_data_3 : _GEN_1237; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1239 = 14'h4 == parameter_2_26 ? phv_data_4 : _GEN_1238; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1240 = 14'h5 == parameter_2_26 ? phv_data_5 : _GEN_1239; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1241 = 14'h6 == parameter_2_26 ? phv_data_6 : _GEN_1240; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1242 = 14'h7 == parameter_2_26 ? phv_data_7 : _GEN_1241; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1243 = 14'h8 == parameter_2_26 ? phv_data_8 : _GEN_1242; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1244 = 14'h9 == parameter_2_26 ? phv_data_9 : _GEN_1243; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1245 = 14'ha == parameter_2_26 ? phv_data_10 : _GEN_1244; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1246 = 14'hb == parameter_2_26 ? phv_data_11 : _GEN_1245; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1247 = 14'hc == parameter_2_26 ? phv_data_12 : _GEN_1246; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1248 = 14'hd == parameter_2_26 ? phv_data_13 : _GEN_1247; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1249 = 14'he == parameter_2_26 ? phv_data_14 : _GEN_1248; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1250 = 14'hf == parameter_2_26 ? phv_data_15 : _GEN_1249; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1251 = 14'h10 == parameter_2_26 ? phv_data_16 : _GEN_1250; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1252 = 14'h11 == parameter_2_26 ? phv_data_17 : _GEN_1251; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1253 = 14'h12 == parameter_2_26 ? phv_data_18 : _GEN_1252; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1254 = 14'h13 == parameter_2_26 ? phv_data_19 : _GEN_1253; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1255 = 14'h14 == parameter_2_26 ? phv_data_20 : _GEN_1254; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1256 = 14'h15 == parameter_2_26 ? phv_data_21 : _GEN_1255; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1257 = 14'h16 == parameter_2_26 ? phv_data_22 : _GEN_1256; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1258 = 14'h17 == parameter_2_26 ? phv_data_23 : _GEN_1257; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1259 = 14'h18 == parameter_2_26 ? phv_data_24 : _GEN_1258; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1260 = 14'h19 == parameter_2_26 ? phv_data_25 : _GEN_1259; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1261 = 14'h1a == parameter_2_26 ? phv_data_26 : _GEN_1260; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1262 = 14'h1b == parameter_2_26 ? phv_data_27 : _GEN_1261; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1263 = 14'h1c == parameter_2_26 ? phv_data_28 : _GEN_1262; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1264 = 14'h1d == parameter_2_26 ? phv_data_29 : _GEN_1263; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1265 = 14'h1e == parameter_2_26 ? phv_data_30 : _GEN_1264; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1266 = 14'h1f == parameter_2_26 ? phv_data_31 : _GEN_1265; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_27 = vliw_27[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_27 = vliw_27[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_27 = parameter_2_27[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_27 = parameter_2_27[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_27 = {{1'd0}, args_offset_27}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_27 = _total_offset_T_27[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1270 = 3'h1 == total_offset_27 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1271 = 3'h2 == total_offset_27 ? args_2 : _GEN_1270; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1272 = 3'h3 == total_offset_27 ? args_3 : _GEN_1271; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1273 = 3'h4 == total_offset_27 ? args_4 : _GEN_1272; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1274 = 3'h5 == total_offset_27 ? args_5 : _GEN_1273; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1275 = 3'h6 == total_offset_27 ? args_6 : _GEN_1274; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1276 = total_offset_27 < 3'h7 ? _GEN_1275 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_27_0 = 3'h0 < args_length_27 ? _GEN_1276 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1278 = opcode_27 == 4'ha ? field_bytes_27_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1279 = opcode_27 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1056 = opcode_27 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_55 = _T_1056 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1280 = opcode_27 == 4'h8 | opcode_27 == 4'hb ? parameter_2_27[7:0] : _GEN_1278; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1281 = opcode_27 == 4'h8 | opcode_27 == 4'hb ? _field_tag_T_55 : _GEN_1279; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1282 = 14'h0 == parameter_2_27 ? phv_data_0 : _GEN_1280; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1283 = 14'h1 == parameter_2_27 ? phv_data_1 : _GEN_1282; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1284 = 14'h2 == parameter_2_27 ? phv_data_2 : _GEN_1283; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1285 = 14'h3 == parameter_2_27 ? phv_data_3 : _GEN_1284; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1286 = 14'h4 == parameter_2_27 ? phv_data_4 : _GEN_1285; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1287 = 14'h5 == parameter_2_27 ? phv_data_5 : _GEN_1286; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1288 = 14'h6 == parameter_2_27 ? phv_data_6 : _GEN_1287; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1289 = 14'h7 == parameter_2_27 ? phv_data_7 : _GEN_1288; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1290 = 14'h8 == parameter_2_27 ? phv_data_8 : _GEN_1289; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1291 = 14'h9 == parameter_2_27 ? phv_data_9 : _GEN_1290; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1292 = 14'ha == parameter_2_27 ? phv_data_10 : _GEN_1291; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1293 = 14'hb == parameter_2_27 ? phv_data_11 : _GEN_1292; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1294 = 14'hc == parameter_2_27 ? phv_data_12 : _GEN_1293; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1295 = 14'hd == parameter_2_27 ? phv_data_13 : _GEN_1294; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1296 = 14'he == parameter_2_27 ? phv_data_14 : _GEN_1295; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1297 = 14'hf == parameter_2_27 ? phv_data_15 : _GEN_1296; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1298 = 14'h10 == parameter_2_27 ? phv_data_16 : _GEN_1297; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1299 = 14'h11 == parameter_2_27 ? phv_data_17 : _GEN_1298; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1300 = 14'h12 == parameter_2_27 ? phv_data_18 : _GEN_1299; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1301 = 14'h13 == parameter_2_27 ? phv_data_19 : _GEN_1300; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1302 = 14'h14 == parameter_2_27 ? phv_data_20 : _GEN_1301; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1303 = 14'h15 == parameter_2_27 ? phv_data_21 : _GEN_1302; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1304 = 14'h16 == parameter_2_27 ? phv_data_22 : _GEN_1303; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1305 = 14'h17 == parameter_2_27 ? phv_data_23 : _GEN_1304; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1306 = 14'h18 == parameter_2_27 ? phv_data_24 : _GEN_1305; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1307 = 14'h19 == parameter_2_27 ? phv_data_25 : _GEN_1306; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1308 = 14'h1a == parameter_2_27 ? phv_data_26 : _GEN_1307; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1309 = 14'h1b == parameter_2_27 ? phv_data_27 : _GEN_1308; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1310 = 14'h1c == parameter_2_27 ? phv_data_28 : _GEN_1309; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1311 = 14'h1d == parameter_2_27 ? phv_data_29 : _GEN_1310; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1312 = 14'h1e == parameter_2_27 ? phv_data_30 : _GEN_1311; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1313 = 14'h1f == parameter_2_27 ? phv_data_31 : _GEN_1312; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_28 = vliw_28[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_28 = vliw_28[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_28 = parameter_2_28[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_28 = parameter_2_28[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_28 = {{1'd0}, args_offset_28}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_28 = _total_offset_T_28[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1317 = 3'h1 == total_offset_28 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1318 = 3'h2 == total_offset_28 ? args_2 : _GEN_1317; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1319 = 3'h3 == total_offset_28 ? args_3 : _GEN_1318; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1320 = 3'h4 == total_offset_28 ? args_4 : _GEN_1319; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1321 = 3'h5 == total_offset_28 ? args_5 : _GEN_1320; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1322 = 3'h6 == total_offset_28 ? args_6 : _GEN_1321; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1323 = total_offset_28 < 3'h7 ? _GEN_1322 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_28_0 = 3'h0 < args_length_28 ? _GEN_1323 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1325 = opcode_28 == 4'ha ? field_bytes_28_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1326 = opcode_28 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1095 = opcode_28 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_57 = _T_1095 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1327 = opcode_28 == 4'h8 | opcode_28 == 4'hb ? parameter_2_28[7:0] : _GEN_1325; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1328 = opcode_28 == 4'h8 | opcode_28 == 4'hb ? _field_tag_T_57 : _GEN_1326; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1329 = 14'h0 == parameter_2_28 ? phv_data_0 : _GEN_1327; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1330 = 14'h1 == parameter_2_28 ? phv_data_1 : _GEN_1329; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1331 = 14'h2 == parameter_2_28 ? phv_data_2 : _GEN_1330; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1332 = 14'h3 == parameter_2_28 ? phv_data_3 : _GEN_1331; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1333 = 14'h4 == parameter_2_28 ? phv_data_4 : _GEN_1332; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1334 = 14'h5 == parameter_2_28 ? phv_data_5 : _GEN_1333; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1335 = 14'h6 == parameter_2_28 ? phv_data_6 : _GEN_1334; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1336 = 14'h7 == parameter_2_28 ? phv_data_7 : _GEN_1335; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1337 = 14'h8 == parameter_2_28 ? phv_data_8 : _GEN_1336; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1338 = 14'h9 == parameter_2_28 ? phv_data_9 : _GEN_1337; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1339 = 14'ha == parameter_2_28 ? phv_data_10 : _GEN_1338; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1340 = 14'hb == parameter_2_28 ? phv_data_11 : _GEN_1339; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1341 = 14'hc == parameter_2_28 ? phv_data_12 : _GEN_1340; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1342 = 14'hd == parameter_2_28 ? phv_data_13 : _GEN_1341; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1343 = 14'he == parameter_2_28 ? phv_data_14 : _GEN_1342; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1344 = 14'hf == parameter_2_28 ? phv_data_15 : _GEN_1343; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1345 = 14'h10 == parameter_2_28 ? phv_data_16 : _GEN_1344; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1346 = 14'h11 == parameter_2_28 ? phv_data_17 : _GEN_1345; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1347 = 14'h12 == parameter_2_28 ? phv_data_18 : _GEN_1346; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1348 = 14'h13 == parameter_2_28 ? phv_data_19 : _GEN_1347; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1349 = 14'h14 == parameter_2_28 ? phv_data_20 : _GEN_1348; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1350 = 14'h15 == parameter_2_28 ? phv_data_21 : _GEN_1349; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1351 = 14'h16 == parameter_2_28 ? phv_data_22 : _GEN_1350; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1352 = 14'h17 == parameter_2_28 ? phv_data_23 : _GEN_1351; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1353 = 14'h18 == parameter_2_28 ? phv_data_24 : _GEN_1352; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1354 = 14'h19 == parameter_2_28 ? phv_data_25 : _GEN_1353; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1355 = 14'h1a == parameter_2_28 ? phv_data_26 : _GEN_1354; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1356 = 14'h1b == parameter_2_28 ? phv_data_27 : _GEN_1355; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1357 = 14'h1c == parameter_2_28 ? phv_data_28 : _GEN_1356; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1358 = 14'h1d == parameter_2_28 ? phv_data_29 : _GEN_1357; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1359 = 14'h1e == parameter_2_28 ? phv_data_30 : _GEN_1358; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1360 = 14'h1f == parameter_2_28 ? phv_data_31 : _GEN_1359; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_29 = vliw_29[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_29 = vliw_29[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_29 = parameter_2_29[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_29 = parameter_2_29[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_29 = {{1'd0}, args_offset_29}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_29 = _total_offset_T_29[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1364 = 3'h1 == total_offset_29 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1365 = 3'h2 == total_offset_29 ? args_2 : _GEN_1364; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1366 = 3'h3 == total_offset_29 ? args_3 : _GEN_1365; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1367 = 3'h4 == total_offset_29 ? args_4 : _GEN_1366; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1368 = 3'h5 == total_offset_29 ? args_5 : _GEN_1367; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1369 = 3'h6 == total_offset_29 ? args_6 : _GEN_1368; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1370 = total_offset_29 < 3'h7 ? _GEN_1369 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_29_0 = 3'h0 < args_length_29 ? _GEN_1370 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1372 = opcode_29 == 4'ha ? field_bytes_29_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1373 = opcode_29 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1134 = opcode_29 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_59 = _T_1134 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1374 = opcode_29 == 4'h8 | opcode_29 == 4'hb ? parameter_2_29[7:0] : _GEN_1372; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1375 = opcode_29 == 4'h8 | opcode_29 == 4'hb ? _field_tag_T_59 : _GEN_1373; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1376 = 14'h0 == parameter_2_29 ? phv_data_0 : _GEN_1374; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1377 = 14'h1 == parameter_2_29 ? phv_data_1 : _GEN_1376; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1378 = 14'h2 == parameter_2_29 ? phv_data_2 : _GEN_1377; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1379 = 14'h3 == parameter_2_29 ? phv_data_3 : _GEN_1378; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1380 = 14'h4 == parameter_2_29 ? phv_data_4 : _GEN_1379; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1381 = 14'h5 == parameter_2_29 ? phv_data_5 : _GEN_1380; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1382 = 14'h6 == parameter_2_29 ? phv_data_6 : _GEN_1381; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1383 = 14'h7 == parameter_2_29 ? phv_data_7 : _GEN_1382; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1384 = 14'h8 == parameter_2_29 ? phv_data_8 : _GEN_1383; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1385 = 14'h9 == parameter_2_29 ? phv_data_9 : _GEN_1384; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1386 = 14'ha == parameter_2_29 ? phv_data_10 : _GEN_1385; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1387 = 14'hb == parameter_2_29 ? phv_data_11 : _GEN_1386; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1388 = 14'hc == parameter_2_29 ? phv_data_12 : _GEN_1387; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1389 = 14'hd == parameter_2_29 ? phv_data_13 : _GEN_1388; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1390 = 14'he == parameter_2_29 ? phv_data_14 : _GEN_1389; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1391 = 14'hf == parameter_2_29 ? phv_data_15 : _GEN_1390; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1392 = 14'h10 == parameter_2_29 ? phv_data_16 : _GEN_1391; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1393 = 14'h11 == parameter_2_29 ? phv_data_17 : _GEN_1392; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1394 = 14'h12 == parameter_2_29 ? phv_data_18 : _GEN_1393; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1395 = 14'h13 == parameter_2_29 ? phv_data_19 : _GEN_1394; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1396 = 14'h14 == parameter_2_29 ? phv_data_20 : _GEN_1395; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1397 = 14'h15 == parameter_2_29 ? phv_data_21 : _GEN_1396; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1398 = 14'h16 == parameter_2_29 ? phv_data_22 : _GEN_1397; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1399 = 14'h17 == parameter_2_29 ? phv_data_23 : _GEN_1398; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1400 = 14'h18 == parameter_2_29 ? phv_data_24 : _GEN_1399; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1401 = 14'h19 == parameter_2_29 ? phv_data_25 : _GEN_1400; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1402 = 14'h1a == parameter_2_29 ? phv_data_26 : _GEN_1401; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1403 = 14'h1b == parameter_2_29 ? phv_data_27 : _GEN_1402; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1404 = 14'h1c == parameter_2_29 ? phv_data_28 : _GEN_1403; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1405 = 14'h1d == parameter_2_29 ? phv_data_29 : _GEN_1404; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1406 = 14'h1e == parameter_2_29 ? phv_data_30 : _GEN_1405; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1407 = 14'h1f == parameter_2_29 ? phv_data_31 : _GEN_1406; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_30 = vliw_30[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_30 = vliw_30[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_30 = parameter_2_30[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_30 = parameter_2_30[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_30 = {{1'd0}, args_offset_30}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_30 = _total_offset_T_30[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1411 = 3'h1 == total_offset_30 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1412 = 3'h2 == total_offset_30 ? args_2 : _GEN_1411; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1413 = 3'h3 == total_offset_30 ? args_3 : _GEN_1412; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1414 = 3'h4 == total_offset_30 ? args_4 : _GEN_1413; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1415 = 3'h5 == total_offset_30 ? args_5 : _GEN_1414; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1416 = 3'h6 == total_offset_30 ? args_6 : _GEN_1415; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1417 = total_offset_30 < 3'h7 ? _GEN_1416 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_30_0 = 3'h0 < args_length_30 ? _GEN_1417 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1419 = opcode_30 == 4'ha ? field_bytes_30_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1420 = opcode_30 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1173 = opcode_30 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_61 = _T_1173 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1421 = opcode_30 == 4'h8 | opcode_30 == 4'hb ? parameter_2_30[7:0] : _GEN_1419; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1422 = opcode_30 == 4'h8 | opcode_30 == 4'hb ? _field_tag_T_61 : _GEN_1420; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1423 = 14'h0 == parameter_2_30 ? phv_data_0 : _GEN_1421; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1424 = 14'h1 == parameter_2_30 ? phv_data_1 : _GEN_1423; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1425 = 14'h2 == parameter_2_30 ? phv_data_2 : _GEN_1424; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1426 = 14'h3 == parameter_2_30 ? phv_data_3 : _GEN_1425; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1427 = 14'h4 == parameter_2_30 ? phv_data_4 : _GEN_1426; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1428 = 14'h5 == parameter_2_30 ? phv_data_5 : _GEN_1427; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1429 = 14'h6 == parameter_2_30 ? phv_data_6 : _GEN_1428; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1430 = 14'h7 == parameter_2_30 ? phv_data_7 : _GEN_1429; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1431 = 14'h8 == parameter_2_30 ? phv_data_8 : _GEN_1430; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1432 = 14'h9 == parameter_2_30 ? phv_data_9 : _GEN_1431; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1433 = 14'ha == parameter_2_30 ? phv_data_10 : _GEN_1432; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1434 = 14'hb == parameter_2_30 ? phv_data_11 : _GEN_1433; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1435 = 14'hc == parameter_2_30 ? phv_data_12 : _GEN_1434; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1436 = 14'hd == parameter_2_30 ? phv_data_13 : _GEN_1435; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1437 = 14'he == parameter_2_30 ? phv_data_14 : _GEN_1436; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1438 = 14'hf == parameter_2_30 ? phv_data_15 : _GEN_1437; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1439 = 14'h10 == parameter_2_30 ? phv_data_16 : _GEN_1438; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1440 = 14'h11 == parameter_2_30 ? phv_data_17 : _GEN_1439; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1441 = 14'h12 == parameter_2_30 ? phv_data_18 : _GEN_1440; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1442 = 14'h13 == parameter_2_30 ? phv_data_19 : _GEN_1441; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1443 = 14'h14 == parameter_2_30 ? phv_data_20 : _GEN_1442; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1444 = 14'h15 == parameter_2_30 ? phv_data_21 : _GEN_1443; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1445 = 14'h16 == parameter_2_30 ? phv_data_22 : _GEN_1444; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1446 = 14'h17 == parameter_2_30 ? phv_data_23 : _GEN_1445; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1447 = 14'h18 == parameter_2_30 ? phv_data_24 : _GEN_1446; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1448 = 14'h19 == parameter_2_30 ? phv_data_25 : _GEN_1447; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1449 = 14'h1a == parameter_2_30 ? phv_data_26 : _GEN_1448; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1450 = 14'h1b == parameter_2_30 ? phv_data_27 : _GEN_1449; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1451 = 14'h1c == parameter_2_30 ? phv_data_28 : _GEN_1450; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1452 = 14'h1d == parameter_2_30 ? phv_data_29 : _GEN_1451; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1453 = 14'h1e == parameter_2_30 ? phv_data_30 : _GEN_1452; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1454 = 14'h1f == parameter_2_30 ? phv_data_31 : _GEN_1453; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_31 = vliw_31[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_31 = vliw_31[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_31 = parameter_2_31[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_31 = parameter_2_31[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_31 = {{1'd0}, args_offset_31}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_31 = _total_offset_T_31[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1458 = 3'h1 == total_offset_31 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1459 = 3'h2 == total_offset_31 ? args_2 : _GEN_1458; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1460 = 3'h3 == total_offset_31 ? args_3 : _GEN_1459; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1461 = 3'h4 == total_offset_31 ? args_4 : _GEN_1460; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1462 = 3'h5 == total_offset_31 ? args_5 : _GEN_1461; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1463 = 3'h6 == total_offset_31 ? args_6 : _GEN_1462; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1464 = total_offset_31 < 3'h7 ? _GEN_1463 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_31_0 = 3'h0 < args_length_31 ? _GEN_1464 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_1466 = opcode_31 == 4'ha ? field_bytes_31_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1467 = opcode_31 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1212 = opcode_31 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_63 = _T_1212 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_1468 = opcode_31 == 4'h8 | opcode_31 == 4'hb ? parameter_2_31[7:0] : _GEN_1466; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_1469 = opcode_31 == 4'h8 | opcode_31 == 4'hb ? _field_tag_T_63 : _GEN_1467; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_1470 = 14'h0 == parameter_2_31 ? phv_data_0 : _GEN_1468; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1471 = 14'h1 == parameter_2_31 ? phv_data_1 : _GEN_1470; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1472 = 14'h2 == parameter_2_31 ? phv_data_2 : _GEN_1471; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1473 = 14'h3 == parameter_2_31 ? phv_data_3 : _GEN_1472; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1474 = 14'h4 == parameter_2_31 ? phv_data_4 : _GEN_1473; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1475 = 14'h5 == parameter_2_31 ? phv_data_5 : _GEN_1474; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1476 = 14'h6 == parameter_2_31 ? phv_data_6 : _GEN_1475; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1477 = 14'h7 == parameter_2_31 ? phv_data_7 : _GEN_1476; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1478 = 14'h8 == parameter_2_31 ? phv_data_8 : _GEN_1477; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1479 = 14'h9 == parameter_2_31 ? phv_data_9 : _GEN_1478; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1480 = 14'ha == parameter_2_31 ? phv_data_10 : _GEN_1479; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1481 = 14'hb == parameter_2_31 ? phv_data_11 : _GEN_1480; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1482 = 14'hc == parameter_2_31 ? phv_data_12 : _GEN_1481; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1483 = 14'hd == parameter_2_31 ? phv_data_13 : _GEN_1482; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1484 = 14'he == parameter_2_31 ? phv_data_14 : _GEN_1483; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1485 = 14'hf == parameter_2_31 ? phv_data_15 : _GEN_1484; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1486 = 14'h10 == parameter_2_31 ? phv_data_16 : _GEN_1485; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1487 = 14'h11 == parameter_2_31 ? phv_data_17 : _GEN_1486; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1488 = 14'h12 == parameter_2_31 ? phv_data_18 : _GEN_1487; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1489 = 14'h13 == parameter_2_31 ? phv_data_19 : _GEN_1488; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1490 = 14'h14 == parameter_2_31 ? phv_data_20 : _GEN_1489; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1491 = 14'h15 == parameter_2_31 ? phv_data_21 : _GEN_1490; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1492 = 14'h16 == parameter_2_31 ? phv_data_22 : _GEN_1491; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1493 = 14'h17 == parameter_2_31 ? phv_data_23 : _GEN_1492; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1494 = 14'h18 == parameter_2_31 ? phv_data_24 : _GEN_1493; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1495 = 14'h19 == parameter_2_31 ? phv_data_25 : _GEN_1494; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1496 = 14'h1a == parameter_2_31 ? phv_data_26 : _GEN_1495; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1497 = 14'h1b == parameter_2_31 ? phv_data_27 : _GEN_1496; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1498 = 14'h1c == parameter_2_31 ? phv_data_28 : _GEN_1497; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1499 = 14'h1d == parameter_2_31 ? phv_data_29 : _GEN_1498; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1500 = 14'h1e == parameter_2_31 ? phv_data_30 : _GEN_1499; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_1501 = 14'h1f == parameter_2_31 ? phv_data_31 : _GEN_1500; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_32 = vliw_32[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo = vliw_32[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_32 = field_data_lo[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_32 = field_data_lo[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_32 = {{1'd0}, args_offset_32}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_32 = _total_offset_T_32[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1505 = 3'h1 == total_offset_32 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1506 = 3'h2 == total_offset_32 ? args_2 : _GEN_1505; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1507 = 3'h3 == total_offset_32 ? args_3 : _GEN_1506; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1508 = 3'h4 == total_offset_32 ? args_4 : _GEN_1507; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1509 = 3'h5 == total_offset_32 ? args_5 : _GEN_1508; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1510 = 3'h6 == total_offset_32 ? args_6 : _GEN_1509; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1511 = total_offset_32 < 3'h7 ? _GEN_1510 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_32_1 = 3'h0 < args_length_32 ? _GEN_1511 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_33 = args_offset_32 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1514 = 3'h1 == total_offset_33 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1515 = 3'h2 == total_offset_33 ? args_2 : _GEN_1514; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1516 = 3'h3 == total_offset_33 ? args_3 : _GEN_1515; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1517 = 3'h4 == total_offset_33 ? args_4 : _GEN_1516; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1518 = 3'h5 == total_offset_33 ? args_5 : _GEN_1517; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1519 = 3'h6 == total_offset_33 ? args_6 : _GEN_1518; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1520 = total_offset_33 < 3'h7 ? _GEN_1519 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_32_0 = 3'h1 < args_length_32 ? _GEN_1520 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_32 = {field_bytes_32_0,field_bytes_32_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1522 = opcode_32 == 4'ha ? _field_data_T_32 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1523 = opcode_32 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1253 = opcode_32 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi = field_data_lo[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_35 = {field_data_hi,field_data_lo}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_65 = _T_1253 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1524 = opcode_32 == 4'h8 | opcode_32 == 4'hb ? _field_data_T_35 : _GEN_1522; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1525 = opcode_32 == 4'h8 | opcode_32 == 4'hb ? _field_tag_T_65 : _GEN_1523; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _field_data_T_36 = {phv_data_32,phv_data_33}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1526 = 14'h20 == field_data_lo ? _field_data_T_36 : _GEN_1524; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_37 = {phv_data_34,phv_data_35}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1527 = 14'h21 == field_data_lo ? _field_data_T_37 : _GEN_1526; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_38 = {phv_data_36,phv_data_37}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1528 = 14'h22 == field_data_lo ? _field_data_T_38 : _GEN_1527; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_39 = {phv_data_38,phv_data_39}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1529 = 14'h23 == field_data_lo ? _field_data_T_39 : _GEN_1528; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_40 = {phv_data_40,phv_data_41}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1530 = 14'h24 == field_data_lo ? _field_data_T_40 : _GEN_1529; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_41 = {phv_data_42,phv_data_43}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1531 = 14'h25 == field_data_lo ? _field_data_T_41 : _GEN_1530; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_42 = {phv_data_44,phv_data_45}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1532 = 14'h26 == field_data_lo ? _field_data_T_42 : _GEN_1531; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_43 = {phv_data_46,phv_data_47}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1533 = 14'h27 == field_data_lo ? _field_data_T_43 : _GEN_1532; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_44 = {phv_data_48,phv_data_49}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1534 = 14'h28 == field_data_lo ? _field_data_T_44 : _GEN_1533; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_45 = {phv_data_50,phv_data_51}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1535 = 14'h29 == field_data_lo ? _field_data_T_45 : _GEN_1534; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_46 = {phv_data_52,phv_data_53}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1536 = 14'h2a == field_data_lo ? _field_data_T_46 : _GEN_1535; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_47 = {phv_data_54,phv_data_55}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1537 = 14'h2b == field_data_lo ? _field_data_T_47 : _GEN_1536; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_48 = {phv_data_56,phv_data_57}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1538 = 14'h2c == field_data_lo ? _field_data_T_48 : _GEN_1537; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_49 = {phv_data_58,phv_data_59}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1539 = 14'h2d == field_data_lo ? _field_data_T_49 : _GEN_1538; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_50 = {phv_data_60,phv_data_61}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1540 = 14'h2e == field_data_lo ? _field_data_T_50 : _GEN_1539; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_51 = {phv_data_62,phv_data_63}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1541 = 14'h2f == field_data_lo ? _field_data_T_51 : _GEN_1540; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_52 = {phv_data_64,phv_data_65}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1542 = 14'h30 == field_data_lo ? _field_data_T_52 : _GEN_1541; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_53 = {phv_data_66,phv_data_67}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1543 = 14'h31 == field_data_lo ? _field_data_T_53 : _GEN_1542; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_54 = {phv_data_68,phv_data_69}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1544 = 14'h32 == field_data_lo ? _field_data_T_54 : _GEN_1543; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_55 = {phv_data_70,phv_data_71}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1545 = 14'h33 == field_data_lo ? _field_data_T_55 : _GEN_1544; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_56 = {phv_data_72,phv_data_73}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1546 = 14'h34 == field_data_lo ? _field_data_T_56 : _GEN_1545; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_57 = {phv_data_74,phv_data_75}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1547 = 14'h35 == field_data_lo ? _field_data_T_57 : _GEN_1546; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_58 = {phv_data_76,phv_data_77}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1548 = 14'h36 == field_data_lo ? _field_data_T_58 : _GEN_1547; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_59 = {phv_data_78,phv_data_79}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1549 = 14'h37 == field_data_lo ? _field_data_T_59 : _GEN_1548; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_60 = {phv_data_80,phv_data_81}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1550 = 14'h38 == field_data_lo ? _field_data_T_60 : _GEN_1549; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_61 = {phv_data_82,phv_data_83}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1551 = 14'h39 == field_data_lo ? _field_data_T_61 : _GEN_1550; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_62 = {phv_data_84,phv_data_85}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1552 = 14'h3a == field_data_lo ? _field_data_T_62 : _GEN_1551; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_63 = {phv_data_86,phv_data_87}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1553 = 14'h3b == field_data_lo ? _field_data_T_63 : _GEN_1552; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_64 = {phv_data_88,phv_data_89}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1554 = 14'h3c == field_data_lo ? _field_data_T_64 : _GEN_1553; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_65 = {phv_data_90,phv_data_91}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1555 = 14'h3d == field_data_lo ? _field_data_T_65 : _GEN_1554; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_66 = {phv_data_92,phv_data_93}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1556 = 14'h3e == field_data_lo ? _field_data_T_66 : _GEN_1555; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_67 = {phv_data_94,phv_data_95}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1557 = 14'h3f == field_data_lo ? _field_data_T_67 : _GEN_1556; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_68 = {phv_data_96,phv_data_97}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1558 = 14'h40 == field_data_lo ? _field_data_T_68 : _GEN_1557; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_69 = {phv_data_98,phv_data_99}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1559 = 14'h41 == field_data_lo ? _field_data_T_69 : _GEN_1558; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_70 = {phv_data_100,phv_data_101}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1560 = 14'h42 == field_data_lo ? _field_data_T_70 : _GEN_1559; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_71 = {phv_data_102,phv_data_103}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1561 = 14'h43 == field_data_lo ? _field_data_T_71 : _GEN_1560; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_72 = {phv_data_104,phv_data_105}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1562 = 14'h44 == field_data_lo ? _field_data_T_72 : _GEN_1561; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_73 = {phv_data_106,phv_data_107}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1563 = 14'h45 == field_data_lo ? _field_data_T_73 : _GEN_1562; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_74 = {phv_data_108,phv_data_109}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1564 = 14'h46 == field_data_lo ? _field_data_T_74 : _GEN_1563; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_75 = {phv_data_110,phv_data_111}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1565 = 14'h47 == field_data_lo ? _field_data_T_75 : _GEN_1564; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_76 = {phv_data_112,phv_data_113}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1566 = 14'h48 == field_data_lo ? _field_data_T_76 : _GEN_1565; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_77 = {phv_data_114,phv_data_115}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1567 = 14'h49 == field_data_lo ? _field_data_T_77 : _GEN_1566; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_78 = {phv_data_116,phv_data_117}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1568 = 14'h4a == field_data_lo ? _field_data_T_78 : _GEN_1567; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_79 = {phv_data_118,phv_data_119}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1569 = 14'h4b == field_data_lo ? _field_data_T_79 : _GEN_1568; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_80 = {phv_data_120,phv_data_121}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1570 = 14'h4c == field_data_lo ? _field_data_T_80 : _GEN_1569; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_81 = {phv_data_122,phv_data_123}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1571 = 14'h4d == field_data_lo ? _field_data_T_81 : _GEN_1570; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_82 = {phv_data_124,phv_data_125}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1572 = 14'h4e == field_data_lo ? _field_data_T_82 : _GEN_1571; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_83 = {phv_data_126,phv_data_127}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1573 = 14'h4f == field_data_lo ? _field_data_T_83 : _GEN_1572; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_33 = vliw_33[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_1 = vliw_33[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_33 = field_data_lo_1[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_33 = field_data_lo_1[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_34 = {{1'd0}, args_offset_33}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_34 = _total_offset_T_34[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1577 = 3'h1 == total_offset_34 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1578 = 3'h2 == total_offset_34 ? args_2 : _GEN_1577; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1579 = 3'h3 == total_offset_34 ? args_3 : _GEN_1578; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1580 = 3'h4 == total_offset_34 ? args_4 : _GEN_1579; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1581 = 3'h5 == total_offset_34 ? args_5 : _GEN_1580; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1582 = 3'h6 == total_offset_34 ? args_6 : _GEN_1581; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1583 = total_offset_34 < 3'h7 ? _GEN_1582 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_33_1 = 3'h0 < args_length_33 ? _GEN_1583 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_35 = args_offset_33 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1586 = 3'h1 == total_offset_35 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1587 = 3'h2 == total_offset_35 ? args_2 : _GEN_1586; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1588 = 3'h3 == total_offset_35 ? args_3 : _GEN_1587; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1589 = 3'h4 == total_offset_35 ? args_4 : _GEN_1588; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1590 = 3'h5 == total_offset_35 ? args_5 : _GEN_1589; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1591 = 3'h6 == total_offset_35 ? args_6 : _GEN_1590; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1592 = total_offset_35 < 3'h7 ? _GEN_1591 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_33_0 = 3'h1 < args_length_33 ? _GEN_1592 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_84 = {field_bytes_33_0,field_bytes_33_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1594 = opcode_33 == 4'ha ? _field_data_T_84 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1595 = opcode_33 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1310 = opcode_33 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_1 = field_data_lo_1[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_87 = {field_data_hi_1,field_data_lo_1}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_67 = _T_1310 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1596 = opcode_33 == 4'h8 | opcode_33 == 4'hb ? _field_data_T_87 : _GEN_1594; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1597 = opcode_33 == 4'h8 | opcode_33 == 4'hb ? _field_tag_T_67 : _GEN_1595; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1598 = 14'h20 == field_data_lo_1 ? _field_data_T_36 : _GEN_1596; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1599 = 14'h21 == field_data_lo_1 ? _field_data_T_37 : _GEN_1598; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1600 = 14'h22 == field_data_lo_1 ? _field_data_T_38 : _GEN_1599; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1601 = 14'h23 == field_data_lo_1 ? _field_data_T_39 : _GEN_1600; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1602 = 14'h24 == field_data_lo_1 ? _field_data_T_40 : _GEN_1601; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1603 = 14'h25 == field_data_lo_1 ? _field_data_T_41 : _GEN_1602; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1604 = 14'h26 == field_data_lo_1 ? _field_data_T_42 : _GEN_1603; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1605 = 14'h27 == field_data_lo_1 ? _field_data_T_43 : _GEN_1604; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1606 = 14'h28 == field_data_lo_1 ? _field_data_T_44 : _GEN_1605; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1607 = 14'h29 == field_data_lo_1 ? _field_data_T_45 : _GEN_1606; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1608 = 14'h2a == field_data_lo_1 ? _field_data_T_46 : _GEN_1607; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1609 = 14'h2b == field_data_lo_1 ? _field_data_T_47 : _GEN_1608; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1610 = 14'h2c == field_data_lo_1 ? _field_data_T_48 : _GEN_1609; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1611 = 14'h2d == field_data_lo_1 ? _field_data_T_49 : _GEN_1610; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1612 = 14'h2e == field_data_lo_1 ? _field_data_T_50 : _GEN_1611; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1613 = 14'h2f == field_data_lo_1 ? _field_data_T_51 : _GEN_1612; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1614 = 14'h30 == field_data_lo_1 ? _field_data_T_52 : _GEN_1613; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1615 = 14'h31 == field_data_lo_1 ? _field_data_T_53 : _GEN_1614; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1616 = 14'h32 == field_data_lo_1 ? _field_data_T_54 : _GEN_1615; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1617 = 14'h33 == field_data_lo_1 ? _field_data_T_55 : _GEN_1616; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1618 = 14'h34 == field_data_lo_1 ? _field_data_T_56 : _GEN_1617; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1619 = 14'h35 == field_data_lo_1 ? _field_data_T_57 : _GEN_1618; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1620 = 14'h36 == field_data_lo_1 ? _field_data_T_58 : _GEN_1619; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1621 = 14'h37 == field_data_lo_1 ? _field_data_T_59 : _GEN_1620; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1622 = 14'h38 == field_data_lo_1 ? _field_data_T_60 : _GEN_1621; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1623 = 14'h39 == field_data_lo_1 ? _field_data_T_61 : _GEN_1622; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1624 = 14'h3a == field_data_lo_1 ? _field_data_T_62 : _GEN_1623; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1625 = 14'h3b == field_data_lo_1 ? _field_data_T_63 : _GEN_1624; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1626 = 14'h3c == field_data_lo_1 ? _field_data_T_64 : _GEN_1625; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1627 = 14'h3d == field_data_lo_1 ? _field_data_T_65 : _GEN_1626; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1628 = 14'h3e == field_data_lo_1 ? _field_data_T_66 : _GEN_1627; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1629 = 14'h3f == field_data_lo_1 ? _field_data_T_67 : _GEN_1628; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1630 = 14'h40 == field_data_lo_1 ? _field_data_T_68 : _GEN_1629; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1631 = 14'h41 == field_data_lo_1 ? _field_data_T_69 : _GEN_1630; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1632 = 14'h42 == field_data_lo_1 ? _field_data_T_70 : _GEN_1631; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1633 = 14'h43 == field_data_lo_1 ? _field_data_T_71 : _GEN_1632; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1634 = 14'h44 == field_data_lo_1 ? _field_data_T_72 : _GEN_1633; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1635 = 14'h45 == field_data_lo_1 ? _field_data_T_73 : _GEN_1634; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1636 = 14'h46 == field_data_lo_1 ? _field_data_T_74 : _GEN_1635; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1637 = 14'h47 == field_data_lo_1 ? _field_data_T_75 : _GEN_1636; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1638 = 14'h48 == field_data_lo_1 ? _field_data_T_76 : _GEN_1637; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1639 = 14'h49 == field_data_lo_1 ? _field_data_T_77 : _GEN_1638; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1640 = 14'h4a == field_data_lo_1 ? _field_data_T_78 : _GEN_1639; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1641 = 14'h4b == field_data_lo_1 ? _field_data_T_79 : _GEN_1640; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1642 = 14'h4c == field_data_lo_1 ? _field_data_T_80 : _GEN_1641; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1643 = 14'h4d == field_data_lo_1 ? _field_data_T_81 : _GEN_1642; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1644 = 14'h4e == field_data_lo_1 ? _field_data_T_82 : _GEN_1643; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1645 = 14'h4f == field_data_lo_1 ? _field_data_T_83 : _GEN_1644; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_34 = vliw_34[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_2 = vliw_34[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_34 = field_data_lo_2[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_34 = field_data_lo_2[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_36 = {{1'd0}, args_offset_34}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_36 = _total_offset_T_36[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1649 = 3'h1 == total_offset_36 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1650 = 3'h2 == total_offset_36 ? args_2 : _GEN_1649; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1651 = 3'h3 == total_offset_36 ? args_3 : _GEN_1650; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1652 = 3'h4 == total_offset_36 ? args_4 : _GEN_1651; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1653 = 3'h5 == total_offset_36 ? args_5 : _GEN_1652; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1654 = 3'h6 == total_offset_36 ? args_6 : _GEN_1653; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1655 = total_offset_36 < 3'h7 ? _GEN_1654 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_34_1 = 3'h0 < args_length_34 ? _GEN_1655 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_37 = args_offset_34 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1658 = 3'h1 == total_offset_37 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1659 = 3'h2 == total_offset_37 ? args_2 : _GEN_1658; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1660 = 3'h3 == total_offset_37 ? args_3 : _GEN_1659; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1661 = 3'h4 == total_offset_37 ? args_4 : _GEN_1660; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1662 = 3'h5 == total_offset_37 ? args_5 : _GEN_1661; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1663 = 3'h6 == total_offset_37 ? args_6 : _GEN_1662; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1664 = total_offset_37 < 3'h7 ? _GEN_1663 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_34_0 = 3'h1 < args_length_34 ? _GEN_1664 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_136 = {field_bytes_34_0,field_bytes_34_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1666 = opcode_34 == 4'ha ? _field_data_T_136 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1667 = opcode_34 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1367 = opcode_34 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_2 = field_data_lo_2[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_139 = {field_data_hi_2,field_data_lo_2}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_69 = _T_1367 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1668 = opcode_34 == 4'h8 | opcode_34 == 4'hb ? _field_data_T_139 : _GEN_1666; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1669 = opcode_34 == 4'h8 | opcode_34 == 4'hb ? _field_tag_T_69 : _GEN_1667; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1670 = 14'h20 == field_data_lo_2 ? _field_data_T_36 : _GEN_1668; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1671 = 14'h21 == field_data_lo_2 ? _field_data_T_37 : _GEN_1670; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1672 = 14'h22 == field_data_lo_2 ? _field_data_T_38 : _GEN_1671; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1673 = 14'h23 == field_data_lo_2 ? _field_data_T_39 : _GEN_1672; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1674 = 14'h24 == field_data_lo_2 ? _field_data_T_40 : _GEN_1673; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1675 = 14'h25 == field_data_lo_2 ? _field_data_T_41 : _GEN_1674; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1676 = 14'h26 == field_data_lo_2 ? _field_data_T_42 : _GEN_1675; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1677 = 14'h27 == field_data_lo_2 ? _field_data_T_43 : _GEN_1676; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1678 = 14'h28 == field_data_lo_2 ? _field_data_T_44 : _GEN_1677; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1679 = 14'h29 == field_data_lo_2 ? _field_data_T_45 : _GEN_1678; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1680 = 14'h2a == field_data_lo_2 ? _field_data_T_46 : _GEN_1679; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1681 = 14'h2b == field_data_lo_2 ? _field_data_T_47 : _GEN_1680; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1682 = 14'h2c == field_data_lo_2 ? _field_data_T_48 : _GEN_1681; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1683 = 14'h2d == field_data_lo_2 ? _field_data_T_49 : _GEN_1682; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1684 = 14'h2e == field_data_lo_2 ? _field_data_T_50 : _GEN_1683; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1685 = 14'h2f == field_data_lo_2 ? _field_data_T_51 : _GEN_1684; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1686 = 14'h30 == field_data_lo_2 ? _field_data_T_52 : _GEN_1685; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1687 = 14'h31 == field_data_lo_2 ? _field_data_T_53 : _GEN_1686; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1688 = 14'h32 == field_data_lo_2 ? _field_data_T_54 : _GEN_1687; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1689 = 14'h33 == field_data_lo_2 ? _field_data_T_55 : _GEN_1688; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1690 = 14'h34 == field_data_lo_2 ? _field_data_T_56 : _GEN_1689; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1691 = 14'h35 == field_data_lo_2 ? _field_data_T_57 : _GEN_1690; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1692 = 14'h36 == field_data_lo_2 ? _field_data_T_58 : _GEN_1691; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1693 = 14'h37 == field_data_lo_2 ? _field_data_T_59 : _GEN_1692; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1694 = 14'h38 == field_data_lo_2 ? _field_data_T_60 : _GEN_1693; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1695 = 14'h39 == field_data_lo_2 ? _field_data_T_61 : _GEN_1694; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1696 = 14'h3a == field_data_lo_2 ? _field_data_T_62 : _GEN_1695; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1697 = 14'h3b == field_data_lo_2 ? _field_data_T_63 : _GEN_1696; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1698 = 14'h3c == field_data_lo_2 ? _field_data_T_64 : _GEN_1697; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1699 = 14'h3d == field_data_lo_2 ? _field_data_T_65 : _GEN_1698; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1700 = 14'h3e == field_data_lo_2 ? _field_data_T_66 : _GEN_1699; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1701 = 14'h3f == field_data_lo_2 ? _field_data_T_67 : _GEN_1700; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1702 = 14'h40 == field_data_lo_2 ? _field_data_T_68 : _GEN_1701; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1703 = 14'h41 == field_data_lo_2 ? _field_data_T_69 : _GEN_1702; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1704 = 14'h42 == field_data_lo_2 ? _field_data_T_70 : _GEN_1703; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1705 = 14'h43 == field_data_lo_2 ? _field_data_T_71 : _GEN_1704; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1706 = 14'h44 == field_data_lo_2 ? _field_data_T_72 : _GEN_1705; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1707 = 14'h45 == field_data_lo_2 ? _field_data_T_73 : _GEN_1706; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1708 = 14'h46 == field_data_lo_2 ? _field_data_T_74 : _GEN_1707; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1709 = 14'h47 == field_data_lo_2 ? _field_data_T_75 : _GEN_1708; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1710 = 14'h48 == field_data_lo_2 ? _field_data_T_76 : _GEN_1709; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1711 = 14'h49 == field_data_lo_2 ? _field_data_T_77 : _GEN_1710; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1712 = 14'h4a == field_data_lo_2 ? _field_data_T_78 : _GEN_1711; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1713 = 14'h4b == field_data_lo_2 ? _field_data_T_79 : _GEN_1712; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1714 = 14'h4c == field_data_lo_2 ? _field_data_T_80 : _GEN_1713; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1715 = 14'h4d == field_data_lo_2 ? _field_data_T_81 : _GEN_1714; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1716 = 14'h4e == field_data_lo_2 ? _field_data_T_82 : _GEN_1715; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1717 = 14'h4f == field_data_lo_2 ? _field_data_T_83 : _GEN_1716; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_35 = vliw_35[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_3 = vliw_35[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_35 = field_data_lo_3[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_35 = field_data_lo_3[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_38 = {{1'd0}, args_offset_35}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_38 = _total_offset_T_38[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1721 = 3'h1 == total_offset_38 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1722 = 3'h2 == total_offset_38 ? args_2 : _GEN_1721; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1723 = 3'h3 == total_offset_38 ? args_3 : _GEN_1722; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1724 = 3'h4 == total_offset_38 ? args_4 : _GEN_1723; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1725 = 3'h5 == total_offset_38 ? args_5 : _GEN_1724; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1726 = 3'h6 == total_offset_38 ? args_6 : _GEN_1725; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1727 = total_offset_38 < 3'h7 ? _GEN_1726 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_35_1 = 3'h0 < args_length_35 ? _GEN_1727 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_39 = args_offset_35 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1730 = 3'h1 == total_offset_39 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1731 = 3'h2 == total_offset_39 ? args_2 : _GEN_1730; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1732 = 3'h3 == total_offset_39 ? args_3 : _GEN_1731; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1733 = 3'h4 == total_offset_39 ? args_4 : _GEN_1732; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1734 = 3'h5 == total_offset_39 ? args_5 : _GEN_1733; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1735 = 3'h6 == total_offset_39 ? args_6 : _GEN_1734; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1736 = total_offset_39 < 3'h7 ? _GEN_1735 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_35_0 = 3'h1 < args_length_35 ? _GEN_1736 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_188 = {field_bytes_35_0,field_bytes_35_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1738 = opcode_35 == 4'ha ? _field_data_T_188 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1739 = opcode_35 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1424 = opcode_35 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_3 = field_data_lo_3[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_191 = {field_data_hi_3,field_data_lo_3}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_71 = _T_1424 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1740 = opcode_35 == 4'h8 | opcode_35 == 4'hb ? _field_data_T_191 : _GEN_1738; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1741 = opcode_35 == 4'h8 | opcode_35 == 4'hb ? _field_tag_T_71 : _GEN_1739; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1742 = 14'h20 == field_data_lo_3 ? _field_data_T_36 : _GEN_1740; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1743 = 14'h21 == field_data_lo_3 ? _field_data_T_37 : _GEN_1742; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1744 = 14'h22 == field_data_lo_3 ? _field_data_T_38 : _GEN_1743; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1745 = 14'h23 == field_data_lo_3 ? _field_data_T_39 : _GEN_1744; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1746 = 14'h24 == field_data_lo_3 ? _field_data_T_40 : _GEN_1745; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1747 = 14'h25 == field_data_lo_3 ? _field_data_T_41 : _GEN_1746; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1748 = 14'h26 == field_data_lo_3 ? _field_data_T_42 : _GEN_1747; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1749 = 14'h27 == field_data_lo_3 ? _field_data_T_43 : _GEN_1748; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1750 = 14'h28 == field_data_lo_3 ? _field_data_T_44 : _GEN_1749; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1751 = 14'h29 == field_data_lo_3 ? _field_data_T_45 : _GEN_1750; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1752 = 14'h2a == field_data_lo_3 ? _field_data_T_46 : _GEN_1751; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1753 = 14'h2b == field_data_lo_3 ? _field_data_T_47 : _GEN_1752; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1754 = 14'h2c == field_data_lo_3 ? _field_data_T_48 : _GEN_1753; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1755 = 14'h2d == field_data_lo_3 ? _field_data_T_49 : _GEN_1754; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1756 = 14'h2e == field_data_lo_3 ? _field_data_T_50 : _GEN_1755; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1757 = 14'h2f == field_data_lo_3 ? _field_data_T_51 : _GEN_1756; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1758 = 14'h30 == field_data_lo_3 ? _field_data_T_52 : _GEN_1757; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1759 = 14'h31 == field_data_lo_3 ? _field_data_T_53 : _GEN_1758; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1760 = 14'h32 == field_data_lo_3 ? _field_data_T_54 : _GEN_1759; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1761 = 14'h33 == field_data_lo_3 ? _field_data_T_55 : _GEN_1760; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1762 = 14'h34 == field_data_lo_3 ? _field_data_T_56 : _GEN_1761; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1763 = 14'h35 == field_data_lo_3 ? _field_data_T_57 : _GEN_1762; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1764 = 14'h36 == field_data_lo_3 ? _field_data_T_58 : _GEN_1763; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1765 = 14'h37 == field_data_lo_3 ? _field_data_T_59 : _GEN_1764; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1766 = 14'h38 == field_data_lo_3 ? _field_data_T_60 : _GEN_1765; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1767 = 14'h39 == field_data_lo_3 ? _field_data_T_61 : _GEN_1766; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1768 = 14'h3a == field_data_lo_3 ? _field_data_T_62 : _GEN_1767; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1769 = 14'h3b == field_data_lo_3 ? _field_data_T_63 : _GEN_1768; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1770 = 14'h3c == field_data_lo_3 ? _field_data_T_64 : _GEN_1769; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1771 = 14'h3d == field_data_lo_3 ? _field_data_T_65 : _GEN_1770; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1772 = 14'h3e == field_data_lo_3 ? _field_data_T_66 : _GEN_1771; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1773 = 14'h3f == field_data_lo_3 ? _field_data_T_67 : _GEN_1772; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1774 = 14'h40 == field_data_lo_3 ? _field_data_T_68 : _GEN_1773; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1775 = 14'h41 == field_data_lo_3 ? _field_data_T_69 : _GEN_1774; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1776 = 14'h42 == field_data_lo_3 ? _field_data_T_70 : _GEN_1775; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1777 = 14'h43 == field_data_lo_3 ? _field_data_T_71 : _GEN_1776; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1778 = 14'h44 == field_data_lo_3 ? _field_data_T_72 : _GEN_1777; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1779 = 14'h45 == field_data_lo_3 ? _field_data_T_73 : _GEN_1778; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1780 = 14'h46 == field_data_lo_3 ? _field_data_T_74 : _GEN_1779; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1781 = 14'h47 == field_data_lo_3 ? _field_data_T_75 : _GEN_1780; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1782 = 14'h48 == field_data_lo_3 ? _field_data_T_76 : _GEN_1781; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1783 = 14'h49 == field_data_lo_3 ? _field_data_T_77 : _GEN_1782; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1784 = 14'h4a == field_data_lo_3 ? _field_data_T_78 : _GEN_1783; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1785 = 14'h4b == field_data_lo_3 ? _field_data_T_79 : _GEN_1784; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1786 = 14'h4c == field_data_lo_3 ? _field_data_T_80 : _GEN_1785; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1787 = 14'h4d == field_data_lo_3 ? _field_data_T_81 : _GEN_1786; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1788 = 14'h4e == field_data_lo_3 ? _field_data_T_82 : _GEN_1787; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1789 = 14'h4f == field_data_lo_3 ? _field_data_T_83 : _GEN_1788; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_36 = vliw_36[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_4 = vliw_36[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_36 = field_data_lo_4[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_36 = field_data_lo_4[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_40 = {{1'd0}, args_offset_36}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_40 = _total_offset_T_40[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1793 = 3'h1 == total_offset_40 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1794 = 3'h2 == total_offset_40 ? args_2 : _GEN_1793; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1795 = 3'h3 == total_offset_40 ? args_3 : _GEN_1794; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1796 = 3'h4 == total_offset_40 ? args_4 : _GEN_1795; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1797 = 3'h5 == total_offset_40 ? args_5 : _GEN_1796; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1798 = 3'h6 == total_offset_40 ? args_6 : _GEN_1797; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1799 = total_offset_40 < 3'h7 ? _GEN_1798 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_36_1 = 3'h0 < args_length_36 ? _GEN_1799 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_41 = args_offset_36 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1802 = 3'h1 == total_offset_41 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1803 = 3'h2 == total_offset_41 ? args_2 : _GEN_1802; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1804 = 3'h3 == total_offset_41 ? args_3 : _GEN_1803; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1805 = 3'h4 == total_offset_41 ? args_4 : _GEN_1804; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1806 = 3'h5 == total_offset_41 ? args_5 : _GEN_1805; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1807 = 3'h6 == total_offset_41 ? args_6 : _GEN_1806; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1808 = total_offset_41 < 3'h7 ? _GEN_1807 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_36_0 = 3'h1 < args_length_36 ? _GEN_1808 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_240 = {field_bytes_36_0,field_bytes_36_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1810 = opcode_36 == 4'ha ? _field_data_T_240 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1811 = opcode_36 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1481 = opcode_36 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_4 = field_data_lo_4[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_243 = {field_data_hi_4,field_data_lo_4}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_73 = _T_1481 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1812 = opcode_36 == 4'h8 | opcode_36 == 4'hb ? _field_data_T_243 : _GEN_1810; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1813 = opcode_36 == 4'h8 | opcode_36 == 4'hb ? _field_tag_T_73 : _GEN_1811; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1814 = 14'h20 == field_data_lo_4 ? _field_data_T_36 : _GEN_1812; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1815 = 14'h21 == field_data_lo_4 ? _field_data_T_37 : _GEN_1814; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1816 = 14'h22 == field_data_lo_4 ? _field_data_T_38 : _GEN_1815; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1817 = 14'h23 == field_data_lo_4 ? _field_data_T_39 : _GEN_1816; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1818 = 14'h24 == field_data_lo_4 ? _field_data_T_40 : _GEN_1817; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1819 = 14'h25 == field_data_lo_4 ? _field_data_T_41 : _GEN_1818; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1820 = 14'h26 == field_data_lo_4 ? _field_data_T_42 : _GEN_1819; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1821 = 14'h27 == field_data_lo_4 ? _field_data_T_43 : _GEN_1820; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1822 = 14'h28 == field_data_lo_4 ? _field_data_T_44 : _GEN_1821; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1823 = 14'h29 == field_data_lo_4 ? _field_data_T_45 : _GEN_1822; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1824 = 14'h2a == field_data_lo_4 ? _field_data_T_46 : _GEN_1823; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1825 = 14'h2b == field_data_lo_4 ? _field_data_T_47 : _GEN_1824; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1826 = 14'h2c == field_data_lo_4 ? _field_data_T_48 : _GEN_1825; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1827 = 14'h2d == field_data_lo_4 ? _field_data_T_49 : _GEN_1826; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1828 = 14'h2e == field_data_lo_4 ? _field_data_T_50 : _GEN_1827; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1829 = 14'h2f == field_data_lo_4 ? _field_data_T_51 : _GEN_1828; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1830 = 14'h30 == field_data_lo_4 ? _field_data_T_52 : _GEN_1829; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1831 = 14'h31 == field_data_lo_4 ? _field_data_T_53 : _GEN_1830; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1832 = 14'h32 == field_data_lo_4 ? _field_data_T_54 : _GEN_1831; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1833 = 14'h33 == field_data_lo_4 ? _field_data_T_55 : _GEN_1832; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1834 = 14'h34 == field_data_lo_4 ? _field_data_T_56 : _GEN_1833; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1835 = 14'h35 == field_data_lo_4 ? _field_data_T_57 : _GEN_1834; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1836 = 14'h36 == field_data_lo_4 ? _field_data_T_58 : _GEN_1835; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1837 = 14'h37 == field_data_lo_4 ? _field_data_T_59 : _GEN_1836; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1838 = 14'h38 == field_data_lo_4 ? _field_data_T_60 : _GEN_1837; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1839 = 14'h39 == field_data_lo_4 ? _field_data_T_61 : _GEN_1838; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1840 = 14'h3a == field_data_lo_4 ? _field_data_T_62 : _GEN_1839; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1841 = 14'h3b == field_data_lo_4 ? _field_data_T_63 : _GEN_1840; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1842 = 14'h3c == field_data_lo_4 ? _field_data_T_64 : _GEN_1841; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1843 = 14'h3d == field_data_lo_4 ? _field_data_T_65 : _GEN_1842; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1844 = 14'h3e == field_data_lo_4 ? _field_data_T_66 : _GEN_1843; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1845 = 14'h3f == field_data_lo_4 ? _field_data_T_67 : _GEN_1844; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1846 = 14'h40 == field_data_lo_4 ? _field_data_T_68 : _GEN_1845; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1847 = 14'h41 == field_data_lo_4 ? _field_data_T_69 : _GEN_1846; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1848 = 14'h42 == field_data_lo_4 ? _field_data_T_70 : _GEN_1847; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1849 = 14'h43 == field_data_lo_4 ? _field_data_T_71 : _GEN_1848; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1850 = 14'h44 == field_data_lo_4 ? _field_data_T_72 : _GEN_1849; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1851 = 14'h45 == field_data_lo_4 ? _field_data_T_73 : _GEN_1850; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1852 = 14'h46 == field_data_lo_4 ? _field_data_T_74 : _GEN_1851; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1853 = 14'h47 == field_data_lo_4 ? _field_data_T_75 : _GEN_1852; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1854 = 14'h48 == field_data_lo_4 ? _field_data_T_76 : _GEN_1853; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1855 = 14'h49 == field_data_lo_4 ? _field_data_T_77 : _GEN_1854; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1856 = 14'h4a == field_data_lo_4 ? _field_data_T_78 : _GEN_1855; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1857 = 14'h4b == field_data_lo_4 ? _field_data_T_79 : _GEN_1856; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1858 = 14'h4c == field_data_lo_4 ? _field_data_T_80 : _GEN_1857; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1859 = 14'h4d == field_data_lo_4 ? _field_data_T_81 : _GEN_1858; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1860 = 14'h4e == field_data_lo_4 ? _field_data_T_82 : _GEN_1859; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1861 = 14'h4f == field_data_lo_4 ? _field_data_T_83 : _GEN_1860; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_37 = vliw_37[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_5 = vliw_37[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_37 = field_data_lo_5[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_37 = field_data_lo_5[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_42 = {{1'd0}, args_offset_37}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_42 = _total_offset_T_42[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1865 = 3'h1 == total_offset_42 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1866 = 3'h2 == total_offset_42 ? args_2 : _GEN_1865; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1867 = 3'h3 == total_offset_42 ? args_3 : _GEN_1866; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1868 = 3'h4 == total_offset_42 ? args_4 : _GEN_1867; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1869 = 3'h5 == total_offset_42 ? args_5 : _GEN_1868; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1870 = 3'h6 == total_offset_42 ? args_6 : _GEN_1869; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1871 = total_offset_42 < 3'h7 ? _GEN_1870 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_37_1 = 3'h0 < args_length_37 ? _GEN_1871 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_43 = args_offset_37 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1874 = 3'h1 == total_offset_43 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1875 = 3'h2 == total_offset_43 ? args_2 : _GEN_1874; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1876 = 3'h3 == total_offset_43 ? args_3 : _GEN_1875; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1877 = 3'h4 == total_offset_43 ? args_4 : _GEN_1876; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1878 = 3'h5 == total_offset_43 ? args_5 : _GEN_1877; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1879 = 3'h6 == total_offset_43 ? args_6 : _GEN_1878; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1880 = total_offset_43 < 3'h7 ? _GEN_1879 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_37_0 = 3'h1 < args_length_37 ? _GEN_1880 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_292 = {field_bytes_37_0,field_bytes_37_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1882 = opcode_37 == 4'ha ? _field_data_T_292 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1883 = opcode_37 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1538 = opcode_37 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_5 = field_data_lo_5[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_295 = {field_data_hi_5,field_data_lo_5}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_75 = _T_1538 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1884 = opcode_37 == 4'h8 | opcode_37 == 4'hb ? _field_data_T_295 : _GEN_1882; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1885 = opcode_37 == 4'h8 | opcode_37 == 4'hb ? _field_tag_T_75 : _GEN_1883; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1886 = 14'h20 == field_data_lo_5 ? _field_data_T_36 : _GEN_1884; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1887 = 14'h21 == field_data_lo_5 ? _field_data_T_37 : _GEN_1886; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1888 = 14'h22 == field_data_lo_5 ? _field_data_T_38 : _GEN_1887; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1889 = 14'h23 == field_data_lo_5 ? _field_data_T_39 : _GEN_1888; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1890 = 14'h24 == field_data_lo_5 ? _field_data_T_40 : _GEN_1889; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1891 = 14'h25 == field_data_lo_5 ? _field_data_T_41 : _GEN_1890; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1892 = 14'h26 == field_data_lo_5 ? _field_data_T_42 : _GEN_1891; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1893 = 14'h27 == field_data_lo_5 ? _field_data_T_43 : _GEN_1892; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1894 = 14'h28 == field_data_lo_5 ? _field_data_T_44 : _GEN_1893; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1895 = 14'h29 == field_data_lo_5 ? _field_data_T_45 : _GEN_1894; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1896 = 14'h2a == field_data_lo_5 ? _field_data_T_46 : _GEN_1895; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1897 = 14'h2b == field_data_lo_5 ? _field_data_T_47 : _GEN_1896; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1898 = 14'h2c == field_data_lo_5 ? _field_data_T_48 : _GEN_1897; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1899 = 14'h2d == field_data_lo_5 ? _field_data_T_49 : _GEN_1898; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1900 = 14'h2e == field_data_lo_5 ? _field_data_T_50 : _GEN_1899; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1901 = 14'h2f == field_data_lo_5 ? _field_data_T_51 : _GEN_1900; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1902 = 14'h30 == field_data_lo_5 ? _field_data_T_52 : _GEN_1901; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1903 = 14'h31 == field_data_lo_5 ? _field_data_T_53 : _GEN_1902; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1904 = 14'h32 == field_data_lo_5 ? _field_data_T_54 : _GEN_1903; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1905 = 14'h33 == field_data_lo_5 ? _field_data_T_55 : _GEN_1904; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1906 = 14'h34 == field_data_lo_5 ? _field_data_T_56 : _GEN_1905; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1907 = 14'h35 == field_data_lo_5 ? _field_data_T_57 : _GEN_1906; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1908 = 14'h36 == field_data_lo_5 ? _field_data_T_58 : _GEN_1907; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1909 = 14'h37 == field_data_lo_5 ? _field_data_T_59 : _GEN_1908; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1910 = 14'h38 == field_data_lo_5 ? _field_data_T_60 : _GEN_1909; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1911 = 14'h39 == field_data_lo_5 ? _field_data_T_61 : _GEN_1910; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1912 = 14'h3a == field_data_lo_5 ? _field_data_T_62 : _GEN_1911; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1913 = 14'h3b == field_data_lo_5 ? _field_data_T_63 : _GEN_1912; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1914 = 14'h3c == field_data_lo_5 ? _field_data_T_64 : _GEN_1913; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1915 = 14'h3d == field_data_lo_5 ? _field_data_T_65 : _GEN_1914; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1916 = 14'h3e == field_data_lo_5 ? _field_data_T_66 : _GEN_1915; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1917 = 14'h3f == field_data_lo_5 ? _field_data_T_67 : _GEN_1916; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1918 = 14'h40 == field_data_lo_5 ? _field_data_T_68 : _GEN_1917; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1919 = 14'h41 == field_data_lo_5 ? _field_data_T_69 : _GEN_1918; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1920 = 14'h42 == field_data_lo_5 ? _field_data_T_70 : _GEN_1919; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1921 = 14'h43 == field_data_lo_5 ? _field_data_T_71 : _GEN_1920; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1922 = 14'h44 == field_data_lo_5 ? _field_data_T_72 : _GEN_1921; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1923 = 14'h45 == field_data_lo_5 ? _field_data_T_73 : _GEN_1922; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1924 = 14'h46 == field_data_lo_5 ? _field_data_T_74 : _GEN_1923; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1925 = 14'h47 == field_data_lo_5 ? _field_data_T_75 : _GEN_1924; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1926 = 14'h48 == field_data_lo_5 ? _field_data_T_76 : _GEN_1925; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1927 = 14'h49 == field_data_lo_5 ? _field_data_T_77 : _GEN_1926; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1928 = 14'h4a == field_data_lo_5 ? _field_data_T_78 : _GEN_1927; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1929 = 14'h4b == field_data_lo_5 ? _field_data_T_79 : _GEN_1928; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1930 = 14'h4c == field_data_lo_5 ? _field_data_T_80 : _GEN_1929; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1931 = 14'h4d == field_data_lo_5 ? _field_data_T_81 : _GEN_1930; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1932 = 14'h4e == field_data_lo_5 ? _field_data_T_82 : _GEN_1931; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1933 = 14'h4f == field_data_lo_5 ? _field_data_T_83 : _GEN_1932; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_38 = vliw_38[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_6 = vliw_38[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_38 = field_data_lo_6[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_38 = field_data_lo_6[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_44 = {{1'd0}, args_offset_38}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_44 = _total_offset_T_44[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1937 = 3'h1 == total_offset_44 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1938 = 3'h2 == total_offset_44 ? args_2 : _GEN_1937; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1939 = 3'h3 == total_offset_44 ? args_3 : _GEN_1938; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1940 = 3'h4 == total_offset_44 ? args_4 : _GEN_1939; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1941 = 3'h5 == total_offset_44 ? args_5 : _GEN_1940; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1942 = 3'h6 == total_offset_44 ? args_6 : _GEN_1941; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1943 = total_offset_44 < 3'h7 ? _GEN_1942 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_38_1 = 3'h0 < args_length_38 ? _GEN_1943 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_45 = args_offset_38 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1946 = 3'h1 == total_offset_45 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1947 = 3'h2 == total_offset_45 ? args_2 : _GEN_1946; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1948 = 3'h3 == total_offset_45 ? args_3 : _GEN_1947; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1949 = 3'h4 == total_offset_45 ? args_4 : _GEN_1948; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1950 = 3'h5 == total_offset_45 ? args_5 : _GEN_1949; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1951 = 3'h6 == total_offset_45 ? args_6 : _GEN_1950; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1952 = total_offset_45 < 3'h7 ? _GEN_1951 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_38_0 = 3'h1 < args_length_38 ? _GEN_1952 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_344 = {field_bytes_38_0,field_bytes_38_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1954 = opcode_38 == 4'ha ? _field_data_T_344 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1955 = opcode_38 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1595 = opcode_38 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_6 = field_data_lo_6[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_347 = {field_data_hi_6,field_data_lo_6}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_77 = _T_1595 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1956 = opcode_38 == 4'h8 | opcode_38 == 4'hb ? _field_data_T_347 : _GEN_1954; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1957 = opcode_38 == 4'h8 | opcode_38 == 4'hb ? _field_tag_T_77 : _GEN_1955; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1958 = 14'h20 == field_data_lo_6 ? _field_data_T_36 : _GEN_1956; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1959 = 14'h21 == field_data_lo_6 ? _field_data_T_37 : _GEN_1958; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1960 = 14'h22 == field_data_lo_6 ? _field_data_T_38 : _GEN_1959; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1961 = 14'h23 == field_data_lo_6 ? _field_data_T_39 : _GEN_1960; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1962 = 14'h24 == field_data_lo_6 ? _field_data_T_40 : _GEN_1961; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1963 = 14'h25 == field_data_lo_6 ? _field_data_T_41 : _GEN_1962; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1964 = 14'h26 == field_data_lo_6 ? _field_data_T_42 : _GEN_1963; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1965 = 14'h27 == field_data_lo_6 ? _field_data_T_43 : _GEN_1964; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1966 = 14'h28 == field_data_lo_6 ? _field_data_T_44 : _GEN_1965; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1967 = 14'h29 == field_data_lo_6 ? _field_data_T_45 : _GEN_1966; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1968 = 14'h2a == field_data_lo_6 ? _field_data_T_46 : _GEN_1967; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1969 = 14'h2b == field_data_lo_6 ? _field_data_T_47 : _GEN_1968; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1970 = 14'h2c == field_data_lo_6 ? _field_data_T_48 : _GEN_1969; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1971 = 14'h2d == field_data_lo_6 ? _field_data_T_49 : _GEN_1970; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1972 = 14'h2e == field_data_lo_6 ? _field_data_T_50 : _GEN_1971; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1973 = 14'h2f == field_data_lo_6 ? _field_data_T_51 : _GEN_1972; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1974 = 14'h30 == field_data_lo_6 ? _field_data_T_52 : _GEN_1973; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1975 = 14'h31 == field_data_lo_6 ? _field_data_T_53 : _GEN_1974; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1976 = 14'h32 == field_data_lo_6 ? _field_data_T_54 : _GEN_1975; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1977 = 14'h33 == field_data_lo_6 ? _field_data_T_55 : _GEN_1976; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1978 = 14'h34 == field_data_lo_6 ? _field_data_T_56 : _GEN_1977; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1979 = 14'h35 == field_data_lo_6 ? _field_data_T_57 : _GEN_1978; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1980 = 14'h36 == field_data_lo_6 ? _field_data_T_58 : _GEN_1979; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1981 = 14'h37 == field_data_lo_6 ? _field_data_T_59 : _GEN_1980; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1982 = 14'h38 == field_data_lo_6 ? _field_data_T_60 : _GEN_1981; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1983 = 14'h39 == field_data_lo_6 ? _field_data_T_61 : _GEN_1982; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1984 = 14'h3a == field_data_lo_6 ? _field_data_T_62 : _GEN_1983; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1985 = 14'h3b == field_data_lo_6 ? _field_data_T_63 : _GEN_1984; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1986 = 14'h3c == field_data_lo_6 ? _field_data_T_64 : _GEN_1985; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1987 = 14'h3d == field_data_lo_6 ? _field_data_T_65 : _GEN_1986; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1988 = 14'h3e == field_data_lo_6 ? _field_data_T_66 : _GEN_1987; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1989 = 14'h3f == field_data_lo_6 ? _field_data_T_67 : _GEN_1988; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1990 = 14'h40 == field_data_lo_6 ? _field_data_T_68 : _GEN_1989; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1991 = 14'h41 == field_data_lo_6 ? _field_data_T_69 : _GEN_1990; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1992 = 14'h42 == field_data_lo_6 ? _field_data_T_70 : _GEN_1991; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1993 = 14'h43 == field_data_lo_6 ? _field_data_T_71 : _GEN_1992; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1994 = 14'h44 == field_data_lo_6 ? _field_data_T_72 : _GEN_1993; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1995 = 14'h45 == field_data_lo_6 ? _field_data_T_73 : _GEN_1994; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1996 = 14'h46 == field_data_lo_6 ? _field_data_T_74 : _GEN_1995; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1997 = 14'h47 == field_data_lo_6 ? _field_data_T_75 : _GEN_1996; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1998 = 14'h48 == field_data_lo_6 ? _field_data_T_76 : _GEN_1997; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1999 = 14'h49 == field_data_lo_6 ? _field_data_T_77 : _GEN_1998; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2000 = 14'h4a == field_data_lo_6 ? _field_data_T_78 : _GEN_1999; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2001 = 14'h4b == field_data_lo_6 ? _field_data_T_79 : _GEN_2000; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2002 = 14'h4c == field_data_lo_6 ? _field_data_T_80 : _GEN_2001; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2003 = 14'h4d == field_data_lo_6 ? _field_data_T_81 : _GEN_2002; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2004 = 14'h4e == field_data_lo_6 ? _field_data_T_82 : _GEN_2003; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2005 = 14'h4f == field_data_lo_6 ? _field_data_T_83 : _GEN_2004; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_39 = vliw_39[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_7 = vliw_39[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_39 = field_data_lo_7[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_39 = field_data_lo_7[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_46 = {{1'd0}, args_offset_39}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_46 = _total_offset_T_46[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2009 = 3'h1 == total_offset_46 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2010 = 3'h2 == total_offset_46 ? args_2 : _GEN_2009; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2011 = 3'h3 == total_offset_46 ? args_3 : _GEN_2010; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2012 = 3'h4 == total_offset_46 ? args_4 : _GEN_2011; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2013 = 3'h5 == total_offset_46 ? args_5 : _GEN_2012; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2014 = 3'h6 == total_offset_46 ? args_6 : _GEN_2013; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2015 = total_offset_46 < 3'h7 ? _GEN_2014 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_39_1 = 3'h0 < args_length_39 ? _GEN_2015 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_47 = args_offset_39 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2018 = 3'h1 == total_offset_47 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2019 = 3'h2 == total_offset_47 ? args_2 : _GEN_2018; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2020 = 3'h3 == total_offset_47 ? args_3 : _GEN_2019; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2021 = 3'h4 == total_offset_47 ? args_4 : _GEN_2020; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2022 = 3'h5 == total_offset_47 ? args_5 : _GEN_2021; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2023 = 3'h6 == total_offset_47 ? args_6 : _GEN_2022; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2024 = total_offset_47 < 3'h7 ? _GEN_2023 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_39_0 = 3'h1 < args_length_39 ? _GEN_2024 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_396 = {field_bytes_39_0,field_bytes_39_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2026 = opcode_39 == 4'ha ? _field_data_T_396 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2027 = opcode_39 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1652 = opcode_39 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_7 = field_data_lo_7[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_399 = {field_data_hi_7,field_data_lo_7}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_79 = _T_1652 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2028 = opcode_39 == 4'h8 | opcode_39 == 4'hb ? _field_data_T_399 : _GEN_2026; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2029 = opcode_39 == 4'h8 | opcode_39 == 4'hb ? _field_tag_T_79 : _GEN_2027; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2030 = 14'h20 == field_data_lo_7 ? _field_data_T_36 : _GEN_2028; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2031 = 14'h21 == field_data_lo_7 ? _field_data_T_37 : _GEN_2030; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2032 = 14'h22 == field_data_lo_7 ? _field_data_T_38 : _GEN_2031; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2033 = 14'h23 == field_data_lo_7 ? _field_data_T_39 : _GEN_2032; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2034 = 14'h24 == field_data_lo_7 ? _field_data_T_40 : _GEN_2033; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2035 = 14'h25 == field_data_lo_7 ? _field_data_T_41 : _GEN_2034; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2036 = 14'h26 == field_data_lo_7 ? _field_data_T_42 : _GEN_2035; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2037 = 14'h27 == field_data_lo_7 ? _field_data_T_43 : _GEN_2036; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2038 = 14'h28 == field_data_lo_7 ? _field_data_T_44 : _GEN_2037; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2039 = 14'h29 == field_data_lo_7 ? _field_data_T_45 : _GEN_2038; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2040 = 14'h2a == field_data_lo_7 ? _field_data_T_46 : _GEN_2039; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2041 = 14'h2b == field_data_lo_7 ? _field_data_T_47 : _GEN_2040; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2042 = 14'h2c == field_data_lo_7 ? _field_data_T_48 : _GEN_2041; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2043 = 14'h2d == field_data_lo_7 ? _field_data_T_49 : _GEN_2042; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2044 = 14'h2e == field_data_lo_7 ? _field_data_T_50 : _GEN_2043; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2045 = 14'h2f == field_data_lo_7 ? _field_data_T_51 : _GEN_2044; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2046 = 14'h30 == field_data_lo_7 ? _field_data_T_52 : _GEN_2045; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2047 = 14'h31 == field_data_lo_7 ? _field_data_T_53 : _GEN_2046; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2048 = 14'h32 == field_data_lo_7 ? _field_data_T_54 : _GEN_2047; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2049 = 14'h33 == field_data_lo_7 ? _field_data_T_55 : _GEN_2048; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2050 = 14'h34 == field_data_lo_7 ? _field_data_T_56 : _GEN_2049; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2051 = 14'h35 == field_data_lo_7 ? _field_data_T_57 : _GEN_2050; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2052 = 14'h36 == field_data_lo_7 ? _field_data_T_58 : _GEN_2051; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2053 = 14'h37 == field_data_lo_7 ? _field_data_T_59 : _GEN_2052; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2054 = 14'h38 == field_data_lo_7 ? _field_data_T_60 : _GEN_2053; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2055 = 14'h39 == field_data_lo_7 ? _field_data_T_61 : _GEN_2054; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2056 = 14'h3a == field_data_lo_7 ? _field_data_T_62 : _GEN_2055; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2057 = 14'h3b == field_data_lo_7 ? _field_data_T_63 : _GEN_2056; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2058 = 14'h3c == field_data_lo_7 ? _field_data_T_64 : _GEN_2057; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2059 = 14'h3d == field_data_lo_7 ? _field_data_T_65 : _GEN_2058; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2060 = 14'h3e == field_data_lo_7 ? _field_data_T_66 : _GEN_2059; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2061 = 14'h3f == field_data_lo_7 ? _field_data_T_67 : _GEN_2060; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2062 = 14'h40 == field_data_lo_7 ? _field_data_T_68 : _GEN_2061; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2063 = 14'h41 == field_data_lo_7 ? _field_data_T_69 : _GEN_2062; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2064 = 14'h42 == field_data_lo_7 ? _field_data_T_70 : _GEN_2063; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2065 = 14'h43 == field_data_lo_7 ? _field_data_T_71 : _GEN_2064; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2066 = 14'h44 == field_data_lo_7 ? _field_data_T_72 : _GEN_2065; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2067 = 14'h45 == field_data_lo_7 ? _field_data_T_73 : _GEN_2066; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2068 = 14'h46 == field_data_lo_7 ? _field_data_T_74 : _GEN_2067; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2069 = 14'h47 == field_data_lo_7 ? _field_data_T_75 : _GEN_2068; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2070 = 14'h48 == field_data_lo_7 ? _field_data_T_76 : _GEN_2069; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2071 = 14'h49 == field_data_lo_7 ? _field_data_T_77 : _GEN_2070; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2072 = 14'h4a == field_data_lo_7 ? _field_data_T_78 : _GEN_2071; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2073 = 14'h4b == field_data_lo_7 ? _field_data_T_79 : _GEN_2072; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2074 = 14'h4c == field_data_lo_7 ? _field_data_T_80 : _GEN_2073; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2075 = 14'h4d == field_data_lo_7 ? _field_data_T_81 : _GEN_2074; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2076 = 14'h4e == field_data_lo_7 ? _field_data_T_82 : _GEN_2075; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2077 = 14'h4f == field_data_lo_7 ? _field_data_T_83 : _GEN_2076; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_40 = vliw_40[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_8 = vliw_40[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_40 = field_data_lo_8[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_40 = field_data_lo_8[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_48 = {{1'd0}, args_offset_40}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_48 = _total_offset_T_48[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2081 = 3'h1 == total_offset_48 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2082 = 3'h2 == total_offset_48 ? args_2 : _GEN_2081; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2083 = 3'h3 == total_offset_48 ? args_3 : _GEN_2082; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2084 = 3'h4 == total_offset_48 ? args_4 : _GEN_2083; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2085 = 3'h5 == total_offset_48 ? args_5 : _GEN_2084; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2086 = 3'h6 == total_offset_48 ? args_6 : _GEN_2085; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2087 = total_offset_48 < 3'h7 ? _GEN_2086 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_40_1 = 3'h0 < args_length_40 ? _GEN_2087 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_49 = args_offset_40 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2090 = 3'h1 == total_offset_49 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2091 = 3'h2 == total_offset_49 ? args_2 : _GEN_2090; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2092 = 3'h3 == total_offset_49 ? args_3 : _GEN_2091; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2093 = 3'h4 == total_offset_49 ? args_4 : _GEN_2092; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2094 = 3'h5 == total_offset_49 ? args_5 : _GEN_2093; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2095 = 3'h6 == total_offset_49 ? args_6 : _GEN_2094; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2096 = total_offset_49 < 3'h7 ? _GEN_2095 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_40_0 = 3'h1 < args_length_40 ? _GEN_2096 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_448 = {field_bytes_40_0,field_bytes_40_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2098 = opcode_40 == 4'ha ? _field_data_T_448 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2099 = opcode_40 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1709 = opcode_40 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_8 = field_data_lo_8[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_451 = {field_data_hi_8,field_data_lo_8}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_81 = _T_1709 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2100 = opcode_40 == 4'h8 | opcode_40 == 4'hb ? _field_data_T_451 : _GEN_2098; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2101 = opcode_40 == 4'h8 | opcode_40 == 4'hb ? _field_tag_T_81 : _GEN_2099; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2102 = 14'h20 == field_data_lo_8 ? _field_data_T_36 : _GEN_2100; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2103 = 14'h21 == field_data_lo_8 ? _field_data_T_37 : _GEN_2102; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2104 = 14'h22 == field_data_lo_8 ? _field_data_T_38 : _GEN_2103; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2105 = 14'h23 == field_data_lo_8 ? _field_data_T_39 : _GEN_2104; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2106 = 14'h24 == field_data_lo_8 ? _field_data_T_40 : _GEN_2105; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2107 = 14'h25 == field_data_lo_8 ? _field_data_T_41 : _GEN_2106; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2108 = 14'h26 == field_data_lo_8 ? _field_data_T_42 : _GEN_2107; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2109 = 14'h27 == field_data_lo_8 ? _field_data_T_43 : _GEN_2108; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2110 = 14'h28 == field_data_lo_8 ? _field_data_T_44 : _GEN_2109; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2111 = 14'h29 == field_data_lo_8 ? _field_data_T_45 : _GEN_2110; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2112 = 14'h2a == field_data_lo_8 ? _field_data_T_46 : _GEN_2111; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2113 = 14'h2b == field_data_lo_8 ? _field_data_T_47 : _GEN_2112; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2114 = 14'h2c == field_data_lo_8 ? _field_data_T_48 : _GEN_2113; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2115 = 14'h2d == field_data_lo_8 ? _field_data_T_49 : _GEN_2114; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2116 = 14'h2e == field_data_lo_8 ? _field_data_T_50 : _GEN_2115; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2117 = 14'h2f == field_data_lo_8 ? _field_data_T_51 : _GEN_2116; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2118 = 14'h30 == field_data_lo_8 ? _field_data_T_52 : _GEN_2117; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2119 = 14'h31 == field_data_lo_8 ? _field_data_T_53 : _GEN_2118; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2120 = 14'h32 == field_data_lo_8 ? _field_data_T_54 : _GEN_2119; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2121 = 14'h33 == field_data_lo_8 ? _field_data_T_55 : _GEN_2120; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2122 = 14'h34 == field_data_lo_8 ? _field_data_T_56 : _GEN_2121; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2123 = 14'h35 == field_data_lo_8 ? _field_data_T_57 : _GEN_2122; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2124 = 14'h36 == field_data_lo_8 ? _field_data_T_58 : _GEN_2123; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2125 = 14'h37 == field_data_lo_8 ? _field_data_T_59 : _GEN_2124; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2126 = 14'h38 == field_data_lo_8 ? _field_data_T_60 : _GEN_2125; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2127 = 14'h39 == field_data_lo_8 ? _field_data_T_61 : _GEN_2126; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2128 = 14'h3a == field_data_lo_8 ? _field_data_T_62 : _GEN_2127; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2129 = 14'h3b == field_data_lo_8 ? _field_data_T_63 : _GEN_2128; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2130 = 14'h3c == field_data_lo_8 ? _field_data_T_64 : _GEN_2129; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2131 = 14'h3d == field_data_lo_8 ? _field_data_T_65 : _GEN_2130; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2132 = 14'h3e == field_data_lo_8 ? _field_data_T_66 : _GEN_2131; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2133 = 14'h3f == field_data_lo_8 ? _field_data_T_67 : _GEN_2132; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2134 = 14'h40 == field_data_lo_8 ? _field_data_T_68 : _GEN_2133; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2135 = 14'h41 == field_data_lo_8 ? _field_data_T_69 : _GEN_2134; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2136 = 14'h42 == field_data_lo_8 ? _field_data_T_70 : _GEN_2135; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2137 = 14'h43 == field_data_lo_8 ? _field_data_T_71 : _GEN_2136; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2138 = 14'h44 == field_data_lo_8 ? _field_data_T_72 : _GEN_2137; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2139 = 14'h45 == field_data_lo_8 ? _field_data_T_73 : _GEN_2138; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2140 = 14'h46 == field_data_lo_8 ? _field_data_T_74 : _GEN_2139; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2141 = 14'h47 == field_data_lo_8 ? _field_data_T_75 : _GEN_2140; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2142 = 14'h48 == field_data_lo_8 ? _field_data_T_76 : _GEN_2141; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2143 = 14'h49 == field_data_lo_8 ? _field_data_T_77 : _GEN_2142; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2144 = 14'h4a == field_data_lo_8 ? _field_data_T_78 : _GEN_2143; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2145 = 14'h4b == field_data_lo_8 ? _field_data_T_79 : _GEN_2144; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2146 = 14'h4c == field_data_lo_8 ? _field_data_T_80 : _GEN_2145; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2147 = 14'h4d == field_data_lo_8 ? _field_data_T_81 : _GEN_2146; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2148 = 14'h4e == field_data_lo_8 ? _field_data_T_82 : _GEN_2147; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2149 = 14'h4f == field_data_lo_8 ? _field_data_T_83 : _GEN_2148; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_41 = vliw_41[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_9 = vliw_41[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_41 = field_data_lo_9[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_41 = field_data_lo_9[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_50 = {{1'd0}, args_offset_41}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_50 = _total_offset_T_50[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2153 = 3'h1 == total_offset_50 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2154 = 3'h2 == total_offset_50 ? args_2 : _GEN_2153; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2155 = 3'h3 == total_offset_50 ? args_3 : _GEN_2154; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2156 = 3'h4 == total_offset_50 ? args_4 : _GEN_2155; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2157 = 3'h5 == total_offset_50 ? args_5 : _GEN_2156; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2158 = 3'h6 == total_offset_50 ? args_6 : _GEN_2157; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2159 = total_offset_50 < 3'h7 ? _GEN_2158 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_41_1 = 3'h0 < args_length_41 ? _GEN_2159 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_51 = args_offset_41 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2162 = 3'h1 == total_offset_51 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2163 = 3'h2 == total_offset_51 ? args_2 : _GEN_2162; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2164 = 3'h3 == total_offset_51 ? args_3 : _GEN_2163; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2165 = 3'h4 == total_offset_51 ? args_4 : _GEN_2164; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2166 = 3'h5 == total_offset_51 ? args_5 : _GEN_2165; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2167 = 3'h6 == total_offset_51 ? args_6 : _GEN_2166; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2168 = total_offset_51 < 3'h7 ? _GEN_2167 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_41_0 = 3'h1 < args_length_41 ? _GEN_2168 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_500 = {field_bytes_41_0,field_bytes_41_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2170 = opcode_41 == 4'ha ? _field_data_T_500 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2171 = opcode_41 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1766 = opcode_41 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_9 = field_data_lo_9[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_503 = {field_data_hi_9,field_data_lo_9}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_83 = _T_1766 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2172 = opcode_41 == 4'h8 | opcode_41 == 4'hb ? _field_data_T_503 : _GEN_2170; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2173 = opcode_41 == 4'h8 | opcode_41 == 4'hb ? _field_tag_T_83 : _GEN_2171; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2174 = 14'h20 == field_data_lo_9 ? _field_data_T_36 : _GEN_2172; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2175 = 14'h21 == field_data_lo_9 ? _field_data_T_37 : _GEN_2174; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2176 = 14'h22 == field_data_lo_9 ? _field_data_T_38 : _GEN_2175; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2177 = 14'h23 == field_data_lo_9 ? _field_data_T_39 : _GEN_2176; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2178 = 14'h24 == field_data_lo_9 ? _field_data_T_40 : _GEN_2177; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2179 = 14'h25 == field_data_lo_9 ? _field_data_T_41 : _GEN_2178; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2180 = 14'h26 == field_data_lo_9 ? _field_data_T_42 : _GEN_2179; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2181 = 14'h27 == field_data_lo_9 ? _field_data_T_43 : _GEN_2180; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2182 = 14'h28 == field_data_lo_9 ? _field_data_T_44 : _GEN_2181; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2183 = 14'h29 == field_data_lo_9 ? _field_data_T_45 : _GEN_2182; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2184 = 14'h2a == field_data_lo_9 ? _field_data_T_46 : _GEN_2183; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2185 = 14'h2b == field_data_lo_9 ? _field_data_T_47 : _GEN_2184; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2186 = 14'h2c == field_data_lo_9 ? _field_data_T_48 : _GEN_2185; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2187 = 14'h2d == field_data_lo_9 ? _field_data_T_49 : _GEN_2186; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2188 = 14'h2e == field_data_lo_9 ? _field_data_T_50 : _GEN_2187; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2189 = 14'h2f == field_data_lo_9 ? _field_data_T_51 : _GEN_2188; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2190 = 14'h30 == field_data_lo_9 ? _field_data_T_52 : _GEN_2189; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2191 = 14'h31 == field_data_lo_9 ? _field_data_T_53 : _GEN_2190; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2192 = 14'h32 == field_data_lo_9 ? _field_data_T_54 : _GEN_2191; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2193 = 14'h33 == field_data_lo_9 ? _field_data_T_55 : _GEN_2192; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2194 = 14'h34 == field_data_lo_9 ? _field_data_T_56 : _GEN_2193; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2195 = 14'h35 == field_data_lo_9 ? _field_data_T_57 : _GEN_2194; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2196 = 14'h36 == field_data_lo_9 ? _field_data_T_58 : _GEN_2195; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2197 = 14'h37 == field_data_lo_9 ? _field_data_T_59 : _GEN_2196; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2198 = 14'h38 == field_data_lo_9 ? _field_data_T_60 : _GEN_2197; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2199 = 14'h39 == field_data_lo_9 ? _field_data_T_61 : _GEN_2198; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2200 = 14'h3a == field_data_lo_9 ? _field_data_T_62 : _GEN_2199; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2201 = 14'h3b == field_data_lo_9 ? _field_data_T_63 : _GEN_2200; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2202 = 14'h3c == field_data_lo_9 ? _field_data_T_64 : _GEN_2201; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2203 = 14'h3d == field_data_lo_9 ? _field_data_T_65 : _GEN_2202; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2204 = 14'h3e == field_data_lo_9 ? _field_data_T_66 : _GEN_2203; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2205 = 14'h3f == field_data_lo_9 ? _field_data_T_67 : _GEN_2204; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2206 = 14'h40 == field_data_lo_9 ? _field_data_T_68 : _GEN_2205; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2207 = 14'h41 == field_data_lo_9 ? _field_data_T_69 : _GEN_2206; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2208 = 14'h42 == field_data_lo_9 ? _field_data_T_70 : _GEN_2207; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2209 = 14'h43 == field_data_lo_9 ? _field_data_T_71 : _GEN_2208; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2210 = 14'h44 == field_data_lo_9 ? _field_data_T_72 : _GEN_2209; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2211 = 14'h45 == field_data_lo_9 ? _field_data_T_73 : _GEN_2210; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2212 = 14'h46 == field_data_lo_9 ? _field_data_T_74 : _GEN_2211; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2213 = 14'h47 == field_data_lo_9 ? _field_data_T_75 : _GEN_2212; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2214 = 14'h48 == field_data_lo_9 ? _field_data_T_76 : _GEN_2213; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2215 = 14'h49 == field_data_lo_9 ? _field_data_T_77 : _GEN_2214; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2216 = 14'h4a == field_data_lo_9 ? _field_data_T_78 : _GEN_2215; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2217 = 14'h4b == field_data_lo_9 ? _field_data_T_79 : _GEN_2216; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2218 = 14'h4c == field_data_lo_9 ? _field_data_T_80 : _GEN_2217; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2219 = 14'h4d == field_data_lo_9 ? _field_data_T_81 : _GEN_2218; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2220 = 14'h4e == field_data_lo_9 ? _field_data_T_82 : _GEN_2219; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2221 = 14'h4f == field_data_lo_9 ? _field_data_T_83 : _GEN_2220; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_42 = vliw_42[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_10 = vliw_42[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_42 = field_data_lo_10[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_42 = field_data_lo_10[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_52 = {{1'd0}, args_offset_42}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_52 = _total_offset_T_52[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2225 = 3'h1 == total_offset_52 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2226 = 3'h2 == total_offset_52 ? args_2 : _GEN_2225; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2227 = 3'h3 == total_offset_52 ? args_3 : _GEN_2226; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2228 = 3'h4 == total_offset_52 ? args_4 : _GEN_2227; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2229 = 3'h5 == total_offset_52 ? args_5 : _GEN_2228; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2230 = 3'h6 == total_offset_52 ? args_6 : _GEN_2229; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2231 = total_offset_52 < 3'h7 ? _GEN_2230 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_42_1 = 3'h0 < args_length_42 ? _GEN_2231 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_53 = args_offset_42 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2234 = 3'h1 == total_offset_53 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2235 = 3'h2 == total_offset_53 ? args_2 : _GEN_2234; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2236 = 3'h3 == total_offset_53 ? args_3 : _GEN_2235; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2237 = 3'h4 == total_offset_53 ? args_4 : _GEN_2236; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2238 = 3'h5 == total_offset_53 ? args_5 : _GEN_2237; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2239 = 3'h6 == total_offset_53 ? args_6 : _GEN_2238; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2240 = total_offset_53 < 3'h7 ? _GEN_2239 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_42_0 = 3'h1 < args_length_42 ? _GEN_2240 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_552 = {field_bytes_42_0,field_bytes_42_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2242 = opcode_42 == 4'ha ? _field_data_T_552 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2243 = opcode_42 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1823 = opcode_42 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_10 = field_data_lo_10[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_555 = {field_data_hi_10,field_data_lo_10}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_85 = _T_1823 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2244 = opcode_42 == 4'h8 | opcode_42 == 4'hb ? _field_data_T_555 : _GEN_2242; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2245 = opcode_42 == 4'h8 | opcode_42 == 4'hb ? _field_tag_T_85 : _GEN_2243; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2246 = 14'h20 == field_data_lo_10 ? _field_data_T_36 : _GEN_2244; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2247 = 14'h21 == field_data_lo_10 ? _field_data_T_37 : _GEN_2246; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2248 = 14'h22 == field_data_lo_10 ? _field_data_T_38 : _GEN_2247; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2249 = 14'h23 == field_data_lo_10 ? _field_data_T_39 : _GEN_2248; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2250 = 14'h24 == field_data_lo_10 ? _field_data_T_40 : _GEN_2249; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2251 = 14'h25 == field_data_lo_10 ? _field_data_T_41 : _GEN_2250; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2252 = 14'h26 == field_data_lo_10 ? _field_data_T_42 : _GEN_2251; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2253 = 14'h27 == field_data_lo_10 ? _field_data_T_43 : _GEN_2252; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2254 = 14'h28 == field_data_lo_10 ? _field_data_T_44 : _GEN_2253; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2255 = 14'h29 == field_data_lo_10 ? _field_data_T_45 : _GEN_2254; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2256 = 14'h2a == field_data_lo_10 ? _field_data_T_46 : _GEN_2255; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2257 = 14'h2b == field_data_lo_10 ? _field_data_T_47 : _GEN_2256; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2258 = 14'h2c == field_data_lo_10 ? _field_data_T_48 : _GEN_2257; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2259 = 14'h2d == field_data_lo_10 ? _field_data_T_49 : _GEN_2258; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2260 = 14'h2e == field_data_lo_10 ? _field_data_T_50 : _GEN_2259; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2261 = 14'h2f == field_data_lo_10 ? _field_data_T_51 : _GEN_2260; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2262 = 14'h30 == field_data_lo_10 ? _field_data_T_52 : _GEN_2261; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2263 = 14'h31 == field_data_lo_10 ? _field_data_T_53 : _GEN_2262; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2264 = 14'h32 == field_data_lo_10 ? _field_data_T_54 : _GEN_2263; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2265 = 14'h33 == field_data_lo_10 ? _field_data_T_55 : _GEN_2264; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2266 = 14'h34 == field_data_lo_10 ? _field_data_T_56 : _GEN_2265; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2267 = 14'h35 == field_data_lo_10 ? _field_data_T_57 : _GEN_2266; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2268 = 14'h36 == field_data_lo_10 ? _field_data_T_58 : _GEN_2267; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2269 = 14'h37 == field_data_lo_10 ? _field_data_T_59 : _GEN_2268; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2270 = 14'h38 == field_data_lo_10 ? _field_data_T_60 : _GEN_2269; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2271 = 14'h39 == field_data_lo_10 ? _field_data_T_61 : _GEN_2270; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2272 = 14'h3a == field_data_lo_10 ? _field_data_T_62 : _GEN_2271; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2273 = 14'h3b == field_data_lo_10 ? _field_data_T_63 : _GEN_2272; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2274 = 14'h3c == field_data_lo_10 ? _field_data_T_64 : _GEN_2273; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2275 = 14'h3d == field_data_lo_10 ? _field_data_T_65 : _GEN_2274; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2276 = 14'h3e == field_data_lo_10 ? _field_data_T_66 : _GEN_2275; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2277 = 14'h3f == field_data_lo_10 ? _field_data_T_67 : _GEN_2276; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2278 = 14'h40 == field_data_lo_10 ? _field_data_T_68 : _GEN_2277; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2279 = 14'h41 == field_data_lo_10 ? _field_data_T_69 : _GEN_2278; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2280 = 14'h42 == field_data_lo_10 ? _field_data_T_70 : _GEN_2279; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2281 = 14'h43 == field_data_lo_10 ? _field_data_T_71 : _GEN_2280; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2282 = 14'h44 == field_data_lo_10 ? _field_data_T_72 : _GEN_2281; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2283 = 14'h45 == field_data_lo_10 ? _field_data_T_73 : _GEN_2282; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2284 = 14'h46 == field_data_lo_10 ? _field_data_T_74 : _GEN_2283; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2285 = 14'h47 == field_data_lo_10 ? _field_data_T_75 : _GEN_2284; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2286 = 14'h48 == field_data_lo_10 ? _field_data_T_76 : _GEN_2285; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2287 = 14'h49 == field_data_lo_10 ? _field_data_T_77 : _GEN_2286; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2288 = 14'h4a == field_data_lo_10 ? _field_data_T_78 : _GEN_2287; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2289 = 14'h4b == field_data_lo_10 ? _field_data_T_79 : _GEN_2288; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2290 = 14'h4c == field_data_lo_10 ? _field_data_T_80 : _GEN_2289; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2291 = 14'h4d == field_data_lo_10 ? _field_data_T_81 : _GEN_2290; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2292 = 14'h4e == field_data_lo_10 ? _field_data_T_82 : _GEN_2291; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2293 = 14'h4f == field_data_lo_10 ? _field_data_T_83 : _GEN_2292; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_43 = vliw_43[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_11 = vliw_43[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_43 = field_data_lo_11[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_43 = field_data_lo_11[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_54 = {{1'd0}, args_offset_43}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_54 = _total_offset_T_54[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2297 = 3'h1 == total_offset_54 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2298 = 3'h2 == total_offset_54 ? args_2 : _GEN_2297; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2299 = 3'h3 == total_offset_54 ? args_3 : _GEN_2298; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2300 = 3'h4 == total_offset_54 ? args_4 : _GEN_2299; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2301 = 3'h5 == total_offset_54 ? args_5 : _GEN_2300; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2302 = 3'h6 == total_offset_54 ? args_6 : _GEN_2301; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2303 = total_offset_54 < 3'h7 ? _GEN_2302 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_43_1 = 3'h0 < args_length_43 ? _GEN_2303 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_55 = args_offset_43 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2306 = 3'h1 == total_offset_55 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2307 = 3'h2 == total_offset_55 ? args_2 : _GEN_2306; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2308 = 3'h3 == total_offset_55 ? args_3 : _GEN_2307; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2309 = 3'h4 == total_offset_55 ? args_4 : _GEN_2308; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2310 = 3'h5 == total_offset_55 ? args_5 : _GEN_2309; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2311 = 3'h6 == total_offset_55 ? args_6 : _GEN_2310; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2312 = total_offset_55 < 3'h7 ? _GEN_2311 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_43_0 = 3'h1 < args_length_43 ? _GEN_2312 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_604 = {field_bytes_43_0,field_bytes_43_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2314 = opcode_43 == 4'ha ? _field_data_T_604 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2315 = opcode_43 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1880 = opcode_43 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_11 = field_data_lo_11[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_607 = {field_data_hi_11,field_data_lo_11}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_87 = _T_1880 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2316 = opcode_43 == 4'h8 | opcode_43 == 4'hb ? _field_data_T_607 : _GEN_2314; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2317 = opcode_43 == 4'h8 | opcode_43 == 4'hb ? _field_tag_T_87 : _GEN_2315; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2318 = 14'h20 == field_data_lo_11 ? _field_data_T_36 : _GEN_2316; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2319 = 14'h21 == field_data_lo_11 ? _field_data_T_37 : _GEN_2318; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2320 = 14'h22 == field_data_lo_11 ? _field_data_T_38 : _GEN_2319; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2321 = 14'h23 == field_data_lo_11 ? _field_data_T_39 : _GEN_2320; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2322 = 14'h24 == field_data_lo_11 ? _field_data_T_40 : _GEN_2321; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2323 = 14'h25 == field_data_lo_11 ? _field_data_T_41 : _GEN_2322; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2324 = 14'h26 == field_data_lo_11 ? _field_data_T_42 : _GEN_2323; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2325 = 14'h27 == field_data_lo_11 ? _field_data_T_43 : _GEN_2324; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2326 = 14'h28 == field_data_lo_11 ? _field_data_T_44 : _GEN_2325; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2327 = 14'h29 == field_data_lo_11 ? _field_data_T_45 : _GEN_2326; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2328 = 14'h2a == field_data_lo_11 ? _field_data_T_46 : _GEN_2327; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2329 = 14'h2b == field_data_lo_11 ? _field_data_T_47 : _GEN_2328; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2330 = 14'h2c == field_data_lo_11 ? _field_data_T_48 : _GEN_2329; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2331 = 14'h2d == field_data_lo_11 ? _field_data_T_49 : _GEN_2330; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2332 = 14'h2e == field_data_lo_11 ? _field_data_T_50 : _GEN_2331; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2333 = 14'h2f == field_data_lo_11 ? _field_data_T_51 : _GEN_2332; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2334 = 14'h30 == field_data_lo_11 ? _field_data_T_52 : _GEN_2333; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2335 = 14'h31 == field_data_lo_11 ? _field_data_T_53 : _GEN_2334; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2336 = 14'h32 == field_data_lo_11 ? _field_data_T_54 : _GEN_2335; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2337 = 14'h33 == field_data_lo_11 ? _field_data_T_55 : _GEN_2336; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2338 = 14'h34 == field_data_lo_11 ? _field_data_T_56 : _GEN_2337; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2339 = 14'h35 == field_data_lo_11 ? _field_data_T_57 : _GEN_2338; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2340 = 14'h36 == field_data_lo_11 ? _field_data_T_58 : _GEN_2339; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2341 = 14'h37 == field_data_lo_11 ? _field_data_T_59 : _GEN_2340; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2342 = 14'h38 == field_data_lo_11 ? _field_data_T_60 : _GEN_2341; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2343 = 14'h39 == field_data_lo_11 ? _field_data_T_61 : _GEN_2342; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2344 = 14'h3a == field_data_lo_11 ? _field_data_T_62 : _GEN_2343; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2345 = 14'h3b == field_data_lo_11 ? _field_data_T_63 : _GEN_2344; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2346 = 14'h3c == field_data_lo_11 ? _field_data_T_64 : _GEN_2345; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2347 = 14'h3d == field_data_lo_11 ? _field_data_T_65 : _GEN_2346; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2348 = 14'h3e == field_data_lo_11 ? _field_data_T_66 : _GEN_2347; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2349 = 14'h3f == field_data_lo_11 ? _field_data_T_67 : _GEN_2348; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2350 = 14'h40 == field_data_lo_11 ? _field_data_T_68 : _GEN_2349; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2351 = 14'h41 == field_data_lo_11 ? _field_data_T_69 : _GEN_2350; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2352 = 14'h42 == field_data_lo_11 ? _field_data_T_70 : _GEN_2351; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2353 = 14'h43 == field_data_lo_11 ? _field_data_T_71 : _GEN_2352; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2354 = 14'h44 == field_data_lo_11 ? _field_data_T_72 : _GEN_2353; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2355 = 14'h45 == field_data_lo_11 ? _field_data_T_73 : _GEN_2354; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2356 = 14'h46 == field_data_lo_11 ? _field_data_T_74 : _GEN_2355; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2357 = 14'h47 == field_data_lo_11 ? _field_data_T_75 : _GEN_2356; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2358 = 14'h48 == field_data_lo_11 ? _field_data_T_76 : _GEN_2357; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2359 = 14'h49 == field_data_lo_11 ? _field_data_T_77 : _GEN_2358; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2360 = 14'h4a == field_data_lo_11 ? _field_data_T_78 : _GEN_2359; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2361 = 14'h4b == field_data_lo_11 ? _field_data_T_79 : _GEN_2360; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2362 = 14'h4c == field_data_lo_11 ? _field_data_T_80 : _GEN_2361; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2363 = 14'h4d == field_data_lo_11 ? _field_data_T_81 : _GEN_2362; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2364 = 14'h4e == field_data_lo_11 ? _field_data_T_82 : _GEN_2363; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2365 = 14'h4f == field_data_lo_11 ? _field_data_T_83 : _GEN_2364; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_44 = vliw_44[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_12 = vliw_44[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_44 = field_data_lo_12[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_44 = field_data_lo_12[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_56 = {{1'd0}, args_offset_44}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_56 = _total_offset_T_56[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2369 = 3'h1 == total_offset_56 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2370 = 3'h2 == total_offset_56 ? args_2 : _GEN_2369; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2371 = 3'h3 == total_offset_56 ? args_3 : _GEN_2370; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2372 = 3'h4 == total_offset_56 ? args_4 : _GEN_2371; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2373 = 3'h5 == total_offset_56 ? args_5 : _GEN_2372; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2374 = 3'h6 == total_offset_56 ? args_6 : _GEN_2373; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2375 = total_offset_56 < 3'h7 ? _GEN_2374 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_44_1 = 3'h0 < args_length_44 ? _GEN_2375 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_57 = args_offset_44 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2378 = 3'h1 == total_offset_57 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2379 = 3'h2 == total_offset_57 ? args_2 : _GEN_2378; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2380 = 3'h3 == total_offset_57 ? args_3 : _GEN_2379; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2381 = 3'h4 == total_offset_57 ? args_4 : _GEN_2380; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2382 = 3'h5 == total_offset_57 ? args_5 : _GEN_2381; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2383 = 3'h6 == total_offset_57 ? args_6 : _GEN_2382; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2384 = total_offset_57 < 3'h7 ? _GEN_2383 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_44_0 = 3'h1 < args_length_44 ? _GEN_2384 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_656 = {field_bytes_44_0,field_bytes_44_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2386 = opcode_44 == 4'ha ? _field_data_T_656 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2387 = opcode_44 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1937 = opcode_44 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_12 = field_data_lo_12[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_659 = {field_data_hi_12,field_data_lo_12}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_89 = _T_1937 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2388 = opcode_44 == 4'h8 | opcode_44 == 4'hb ? _field_data_T_659 : _GEN_2386; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2389 = opcode_44 == 4'h8 | opcode_44 == 4'hb ? _field_tag_T_89 : _GEN_2387; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2390 = 14'h20 == field_data_lo_12 ? _field_data_T_36 : _GEN_2388; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2391 = 14'h21 == field_data_lo_12 ? _field_data_T_37 : _GEN_2390; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2392 = 14'h22 == field_data_lo_12 ? _field_data_T_38 : _GEN_2391; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2393 = 14'h23 == field_data_lo_12 ? _field_data_T_39 : _GEN_2392; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2394 = 14'h24 == field_data_lo_12 ? _field_data_T_40 : _GEN_2393; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2395 = 14'h25 == field_data_lo_12 ? _field_data_T_41 : _GEN_2394; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2396 = 14'h26 == field_data_lo_12 ? _field_data_T_42 : _GEN_2395; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2397 = 14'h27 == field_data_lo_12 ? _field_data_T_43 : _GEN_2396; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2398 = 14'h28 == field_data_lo_12 ? _field_data_T_44 : _GEN_2397; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2399 = 14'h29 == field_data_lo_12 ? _field_data_T_45 : _GEN_2398; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2400 = 14'h2a == field_data_lo_12 ? _field_data_T_46 : _GEN_2399; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2401 = 14'h2b == field_data_lo_12 ? _field_data_T_47 : _GEN_2400; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2402 = 14'h2c == field_data_lo_12 ? _field_data_T_48 : _GEN_2401; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2403 = 14'h2d == field_data_lo_12 ? _field_data_T_49 : _GEN_2402; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2404 = 14'h2e == field_data_lo_12 ? _field_data_T_50 : _GEN_2403; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2405 = 14'h2f == field_data_lo_12 ? _field_data_T_51 : _GEN_2404; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2406 = 14'h30 == field_data_lo_12 ? _field_data_T_52 : _GEN_2405; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2407 = 14'h31 == field_data_lo_12 ? _field_data_T_53 : _GEN_2406; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2408 = 14'h32 == field_data_lo_12 ? _field_data_T_54 : _GEN_2407; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2409 = 14'h33 == field_data_lo_12 ? _field_data_T_55 : _GEN_2408; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2410 = 14'h34 == field_data_lo_12 ? _field_data_T_56 : _GEN_2409; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2411 = 14'h35 == field_data_lo_12 ? _field_data_T_57 : _GEN_2410; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2412 = 14'h36 == field_data_lo_12 ? _field_data_T_58 : _GEN_2411; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2413 = 14'h37 == field_data_lo_12 ? _field_data_T_59 : _GEN_2412; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2414 = 14'h38 == field_data_lo_12 ? _field_data_T_60 : _GEN_2413; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2415 = 14'h39 == field_data_lo_12 ? _field_data_T_61 : _GEN_2414; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2416 = 14'h3a == field_data_lo_12 ? _field_data_T_62 : _GEN_2415; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2417 = 14'h3b == field_data_lo_12 ? _field_data_T_63 : _GEN_2416; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2418 = 14'h3c == field_data_lo_12 ? _field_data_T_64 : _GEN_2417; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2419 = 14'h3d == field_data_lo_12 ? _field_data_T_65 : _GEN_2418; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2420 = 14'h3e == field_data_lo_12 ? _field_data_T_66 : _GEN_2419; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2421 = 14'h3f == field_data_lo_12 ? _field_data_T_67 : _GEN_2420; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2422 = 14'h40 == field_data_lo_12 ? _field_data_T_68 : _GEN_2421; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2423 = 14'h41 == field_data_lo_12 ? _field_data_T_69 : _GEN_2422; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2424 = 14'h42 == field_data_lo_12 ? _field_data_T_70 : _GEN_2423; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2425 = 14'h43 == field_data_lo_12 ? _field_data_T_71 : _GEN_2424; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2426 = 14'h44 == field_data_lo_12 ? _field_data_T_72 : _GEN_2425; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2427 = 14'h45 == field_data_lo_12 ? _field_data_T_73 : _GEN_2426; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2428 = 14'h46 == field_data_lo_12 ? _field_data_T_74 : _GEN_2427; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2429 = 14'h47 == field_data_lo_12 ? _field_data_T_75 : _GEN_2428; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2430 = 14'h48 == field_data_lo_12 ? _field_data_T_76 : _GEN_2429; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2431 = 14'h49 == field_data_lo_12 ? _field_data_T_77 : _GEN_2430; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2432 = 14'h4a == field_data_lo_12 ? _field_data_T_78 : _GEN_2431; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2433 = 14'h4b == field_data_lo_12 ? _field_data_T_79 : _GEN_2432; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2434 = 14'h4c == field_data_lo_12 ? _field_data_T_80 : _GEN_2433; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2435 = 14'h4d == field_data_lo_12 ? _field_data_T_81 : _GEN_2434; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2436 = 14'h4e == field_data_lo_12 ? _field_data_T_82 : _GEN_2435; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2437 = 14'h4f == field_data_lo_12 ? _field_data_T_83 : _GEN_2436; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_45 = vliw_45[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_13 = vliw_45[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_45 = field_data_lo_13[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_45 = field_data_lo_13[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_58 = {{1'd0}, args_offset_45}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_58 = _total_offset_T_58[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2441 = 3'h1 == total_offset_58 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2442 = 3'h2 == total_offset_58 ? args_2 : _GEN_2441; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2443 = 3'h3 == total_offset_58 ? args_3 : _GEN_2442; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2444 = 3'h4 == total_offset_58 ? args_4 : _GEN_2443; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2445 = 3'h5 == total_offset_58 ? args_5 : _GEN_2444; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2446 = 3'h6 == total_offset_58 ? args_6 : _GEN_2445; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2447 = total_offset_58 < 3'h7 ? _GEN_2446 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_45_1 = 3'h0 < args_length_45 ? _GEN_2447 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_59 = args_offset_45 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2450 = 3'h1 == total_offset_59 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2451 = 3'h2 == total_offset_59 ? args_2 : _GEN_2450; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2452 = 3'h3 == total_offset_59 ? args_3 : _GEN_2451; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2453 = 3'h4 == total_offset_59 ? args_4 : _GEN_2452; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2454 = 3'h5 == total_offset_59 ? args_5 : _GEN_2453; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2455 = 3'h6 == total_offset_59 ? args_6 : _GEN_2454; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2456 = total_offset_59 < 3'h7 ? _GEN_2455 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_45_0 = 3'h1 < args_length_45 ? _GEN_2456 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_708 = {field_bytes_45_0,field_bytes_45_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2458 = opcode_45 == 4'ha ? _field_data_T_708 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2459 = opcode_45 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1994 = opcode_45 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_13 = field_data_lo_13[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_711 = {field_data_hi_13,field_data_lo_13}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_91 = _T_1994 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2460 = opcode_45 == 4'h8 | opcode_45 == 4'hb ? _field_data_T_711 : _GEN_2458; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2461 = opcode_45 == 4'h8 | opcode_45 == 4'hb ? _field_tag_T_91 : _GEN_2459; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2462 = 14'h20 == field_data_lo_13 ? _field_data_T_36 : _GEN_2460; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2463 = 14'h21 == field_data_lo_13 ? _field_data_T_37 : _GEN_2462; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2464 = 14'h22 == field_data_lo_13 ? _field_data_T_38 : _GEN_2463; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2465 = 14'h23 == field_data_lo_13 ? _field_data_T_39 : _GEN_2464; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2466 = 14'h24 == field_data_lo_13 ? _field_data_T_40 : _GEN_2465; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2467 = 14'h25 == field_data_lo_13 ? _field_data_T_41 : _GEN_2466; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2468 = 14'h26 == field_data_lo_13 ? _field_data_T_42 : _GEN_2467; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2469 = 14'h27 == field_data_lo_13 ? _field_data_T_43 : _GEN_2468; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2470 = 14'h28 == field_data_lo_13 ? _field_data_T_44 : _GEN_2469; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2471 = 14'h29 == field_data_lo_13 ? _field_data_T_45 : _GEN_2470; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2472 = 14'h2a == field_data_lo_13 ? _field_data_T_46 : _GEN_2471; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2473 = 14'h2b == field_data_lo_13 ? _field_data_T_47 : _GEN_2472; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2474 = 14'h2c == field_data_lo_13 ? _field_data_T_48 : _GEN_2473; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2475 = 14'h2d == field_data_lo_13 ? _field_data_T_49 : _GEN_2474; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2476 = 14'h2e == field_data_lo_13 ? _field_data_T_50 : _GEN_2475; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2477 = 14'h2f == field_data_lo_13 ? _field_data_T_51 : _GEN_2476; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2478 = 14'h30 == field_data_lo_13 ? _field_data_T_52 : _GEN_2477; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2479 = 14'h31 == field_data_lo_13 ? _field_data_T_53 : _GEN_2478; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2480 = 14'h32 == field_data_lo_13 ? _field_data_T_54 : _GEN_2479; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2481 = 14'h33 == field_data_lo_13 ? _field_data_T_55 : _GEN_2480; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2482 = 14'h34 == field_data_lo_13 ? _field_data_T_56 : _GEN_2481; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2483 = 14'h35 == field_data_lo_13 ? _field_data_T_57 : _GEN_2482; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2484 = 14'h36 == field_data_lo_13 ? _field_data_T_58 : _GEN_2483; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2485 = 14'h37 == field_data_lo_13 ? _field_data_T_59 : _GEN_2484; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2486 = 14'h38 == field_data_lo_13 ? _field_data_T_60 : _GEN_2485; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2487 = 14'h39 == field_data_lo_13 ? _field_data_T_61 : _GEN_2486; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2488 = 14'h3a == field_data_lo_13 ? _field_data_T_62 : _GEN_2487; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2489 = 14'h3b == field_data_lo_13 ? _field_data_T_63 : _GEN_2488; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2490 = 14'h3c == field_data_lo_13 ? _field_data_T_64 : _GEN_2489; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2491 = 14'h3d == field_data_lo_13 ? _field_data_T_65 : _GEN_2490; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2492 = 14'h3e == field_data_lo_13 ? _field_data_T_66 : _GEN_2491; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2493 = 14'h3f == field_data_lo_13 ? _field_data_T_67 : _GEN_2492; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2494 = 14'h40 == field_data_lo_13 ? _field_data_T_68 : _GEN_2493; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2495 = 14'h41 == field_data_lo_13 ? _field_data_T_69 : _GEN_2494; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2496 = 14'h42 == field_data_lo_13 ? _field_data_T_70 : _GEN_2495; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2497 = 14'h43 == field_data_lo_13 ? _field_data_T_71 : _GEN_2496; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2498 = 14'h44 == field_data_lo_13 ? _field_data_T_72 : _GEN_2497; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2499 = 14'h45 == field_data_lo_13 ? _field_data_T_73 : _GEN_2498; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2500 = 14'h46 == field_data_lo_13 ? _field_data_T_74 : _GEN_2499; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2501 = 14'h47 == field_data_lo_13 ? _field_data_T_75 : _GEN_2500; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2502 = 14'h48 == field_data_lo_13 ? _field_data_T_76 : _GEN_2501; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2503 = 14'h49 == field_data_lo_13 ? _field_data_T_77 : _GEN_2502; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2504 = 14'h4a == field_data_lo_13 ? _field_data_T_78 : _GEN_2503; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2505 = 14'h4b == field_data_lo_13 ? _field_data_T_79 : _GEN_2504; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2506 = 14'h4c == field_data_lo_13 ? _field_data_T_80 : _GEN_2505; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2507 = 14'h4d == field_data_lo_13 ? _field_data_T_81 : _GEN_2506; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2508 = 14'h4e == field_data_lo_13 ? _field_data_T_82 : _GEN_2507; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2509 = 14'h4f == field_data_lo_13 ? _field_data_T_83 : _GEN_2508; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_46 = vliw_46[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_14 = vliw_46[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_46 = field_data_lo_14[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_46 = field_data_lo_14[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_60 = {{1'd0}, args_offset_46}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_60 = _total_offset_T_60[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2513 = 3'h1 == total_offset_60 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2514 = 3'h2 == total_offset_60 ? args_2 : _GEN_2513; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2515 = 3'h3 == total_offset_60 ? args_3 : _GEN_2514; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2516 = 3'h4 == total_offset_60 ? args_4 : _GEN_2515; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2517 = 3'h5 == total_offset_60 ? args_5 : _GEN_2516; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2518 = 3'h6 == total_offset_60 ? args_6 : _GEN_2517; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2519 = total_offset_60 < 3'h7 ? _GEN_2518 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_46_1 = 3'h0 < args_length_46 ? _GEN_2519 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_61 = args_offset_46 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2522 = 3'h1 == total_offset_61 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2523 = 3'h2 == total_offset_61 ? args_2 : _GEN_2522; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2524 = 3'h3 == total_offset_61 ? args_3 : _GEN_2523; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2525 = 3'h4 == total_offset_61 ? args_4 : _GEN_2524; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2526 = 3'h5 == total_offset_61 ? args_5 : _GEN_2525; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2527 = 3'h6 == total_offset_61 ? args_6 : _GEN_2526; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2528 = total_offset_61 < 3'h7 ? _GEN_2527 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_46_0 = 3'h1 < args_length_46 ? _GEN_2528 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_760 = {field_bytes_46_0,field_bytes_46_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2530 = opcode_46 == 4'ha ? _field_data_T_760 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2531 = opcode_46 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2051 = opcode_46 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_14 = field_data_lo_14[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_763 = {field_data_hi_14,field_data_lo_14}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_93 = _T_2051 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2532 = opcode_46 == 4'h8 | opcode_46 == 4'hb ? _field_data_T_763 : _GEN_2530; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2533 = opcode_46 == 4'h8 | opcode_46 == 4'hb ? _field_tag_T_93 : _GEN_2531; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2534 = 14'h20 == field_data_lo_14 ? _field_data_T_36 : _GEN_2532; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2535 = 14'h21 == field_data_lo_14 ? _field_data_T_37 : _GEN_2534; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2536 = 14'h22 == field_data_lo_14 ? _field_data_T_38 : _GEN_2535; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2537 = 14'h23 == field_data_lo_14 ? _field_data_T_39 : _GEN_2536; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2538 = 14'h24 == field_data_lo_14 ? _field_data_T_40 : _GEN_2537; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2539 = 14'h25 == field_data_lo_14 ? _field_data_T_41 : _GEN_2538; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2540 = 14'h26 == field_data_lo_14 ? _field_data_T_42 : _GEN_2539; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2541 = 14'h27 == field_data_lo_14 ? _field_data_T_43 : _GEN_2540; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2542 = 14'h28 == field_data_lo_14 ? _field_data_T_44 : _GEN_2541; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2543 = 14'h29 == field_data_lo_14 ? _field_data_T_45 : _GEN_2542; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2544 = 14'h2a == field_data_lo_14 ? _field_data_T_46 : _GEN_2543; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2545 = 14'h2b == field_data_lo_14 ? _field_data_T_47 : _GEN_2544; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2546 = 14'h2c == field_data_lo_14 ? _field_data_T_48 : _GEN_2545; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2547 = 14'h2d == field_data_lo_14 ? _field_data_T_49 : _GEN_2546; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2548 = 14'h2e == field_data_lo_14 ? _field_data_T_50 : _GEN_2547; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2549 = 14'h2f == field_data_lo_14 ? _field_data_T_51 : _GEN_2548; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2550 = 14'h30 == field_data_lo_14 ? _field_data_T_52 : _GEN_2549; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2551 = 14'h31 == field_data_lo_14 ? _field_data_T_53 : _GEN_2550; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2552 = 14'h32 == field_data_lo_14 ? _field_data_T_54 : _GEN_2551; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2553 = 14'h33 == field_data_lo_14 ? _field_data_T_55 : _GEN_2552; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2554 = 14'h34 == field_data_lo_14 ? _field_data_T_56 : _GEN_2553; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2555 = 14'h35 == field_data_lo_14 ? _field_data_T_57 : _GEN_2554; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2556 = 14'h36 == field_data_lo_14 ? _field_data_T_58 : _GEN_2555; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2557 = 14'h37 == field_data_lo_14 ? _field_data_T_59 : _GEN_2556; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2558 = 14'h38 == field_data_lo_14 ? _field_data_T_60 : _GEN_2557; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2559 = 14'h39 == field_data_lo_14 ? _field_data_T_61 : _GEN_2558; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2560 = 14'h3a == field_data_lo_14 ? _field_data_T_62 : _GEN_2559; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2561 = 14'h3b == field_data_lo_14 ? _field_data_T_63 : _GEN_2560; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2562 = 14'h3c == field_data_lo_14 ? _field_data_T_64 : _GEN_2561; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2563 = 14'h3d == field_data_lo_14 ? _field_data_T_65 : _GEN_2562; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2564 = 14'h3e == field_data_lo_14 ? _field_data_T_66 : _GEN_2563; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2565 = 14'h3f == field_data_lo_14 ? _field_data_T_67 : _GEN_2564; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2566 = 14'h40 == field_data_lo_14 ? _field_data_T_68 : _GEN_2565; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2567 = 14'h41 == field_data_lo_14 ? _field_data_T_69 : _GEN_2566; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2568 = 14'h42 == field_data_lo_14 ? _field_data_T_70 : _GEN_2567; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2569 = 14'h43 == field_data_lo_14 ? _field_data_T_71 : _GEN_2568; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2570 = 14'h44 == field_data_lo_14 ? _field_data_T_72 : _GEN_2569; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2571 = 14'h45 == field_data_lo_14 ? _field_data_T_73 : _GEN_2570; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2572 = 14'h46 == field_data_lo_14 ? _field_data_T_74 : _GEN_2571; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2573 = 14'h47 == field_data_lo_14 ? _field_data_T_75 : _GEN_2572; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2574 = 14'h48 == field_data_lo_14 ? _field_data_T_76 : _GEN_2573; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2575 = 14'h49 == field_data_lo_14 ? _field_data_T_77 : _GEN_2574; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2576 = 14'h4a == field_data_lo_14 ? _field_data_T_78 : _GEN_2575; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2577 = 14'h4b == field_data_lo_14 ? _field_data_T_79 : _GEN_2576; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2578 = 14'h4c == field_data_lo_14 ? _field_data_T_80 : _GEN_2577; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2579 = 14'h4d == field_data_lo_14 ? _field_data_T_81 : _GEN_2578; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2580 = 14'h4e == field_data_lo_14 ? _field_data_T_82 : _GEN_2579; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2581 = 14'h4f == field_data_lo_14 ? _field_data_T_83 : _GEN_2580; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_47 = vliw_47[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_15 = vliw_47[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_47 = field_data_lo_15[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_47 = field_data_lo_15[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_62 = {{1'd0}, args_offset_47}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_62 = _total_offset_T_62[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2585 = 3'h1 == total_offset_62 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2586 = 3'h2 == total_offset_62 ? args_2 : _GEN_2585; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2587 = 3'h3 == total_offset_62 ? args_3 : _GEN_2586; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2588 = 3'h4 == total_offset_62 ? args_4 : _GEN_2587; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2589 = 3'h5 == total_offset_62 ? args_5 : _GEN_2588; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2590 = 3'h6 == total_offset_62 ? args_6 : _GEN_2589; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2591 = total_offset_62 < 3'h7 ? _GEN_2590 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_47_1 = 3'h0 < args_length_47 ? _GEN_2591 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_63 = args_offset_47 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2594 = 3'h1 == total_offset_63 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2595 = 3'h2 == total_offset_63 ? args_2 : _GEN_2594; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2596 = 3'h3 == total_offset_63 ? args_3 : _GEN_2595; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2597 = 3'h4 == total_offset_63 ? args_4 : _GEN_2596; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2598 = 3'h5 == total_offset_63 ? args_5 : _GEN_2597; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2599 = 3'h6 == total_offset_63 ? args_6 : _GEN_2598; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2600 = total_offset_63 < 3'h7 ? _GEN_2599 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_47_0 = 3'h1 < args_length_47 ? _GEN_2600 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_812 = {field_bytes_47_0,field_bytes_47_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2602 = opcode_47 == 4'ha ? _field_data_T_812 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2603 = opcode_47 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2108 = opcode_47 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_15 = field_data_lo_15[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_815 = {field_data_hi_15,field_data_lo_15}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_95 = _T_2108 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2604 = opcode_47 == 4'h8 | opcode_47 == 4'hb ? _field_data_T_815 : _GEN_2602; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2605 = opcode_47 == 4'h8 | opcode_47 == 4'hb ? _field_tag_T_95 : _GEN_2603; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2606 = 14'h20 == field_data_lo_15 ? _field_data_T_36 : _GEN_2604; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2607 = 14'h21 == field_data_lo_15 ? _field_data_T_37 : _GEN_2606; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2608 = 14'h22 == field_data_lo_15 ? _field_data_T_38 : _GEN_2607; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2609 = 14'h23 == field_data_lo_15 ? _field_data_T_39 : _GEN_2608; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2610 = 14'h24 == field_data_lo_15 ? _field_data_T_40 : _GEN_2609; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2611 = 14'h25 == field_data_lo_15 ? _field_data_T_41 : _GEN_2610; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2612 = 14'h26 == field_data_lo_15 ? _field_data_T_42 : _GEN_2611; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2613 = 14'h27 == field_data_lo_15 ? _field_data_T_43 : _GEN_2612; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2614 = 14'h28 == field_data_lo_15 ? _field_data_T_44 : _GEN_2613; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2615 = 14'h29 == field_data_lo_15 ? _field_data_T_45 : _GEN_2614; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2616 = 14'h2a == field_data_lo_15 ? _field_data_T_46 : _GEN_2615; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2617 = 14'h2b == field_data_lo_15 ? _field_data_T_47 : _GEN_2616; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2618 = 14'h2c == field_data_lo_15 ? _field_data_T_48 : _GEN_2617; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2619 = 14'h2d == field_data_lo_15 ? _field_data_T_49 : _GEN_2618; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2620 = 14'h2e == field_data_lo_15 ? _field_data_T_50 : _GEN_2619; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2621 = 14'h2f == field_data_lo_15 ? _field_data_T_51 : _GEN_2620; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2622 = 14'h30 == field_data_lo_15 ? _field_data_T_52 : _GEN_2621; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2623 = 14'h31 == field_data_lo_15 ? _field_data_T_53 : _GEN_2622; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2624 = 14'h32 == field_data_lo_15 ? _field_data_T_54 : _GEN_2623; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2625 = 14'h33 == field_data_lo_15 ? _field_data_T_55 : _GEN_2624; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2626 = 14'h34 == field_data_lo_15 ? _field_data_T_56 : _GEN_2625; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2627 = 14'h35 == field_data_lo_15 ? _field_data_T_57 : _GEN_2626; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2628 = 14'h36 == field_data_lo_15 ? _field_data_T_58 : _GEN_2627; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2629 = 14'h37 == field_data_lo_15 ? _field_data_T_59 : _GEN_2628; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2630 = 14'h38 == field_data_lo_15 ? _field_data_T_60 : _GEN_2629; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2631 = 14'h39 == field_data_lo_15 ? _field_data_T_61 : _GEN_2630; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2632 = 14'h3a == field_data_lo_15 ? _field_data_T_62 : _GEN_2631; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2633 = 14'h3b == field_data_lo_15 ? _field_data_T_63 : _GEN_2632; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2634 = 14'h3c == field_data_lo_15 ? _field_data_T_64 : _GEN_2633; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2635 = 14'h3d == field_data_lo_15 ? _field_data_T_65 : _GEN_2634; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2636 = 14'h3e == field_data_lo_15 ? _field_data_T_66 : _GEN_2635; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2637 = 14'h3f == field_data_lo_15 ? _field_data_T_67 : _GEN_2636; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2638 = 14'h40 == field_data_lo_15 ? _field_data_T_68 : _GEN_2637; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2639 = 14'h41 == field_data_lo_15 ? _field_data_T_69 : _GEN_2638; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2640 = 14'h42 == field_data_lo_15 ? _field_data_T_70 : _GEN_2639; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2641 = 14'h43 == field_data_lo_15 ? _field_data_T_71 : _GEN_2640; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2642 = 14'h44 == field_data_lo_15 ? _field_data_T_72 : _GEN_2641; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2643 = 14'h45 == field_data_lo_15 ? _field_data_T_73 : _GEN_2642; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2644 = 14'h46 == field_data_lo_15 ? _field_data_T_74 : _GEN_2643; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2645 = 14'h47 == field_data_lo_15 ? _field_data_T_75 : _GEN_2644; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2646 = 14'h48 == field_data_lo_15 ? _field_data_T_76 : _GEN_2645; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2647 = 14'h49 == field_data_lo_15 ? _field_data_T_77 : _GEN_2646; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2648 = 14'h4a == field_data_lo_15 ? _field_data_T_78 : _GEN_2647; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2649 = 14'h4b == field_data_lo_15 ? _field_data_T_79 : _GEN_2648; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2650 = 14'h4c == field_data_lo_15 ? _field_data_T_80 : _GEN_2649; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2651 = 14'h4d == field_data_lo_15 ? _field_data_T_81 : _GEN_2650; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2652 = 14'h4e == field_data_lo_15 ? _field_data_T_82 : _GEN_2651; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2653 = 14'h4f == field_data_lo_15 ? _field_data_T_83 : _GEN_2652; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_48 = vliw_48[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_16 = vliw_48[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_48 = field_data_lo_16[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_48 = field_data_lo_16[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_64 = {{1'd0}, args_offset_48}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_64 = _total_offset_T_64[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2657 = 3'h1 == total_offset_64 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2658 = 3'h2 == total_offset_64 ? args_2 : _GEN_2657; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2659 = 3'h3 == total_offset_64 ? args_3 : _GEN_2658; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2660 = 3'h4 == total_offset_64 ? args_4 : _GEN_2659; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2661 = 3'h5 == total_offset_64 ? args_5 : _GEN_2660; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2662 = 3'h6 == total_offset_64 ? args_6 : _GEN_2661; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2663 = total_offset_64 < 3'h7 ? _GEN_2662 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_48_1 = 3'h0 < args_length_48 ? _GEN_2663 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_65 = args_offset_48 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2666 = 3'h1 == total_offset_65 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2667 = 3'h2 == total_offset_65 ? args_2 : _GEN_2666; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2668 = 3'h3 == total_offset_65 ? args_3 : _GEN_2667; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2669 = 3'h4 == total_offset_65 ? args_4 : _GEN_2668; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2670 = 3'h5 == total_offset_65 ? args_5 : _GEN_2669; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2671 = 3'h6 == total_offset_65 ? args_6 : _GEN_2670; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2672 = total_offset_65 < 3'h7 ? _GEN_2671 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_48_0 = 3'h1 < args_length_48 ? _GEN_2672 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_864 = {field_bytes_48_0,field_bytes_48_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2674 = opcode_48 == 4'ha ? _field_data_T_864 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2675 = opcode_48 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2165 = opcode_48 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_16 = field_data_lo_16[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_867 = {field_data_hi_16,field_data_lo_16}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_97 = _T_2165 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2676 = opcode_48 == 4'h8 | opcode_48 == 4'hb ? _field_data_T_867 : _GEN_2674; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2677 = opcode_48 == 4'h8 | opcode_48 == 4'hb ? _field_tag_T_97 : _GEN_2675; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2678 = 14'h20 == field_data_lo_16 ? _field_data_T_36 : _GEN_2676; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2679 = 14'h21 == field_data_lo_16 ? _field_data_T_37 : _GEN_2678; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2680 = 14'h22 == field_data_lo_16 ? _field_data_T_38 : _GEN_2679; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2681 = 14'h23 == field_data_lo_16 ? _field_data_T_39 : _GEN_2680; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2682 = 14'h24 == field_data_lo_16 ? _field_data_T_40 : _GEN_2681; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2683 = 14'h25 == field_data_lo_16 ? _field_data_T_41 : _GEN_2682; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2684 = 14'h26 == field_data_lo_16 ? _field_data_T_42 : _GEN_2683; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2685 = 14'h27 == field_data_lo_16 ? _field_data_T_43 : _GEN_2684; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2686 = 14'h28 == field_data_lo_16 ? _field_data_T_44 : _GEN_2685; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2687 = 14'h29 == field_data_lo_16 ? _field_data_T_45 : _GEN_2686; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2688 = 14'h2a == field_data_lo_16 ? _field_data_T_46 : _GEN_2687; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2689 = 14'h2b == field_data_lo_16 ? _field_data_T_47 : _GEN_2688; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2690 = 14'h2c == field_data_lo_16 ? _field_data_T_48 : _GEN_2689; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2691 = 14'h2d == field_data_lo_16 ? _field_data_T_49 : _GEN_2690; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2692 = 14'h2e == field_data_lo_16 ? _field_data_T_50 : _GEN_2691; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2693 = 14'h2f == field_data_lo_16 ? _field_data_T_51 : _GEN_2692; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2694 = 14'h30 == field_data_lo_16 ? _field_data_T_52 : _GEN_2693; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2695 = 14'h31 == field_data_lo_16 ? _field_data_T_53 : _GEN_2694; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2696 = 14'h32 == field_data_lo_16 ? _field_data_T_54 : _GEN_2695; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2697 = 14'h33 == field_data_lo_16 ? _field_data_T_55 : _GEN_2696; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2698 = 14'h34 == field_data_lo_16 ? _field_data_T_56 : _GEN_2697; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2699 = 14'h35 == field_data_lo_16 ? _field_data_T_57 : _GEN_2698; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2700 = 14'h36 == field_data_lo_16 ? _field_data_T_58 : _GEN_2699; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2701 = 14'h37 == field_data_lo_16 ? _field_data_T_59 : _GEN_2700; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2702 = 14'h38 == field_data_lo_16 ? _field_data_T_60 : _GEN_2701; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2703 = 14'h39 == field_data_lo_16 ? _field_data_T_61 : _GEN_2702; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2704 = 14'h3a == field_data_lo_16 ? _field_data_T_62 : _GEN_2703; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2705 = 14'h3b == field_data_lo_16 ? _field_data_T_63 : _GEN_2704; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2706 = 14'h3c == field_data_lo_16 ? _field_data_T_64 : _GEN_2705; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2707 = 14'h3d == field_data_lo_16 ? _field_data_T_65 : _GEN_2706; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2708 = 14'h3e == field_data_lo_16 ? _field_data_T_66 : _GEN_2707; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2709 = 14'h3f == field_data_lo_16 ? _field_data_T_67 : _GEN_2708; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2710 = 14'h40 == field_data_lo_16 ? _field_data_T_68 : _GEN_2709; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2711 = 14'h41 == field_data_lo_16 ? _field_data_T_69 : _GEN_2710; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2712 = 14'h42 == field_data_lo_16 ? _field_data_T_70 : _GEN_2711; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2713 = 14'h43 == field_data_lo_16 ? _field_data_T_71 : _GEN_2712; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2714 = 14'h44 == field_data_lo_16 ? _field_data_T_72 : _GEN_2713; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2715 = 14'h45 == field_data_lo_16 ? _field_data_T_73 : _GEN_2714; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2716 = 14'h46 == field_data_lo_16 ? _field_data_T_74 : _GEN_2715; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2717 = 14'h47 == field_data_lo_16 ? _field_data_T_75 : _GEN_2716; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2718 = 14'h48 == field_data_lo_16 ? _field_data_T_76 : _GEN_2717; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2719 = 14'h49 == field_data_lo_16 ? _field_data_T_77 : _GEN_2718; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2720 = 14'h4a == field_data_lo_16 ? _field_data_T_78 : _GEN_2719; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2721 = 14'h4b == field_data_lo_16 ? _field_data_T_79 : _GEN_2720; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2722 = 14'h4c == field_data_lo_16 ? _field_data_T_80 : _GEN_2721; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2723 = 14'h4d == field_data_lo_16 ? _field_data_T_81 : _GEN_2722; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2724 = 14'h4e == field_data_lo_16 ? _field_data_T_82 : _GEN_2723; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2725 = 14'h4f == field_data_lo_16 ? _field_data_T_83 : _GEN_2724; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_49 = vliw_49[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_17 = vliw_49[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_49 = field_data_lo_17[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_49 = field_data_lo_17[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_66 = {{1'd0}, args_offset_49}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_66 = _total_offset_T_66[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2729 = 3'h1 == total_offset_66 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2730 = 3'h2 == total_offset_66 ? args_2 : _GEN_2729; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2731 = 3'h3 == total_offset_66 ? args_3 : _GEN_2730; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2732 = 3'h4 == total_offset_66 ? args_4 : _GEN_2731; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2733 = 3'h5 == total_offset_66 ? args_5 : _GEN_2732; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2734 = 3'h6 == total_offset_66 ? args_6 : _GEN_2733; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2735 = total_offset_66 < 3'h7 ? _GEN_2734 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_49_1 = 3'h0 < args_length_49 ? _GEN_2735 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_67 = args_offset_49 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2738 = 3'h1 == total_offset_67 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2739 = 3'h2 == total_offset_67 ? args_2 : _GEN_2738; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2740 = 3'h3 == total_offset_67 ? args_3 : _GEN_2739; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2741 = 3'h4 == total_offset_67 ? args_4 : _GEN_2740; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2742 = 3'h5 == total_offset_67 ? args_5 : _GEN_2741; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2743 = 3'h6 == total_offset_67 ? args_6 : _GEN_2742; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2744 = total_offset_67 < 3'h7 ? _GEN_2743 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_49_0 = 3'h1 < args_length_49 ? _GEN_2744 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_916 = {field_bytes_49_0,field_bytes_49_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2746 = opcode_49 == 4'ha ? _field_data_T_916 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2747 = opcode_49 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2222 = opcode_49 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_17 = field_data_lo_17[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_919 = {field_data_hi_17,field_data_lo_17}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_99 = _T_2222 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2748 = opcode_49 == 4'h8 | opcode_49 == 4'hb ? _field_data_T_919 : _GEN_2746; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2749 = opcode_49 == 4'h8 | opcode_49 == 4'hb ? _field_tag_T_99 : _GEN_2747; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2750 = 14'h20 == field_data_lo_17 ? _field_data_T_36 : _GEN_2748; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2751 = 14'h21 == field_data_lo_17 ? _field_data_T_37 : _GEN_2750; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2752 = 14'h22 == field_data_lo_17 ? _field_data_T_38 : _GEN_2751; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2753 = 14'h23 == field_data_lo_17 ? _field_data_T_39 : _GEN_2752; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2754 = 14'h24 == field_data_lo_17 ? _field_data_T_40 : _GEN_2753; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2755 = 14'h25 == field_data_lo_17 ? _field_data_T_41 : _GEN_2754; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2756 = 14'h26 == field_data_lo_17 ? _field_data_T_42 : _GEN_2755; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2757 = 14'h27 == field_data_lo_17 ? _field_data_T_43 : _GEN_2756; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2758 = 14'h28 == field_data_lo_17 ? _field_data_T_44 : _GEN_2757; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2759 = 14'h29 == field_data_lo_17 ? _field_data_T_45 : _GEN_2758; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2760 = 14'h2a == field_data_lo_17 ? _field_data_T_46 : _GEN_2759; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2761 = 14'h2b == field_data_lo_17 ? _field_data_T_47 : _GEN_2760; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2762 = 14'h2c == field_data_lo_17 ? _field_data_T_48 : _GEN_2761; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2763 = 14'h2d == field_data_lo_17 ? _field_data_T_49 : _GEN_2762; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2764 = 14'h2e == field_data_lo_17 ? _field_data_T_50 : _GEN_2763; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2765 = 14'h2f == field_data_lo_17 ? _field_data_T_51 : _GEN_2764; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2766 = 14'h30 == field_data_lo_17 ? _field_data_T_52 : _GEN_2765; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2767 = 14'h31 == field_data_lo_17 ? _field_data_T_53 : _GEN_2766; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2768 = 14'h32 == field_data_lo_17 ? _field_data_T_54 : _GEN_2767; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2769 = 14'h33 == field_data_lo_17 ? _field_data_T_55 : _GEN_2768; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2770 = 14'h34 == field_data_lo_17 ? _field_data_T_56 : _GEN_2769; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2771 = 14'h35 == field_data_lo_17 ? _field_data_T_57 : _GEN_2770; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2772 = 14'h36 == field_data_lo_17 ? _field_data_T_58 : _GEN_2771; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2773 = 14'h37 == field_data_lo_17 ? _field_data_T_59 : _GEN_2772; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2774 = 14'h38 == field_data_lo_17 ? _field_data_T_60 : _GEN_2773; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2775 = 14'h39 == field_data_lo_17 ? _field_data_T_61 : _GEN_2774; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2776 = 14'h3a == field_data_lo_17 ? _field_data_T_62 : _GEN_2775; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2777 = 14'h3b == field_data_lo_17 ? _field_data_T_63 : _GEN_2776; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2778 = 14'h3c == field_data_lo_17 ? _field_data_T_64 : _GEN_2777; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2779 = 14'h3d == field_data_lo_17 ? _field_data_T_65 : _GEN_2778; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2780 = 14'h3e == field_data_lo_17 ? _field_data_T_66 : _GEN_2779; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2781 = 14'h3f == field_data_lo_17 ? _field_data_T_67 : _GEN_2780; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2782 = 14'h40 == field_data_lo_17 ? _field_data_T_68 : _GEN_2781; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2783 = 14'h41 == field_data_lo_17 ? _field_data_T_69 : _GEN_2782; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2784 = 14'h42 == field_data_lo_17 ? _field_data_T_70 : _GEN_2783; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2785 = 14'h43 == field_data_lo_17 ? _field_data_T_71 : _GEN_2784; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2786 = 14'h44 == field_data_lo_17 ? _field_data_T_72 : _GEN_2785; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2787 = 14'h45 == field_data_lo_17 ? _field_data_T_73 : _GEN_2786; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2788 = 14'h46 == field_data_lo_17 ? _field_data_T_74 : _GEN_2787; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2789 = 14'h47 == field_data_lo_17 ? _field_data_T_75 : _GEN_2788; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2790 = 14'h48 == field_data_lo_17 ? _field_data_T_76 : _GEN_2789; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2791 = 14'h49 == field_data_lo_17 ? _field_data_T_77 : _GEN_2790; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2792 = 14'h4a == field_data_lo_17 ? _field_data_T_78 : _GEN_2791; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2793 = 14'h4b == field_data_lo_17 ? _field_data_T_79 : _GEN_2792; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2794 = 14'h4c == field_data_lo_17 ? _field_data_T_80 : _GEN_2793; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2795 = 14'h4d == field_data_lo_17 ? _field_data_T_81 : _GEN_2794; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2796 = 14'h4e == field_data_lo_17 ? _field_data_T_82 : _GEN_2795; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2797 = 14'h4f == field_data_lo_17 ? _field_data_T_83 : _GEN_2796; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_50 = vliw_50[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_18 = vliw_50[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_50 = field_data_lo_18[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_50 = field_data_lo_18[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_68 = {{1'd0}, args_offset_50}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_68 = _total_offset_T_68[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2801 = 3'h1 == total_offset_68 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2802 = 3'h2 == total_offset_68 ? args_2 : _GEN_2801; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2803 = 3'h3 == total_offset_68 ? args_3 : _GEN_2802; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2804 = 3'h4 == total_offset_68 ? args_4 : _GEN_2803; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2805 = 3'h5 == total_offset_68 ? args_5 : _GEN_2804; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2806 = 3'h6 == total_offset_68 ? args_6 : _GEN_2805; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2807 = total_offset_68 < 3'h7 ? _GEN_2806 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_50_1 = 3'h0 < args_length_50 ? _GEN_2807 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_69 = args_offset_50 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2810 = 3'h1 == total_offset_69 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2811 = 3'h2 == total_offset_69 ? args_2 : _GEN_2810; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2812 = 3'h3 == total_offset_69 ? args_3 : _GEN_2811; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2813 = 3'h4 == total_offset_69 ? args_4 : _GEN_2812; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2814 = 3'h5 == total_offset_69 ? args_5 : _GEN_2813; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2815 = 3'h6 == total_offset_69 ? args_6 : _GEN_2814; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2816 = total_offset_69 < 3'h7 ? _GEN_2815 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_50_0 = 3'h1 < args_length_50 ? _GEN_2816 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_968 = {field_bytes_50_0,field_bytes_50_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2818 = opcode_50 == 4'ha ? _field_data_T_968 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2819 = opcode_50 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2279 = opcode_50 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_18 = field_data_lo_18[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_971 = {field_data_hi_18,field_data_lo_18}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_101 = _T_2279 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2820 = opcode_50 == 4'h8 | opcode_50 == 4'hb ? _field_data_T_971 : _GEN_2818; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2821 = opcode_50 == 4'h8 | opcode_50 == 4'hb ? _field_tag_T_101 : _GEN_2819; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2822 = 14'h20 == field_data_lo_18 ? _field_data_T_36 : _GEN_2820; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2823 = 14'h21 == field_data_lo_18 ? _field_data_T_37 : _GEN_2822; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2824 = 14'h22 == field_data_lo_18 ? _field_data_T_38 : _GEN_2823; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2825 = 14'h23 == field_data_lo_18 ? _field_data_T_39 : _GEN_2824; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2826 = 14'h24 == field_data_lo_18 ? _field_data_T_40 : _GEN_2825; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2827 = 14'h25 == field_data_lo_18 ? _field_data_T_41 : _GEN_2826; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2828 = 14'h26 == field_data_lo_18 ? _field_data_T_42 : _GEN_2827; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2829 = 14'h27 == field_data_lo_18 ? _field_data_T_43 : _GEN_2828; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2830 = 14'h28 == field_data_lo_18 ? _field_data_T_44 : _GEN_2829; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2831 = 14'h29 == field_data_lo_18 ? _field_data_T_45 : _GEN_2830; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2832 = 14'h2a == field_data_lo_18 ? _field_data_T_46 : _GEN_2831; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2833 = 14'h2b == field_data_lo_18 ? _field_data_T_47 : _GEN_2832; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2834 = 14'h2c == field_data_lo_18 ? _field_data_T_48 : _GEN_2833; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2835 = 14'h2d == field_data_lo_18 ? _field_data_T_49 : _GEN_2834; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2836 = 14'h2e == field_data_lo_18 ? _field_data_T_50 : _GEN_2835; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2837 = 14'h2f == field_data_lo_18 ? _field_data_T_51 : _GEN_2836; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2838 = 14'h30 == field_data_lo_18 ? _field_data_T_52 : _GEN_2837; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2839 = 14'h31 == field_data_lo_18 ? _field_data_T_53 : _GEN_2838; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2840 = 14'h32 == field_data_lo_18 ? _field_data_T_54 : _GEN_2839; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2841 = 14'h33 == field_data_lo_18 ? _field_data_T_55 : _GEN_2840; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2842 = 14'h34 == field_data_lo_18 ? _field_data_T_56 : _GEN_2841; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2843 = 14'h35 == field_data_lo_18 ? _field_data_T_57 : _GEN_2842; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2844 = 14'h36 == field_data_lo_18 ? _field_data_T_58 : _GEN_2843; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2845 = 14'h37 == field_data_lo_18 ? _field_data_T_59 : _GEN_2844; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2846 = 14'h38 == field_data_lo_18 ? _field_data_T_60 : _GEN_2845; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2847 = 14'h39 == field_data_lo_18 ? _field_data_T_61 : _GEN_2846; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2848 = 14'h3a == field_data_lo_18 ? _field_data_T_62 : _GEN_2847; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2849 = 14'h3b == field_data_lo_18 ? _field_data_T_63 : _GEN_2848; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2850 = 14'h3c == field_data_lo_18 ? _field_data_T_64 : _GEN_2849; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2851 = 14'h3d == field_data_lo_18 ? _field_data_T_65 : _GEN_2850; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2852 = 14'h3e == field_data_lo_18 ? _field_data_T_66 : _GEN_2851; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2853 = 14'h3f == field_data_lo_18 ? _field_data_T_67 : _GEN_2852; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2854 = 14'h40 == field_data_lo_18 ? _field_data_T_68 : _GEN_2853; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2855 = 14'h41 == field_data_lo_18 ? _field_data_T_69 : _GEN_2854; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2856 = 14'h42 == field_data_lo_18 ? _field_data_T_70 : _GEN_2855; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2857 = 14'h43 == field_data_lo_18 ? _field_data_T_71 : _GEN_2856; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2858 = 14'h44 == field_data_lo_18 ? _field_data_T_72 : _GEN_2857; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2859 = 14'h45 == field_data_lo_18 ? _field_data_T_73 : _GEN_2858; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2860 = 14'h46 == field_data_lo_18 ? _field_data_T_74 : _GEN_2859; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2861 = 14'h47 == field_data_lo_18 ? _field_data_T_75 : _GEN_2860; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2862 = 14'h48 == field_data_lo_18 ? _field_data_T_76 : _GEN_2861; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2863 = 14'h49 == field_data_lo_18 ? _field_data_T_77 : _GEN_2862; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2864 = 14'h4a == field_data_lo_18 ? _field_data_T_78 : _GEN_2863; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2865 = 14'h4b == field_data_lo_18 ? _field_data_T_79 : _GEN_2864; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2866 = 14'h4c == field_data_lo_18 ? _field_data_T_80 : _GEN_2865; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2867 = 14'h4d == field_data_lo_18 ? _field_data_T_81 : _GEN_2866; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2868 = 14'h4e == field_data_lo_18 ? _field_data_T_82 : _GEN_2867; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2869 = 14'h4f == field_data_lo_18 ? _field_data_T_83 : _GEN_2868; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_51 = vliw_51[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_19 = vliw_51[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_51 = field_data_lo_19[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_51 = field_data_lo_19[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_70 = {{1'd0}, args_offset_51}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_70 = _total_offset_T_70[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2873 = 3'h1 == total_offset_70 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2874 = 3'h2 == total_offset_70 ? args_2 : _GEN_2873; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2875 = 3'h3 == total_offset_70 ? args_3 : _GEN_2874; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2876 = 3'h4 == total_offset_70 ? args_4 : _GEN_2875; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2877 = 3'h5 == total_offset_70 ? args_5 : _GEN_2876; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2878 = 3'h6 == total_offset_70 ? args_6 : _GEN_2877; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2879 = total_offset_70 < 3'h7 ? _GEN_2878 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_51_1 = 3'h0 < args_length_51 ? _GEN_2879 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_71 = args_offset_51 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2882 = 3'h1 == total_offset_71 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2883 = 3'h2 == total_offset_71 ? args_2 : _GEN_2882; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2884 = 3'h3 == total_offset_71 ? args_3 : _GEN_2883; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2885 = 3'h4 == total_offset_71 ? args_4 : _GEN_2884; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2886 = 3'h5 == total_offset_71 ? args_5 : _GEN_2885; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2887 = 3'h6 == total_offset_71 ? args_6 : _GEN_2886; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2888 = total_offset_71 < 3'h7 ? _GEN_2887 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_51_0 = 3'h1 < args_length_51 ? _GEN_2888 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1020 = {field_bytes_51_0,field_bytes_51_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2890 = opcode_51 == 4'ha ? _field_data_T_1020 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2891 = opcode_51 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2336 = opcode_51 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_19 = field_data_lo_19[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1023 = {field_data_hi_19,field_data_lo_19}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_103 = _T_2336 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2892 = opcode_51 == 4'h8 | opcode_51 == 4'hb ? _field_data_T_1023 : _GEN_2890; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2893 = opcode_51 == 4'h8 | opcode_51 == 4'hb ? _field_tag_T_103 : _GEN_2891; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2894 = 14'h20 == field_data_lo_19 ? _field_data_T_36 : _GEN_2892; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2895 = 14'h21 == field_data_lo_19 ? _field_data_T_37 : _GEN_2894; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2896 = 14'h22 == field_data_lo_19 ? _field_data_T_38 : _GEN_2895; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2897 = 14'h23 == field_data_lo_19 ? _field_data_T_39 : _GEN_2896; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2898 = 14'h24 == field_data_lo_19 ? _field_data_T_40 : _GEN_2897; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2899 = 14'h25 == field_data_lo_19 ? _field_data_T_41 : _GEN_2898; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2900 = 14'h26 == field_data_lo_19 ? _field_data_T_42 : _GEN_2899; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2901 = 14'h27 == field_data_lo_19 ? _field_data_T_43 : _GEN_2900; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2902 = 14'h28 == field_data_lo_19 ? _field_data_T_44 : _GEN_2901; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2903 = 14'h29 == field_data_lo_19 ? _field_data_T_45 : _GEN_2902; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2904 = 14'h2a == field_data_lo_19 ? _field_data_T_46 : _GEN_2903; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2905 = 14'h2b == field_data_lo_19 ? _field_data_T_47 : _GEN_2904; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2906 = 14'h2c == field_data_lo_19 ? _field_data_T_48 : _GEN_2905; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2907 = 14'h2d == field_data_lo_19 ? _field_data_T_49 : _GEN_2906; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2908 = 14'h2e == field_data_lo_19 ? _field_data_T_50 : _GEN_2907; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2909 = 14'h2f == field_data_lo_19 ? _field_data_T_51 : _GEN_2908; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2910 = 14'h30 == field_data_lo_19 ? _field_data_T_52 : _GEN_2909; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2911 = 14'h31 == field_data_lo_19 ? _field_data_T_53 : _GEN_2910; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2912 = 14'h32 == field_data_lo_19 ? _field_data_T_54 : _GEN_2911; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2913 = 14'h33 == field_data_lo_19 ? _field_data_T_55 : _GEN_2912; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2914 = 14'h34 == field_data_lo_19 ? _field_data_T_56 : _GEN_2913; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2915 = 14'h35 == field_data_lo_19 ? _field_data_T_57 : _GEN_2914; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2916 = 14'h36 == field_data_lo_19 ? _field_data_T_58 : _GEN_2915; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2917 = 14'h37 == field_data_lo_19 ? _field_data_T_59 : _GEN_2916; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2918 = 14'h38 == field_data_lo_19 ? _field_data_T_60 : _GEN_2917; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2919 = 14'h39 == field_data_lo_19 ? _field_data_T_61 : _GEN_2918; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2920 = 14'h3a == field_data_lo_19 ? _field_data_T_62 : _GEN_2919; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2921 = 14'h3b == field_data_lo_19 ? _field_data_T_63 : _GEN_2920; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2922 = 14'h3c == field_data_lo_19 ? _field_data_T_64 : _GEN_2921; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2923 = 14'h3d == field_data_lo_19 ? _field_data_T_65 : _GEN_2922; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2924 = 14'h3e == field_data_lo_19 ? _field_data_T_66 : _GEN_2923; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2925 = 14'h3f == field_data_lo_19 ? _field_data_T_67 : _GEN_2924; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2926 = 14'h40 == field_data_lo_19 ? _field_data_T_68 : _GEN_2925; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2927 = 14'h41 == field_data_lo_19 ? _field_data_T_69 : _GEN_2926; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2928 = 14'h42 == field_data_lo_19 ? _field_data_T_70 : _GEN_2927; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2929 = 14'h43 == field_data_lo_19 ? _field_data_T_71 : _GEN_2928; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2930 = 14'h44 == field_data_lo_19 ? _field_data_T_72 : _GEN_2929; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2931 = 14'h45 == field_data_lo_19 ? _field_data_T_73 : _GEN_2930; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2932 = 14'h46 == field_data_lo_19 ? _field_data_T_74 : _GEN_2931; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2933 = 14'h47 == field_data_lo_19 ? _field_data_T_75 : _GEN_2932; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2934 = 14'h48 == field_data_lo_19 ? _field_data_T_76 : _GEN_2933; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2935 = 14'h49 == field_data_lo_19 ? _field_data_T_77 : _GEN_2934; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2936 = 14'h4a == field_data_lo_19 ? _field_data_T_78 : _GEN_2935; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2937 = 14'h4b == field_data_lo_19 ? _field_data_T_79 : _GEN_2936; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2938 = 14'h4c == field_data_lo_19 ? _field_data_T_80 : _GEN_2937; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2939 = 14'h4d == field_data_lo_19 ? _field_data_T_81 : _GEN_2938; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2940 = 14'h4e == field_data_lo_19 ? _field_data_T_82 : _GEN_2939; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2941 = 14'h4f == field_data_lo_19 ? _field_data_T_83 : _GEN_2940; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_52 = vliw_52[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_20 = vliw_52[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_52 = field_data_lo_20[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_52 = field_data_lo_20[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_72 = {{1'd0}, args_offset_52}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_72 = _total_offset_T_72[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2945 = 3'h1 == total_offset_72 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2946 = 3'h2 == total_offset_72 ? args_2 : _GEN_2945; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2947 = 3'h3 == total_offset_72 ? args_3 : _GEN_2946; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2948 = 3'h4 == total_offset_72 ? args_4 : _GEN_2947; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2949 = 3'h5 == total_offset_72 ? args_5 : _GEN_2948; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2950 = 3'h6 == total_offset_72 ? args_6 : _GEN_2949; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2951 = total_offset_72 < 3'h7 ? _GEN_2950 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_52_1 = 3'h0 < args_length_52 ? _GEN_2951 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_73 = args_offset_52 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2954 = 3'h1 == total_offset_73 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2955 = 3'h2 == total_offset_73 ? args_2 : _GEN_2954; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2956 = 3'h3 == total_offset_73 ? args_3 : _GEN_2955; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2957 = 3'h4 == total_offset_73 ? args_4 : _GEN_2956; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2958 = 3'h5 == total_offset_73 ? args_5 : _GEN_2957; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2959 = 3'h6 == total_offset_73 ? args_6 : _GEN_2958; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2960 = total_offset_73 < 3'h7 ? _GEN_2959 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_52_0 = 3'h1 < args_length_52 ? _GEN_2960 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1072 = {field_bytes_52_0,field_bytes_52_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2962 = opcode_52 == 4'ha ? _field_data_T_1072 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2963 = opcode_52 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2393 = opcode_52 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_20 = field_data_lo_20[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1075 = {field_data_hi_20,field_data_lo_20}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_105 = _T_2393 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2964 = opcode_52 == 4'h8 | opcode_52 == 4'hb ? _field_data_T_1075 : _GEN_2962; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2965 = opcode_52 == 4'h8 | opcode_52 == 4'hb ? _field_tag_T_105 : _GEN_2963; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2966 = 14'h20 == field_data_lo_20 ? _field_data_T_36 : _GEN_2964; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2967 = 14'h21 == field_data_lo_20 ? _field_data_T_37 : _GEN_2966; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2968 = 14'h22 == field_data_lo_20 ? _field_data_T_38 : _GEN_2967; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2969 = 14'h23 == field_data_lo_20 ? _field_data_T_39 : _GEN_2968; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2970 = 14'h24 == field_data_lo_20 ? _field_data_T_40 : _GEN_2969; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2971 = 14'h25 == field_data_lo_20 ? _field_data_T_41 : _GEN_2970; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2972 = 14'h26 == field_data_lo_20 ? _field_data_T_42 : _GEN_2971; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2973 = 14'h27 == field_data_lo_20 ? _field_data_T_43 : _GEN_2972; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2974 = 14'h28 == field_data_lo_20 ? _field_data_T_44 : _GEN_2973; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2975 = 14'h29 == field_data_lo_20 ? _field_data_T_45 : _GEN_2974; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2976 = 14'h2a == field_data_lo_20 ? _field_data_T_46 : _GEN_2975; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2977 = 14'h2b == field_data_lo_20 ? _field_data_T_47 : _GEN_2976; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2978 = 14'h2c == field_data_lo_20 ? _field_data_T_48 : _GEN_2977; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2979 = 14'h2d == field_data_lo_20 ? _field_data_T_49 : _GEN_2978; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2980 = 14'h2e == field_data_lo_20 ? _field_data_T_50 : _GEN_2979; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2981 = 14'h2f == field_data_lo_20 ? _field_data_T_51 : _GEN_2980; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2982 = 14'h30 == field_data_lo_20 ? _field_data_T_52 : _GEN_2981; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2983 = 14'h31 == field_data_lo_20 ? _field_data_T_53 : _GEN_2982; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2984 = 14'h32 == field_data_lo_20 ? _field_data_T_54 : _GEN_2983; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2985 = 14'h33 == field_data_lo_20 ? _field_data_T_55 : _GEN_2984; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2986 = 14'h34 == field_data_lo_20 ? _field_data_T_56 : _GEN_2985; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2987 = 14'h35 == field_data_lo_20 ? _field_data_T_57 : _GEN_2986; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2988 = 14'h36 == field_data_lo_20 ? _field_data_T_58 : _GEN_2987; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2989 = 14'h37 == field_data_lo_20 ? _field_data_T_59 : _GEN_2988; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2990 = 14'h38 == field_data_lo_20 ? _field_data_T_60 : _GEN_2989; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2991 = 14'h39 == field_data_lo_20 ? _field_data_T_61 : _GEN_2990; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2992 = 14'h3a == field_data_lo_20 ? _field_data_T_62 : _GEN_2991; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2993 = 14'h3b == field_data_lo_20 ? _field_data_T_63 : _GEN_2992; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2994 = 14'h3c == field_data_lo_20 ? _field_data_T_64 : _GEN_2993; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2995 = 14'h3d == field_data_lo_20 ? _field_data_T_65 : _GEN_2994; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2996 = 14'h3e == field_data_lo_20 ? _field_data_T_66 : _GEN_2995; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2997 = 14'h3f == field_data_lo_20 ? _field_data_T_67 : _GEN_2996; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2998 = 14'h40 == field_data_lo_20 ? _field_data_T_68 : _GEN_2997; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2999 = 14'h41 == field_data_lo_20 ? _field_data_T_69 : _GEN_2998; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3000 = 14'h42 == field_data_lo_20 ? _field_data_T_70 : _GEN_2999; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3001 = 14'h43 == field_data_lo_20 ? _field_data_T_71 : _GEN_3000; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3002 = 14'h44 == field_data_lo_20 ? _field_data_T_72 : _GEN_3001; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3003 = 14'h45 == field_data_lo_20 ? _field_data_T_73 : _GEN_3002; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3004 = 14'h46 == field_data_lo_20 ? _field_data_T_74 : _GEN_3003; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3005 = 14'h47 == field_data_lo_20 ? _field_data_T_75 : _GEN_3004; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3006 = 14'h48 == field_data_lo_20 ? _field_data_T_76 : _GEN_3005; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3007 = 14'h49 == field_data_lo_20 ? _field_data_T_77 : _GEN_3006; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3008 = 14'h4a == field_data_lo_20 ? _field_data_T_78 : _GEN_3007; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3009 = 14'h4b == field_data_lo_20 ? _field_data_T_79 : _GEN_3008; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3010 = 14'h4c == field_data_lo_20 ? _field_data_T_80 : _GEN_3009; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3011 = 14'h4d == field_data_lo_20 ? _field_data_T_81 : _GEN_3010; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3012 = 14'h4e == field_data_lo_20 ? _field_data_T_82 : _GEN_3011; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3013 = 14'h4f == field_data_lo_20 ? _field_data_T_83 : _GEN_3012; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_53 = vliw_53[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_21 = vliw_53[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_53 = field_data_lo_21[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_53 = field_data_lo_21[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_74 = {{1'd0}, args_offset_53}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_74 = _total_offset_T_74[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3017 = 3'h1 == total_offset_74 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3018 = 3'h2 == total_offset_74 ? args_2 : _GEN_3017; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3019 = 3'h3 == total_offset_74 ? args_3 : _GEN_3018; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3020 = 3'h4 == total_offset_74 ? args_4 : _GEN_3019; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3021 = 3'h5 == total_offset_74 ? args_5 : _GEN_3020; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3022 = 3'h6 == total_offset_74 ? args_6 : _GEN_3021; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3023 = total_offset_74 < 3'h7 ? _GEN_3022 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_53_1 = 3'h0 < args_length_53 ? _GEN_3023 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_75 = args_offset_53 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3026 = 3'h1 == total_offset_75 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3027 = 3'h2 == total_offset_75 ? args_2 : _GEN_3026; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3028 = 3'h3 == total_offset_75 ? args_3 : _GEN_3027; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3029 = 3'h4 == total_offset_75 ? args_4 : _GEN_3028; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3030 = 3'h5 == total_offset_75 ? args_5 : _GEN_3029; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3031 = 3'h6 == total_offset_75 ? args_6 : _GEN_3030; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3032 = total_offset_75 < 3'h7 ? _GEN_3031 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_53_0 = 3'h1 < args_length_53 ? _GEN_3032 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1124 = {field_bytes_53_0,field_bytes_53_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_3034 = opcode_53 == 4'ha ? _field_data_T_1124 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3035 = opcode_53 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2450 = opcode_53 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_21 = field_data_lo_21[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1127 = {field_data_hi_21,field_data_lo_21}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_107 = _T_2450 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_3036 = opcode_53 == 4'h8 | opcode_53 == 4'hb ? _field_data_T_1127 : _GEN_3034; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3037 = opcode_53 == 4'h8 | opcode_53 == 4'hb ? _field_tag_T_107 : _GEN_3035; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_3038 = 14'h20 == field_data_lo_21 ? _field_data_T_36 : _GEN_3036; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3039 = 14'h21 == field_data_lo_21 ? _field_data_T_37 : _GEN_3038; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3040 = 14'h22 == field_data_lo_21 ? _field_data_T_38 : _GEN_3039; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3041 = 14'h23 == field_data_lo_21 ? _field_data_T_39 : _GEN_3040; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3042 = 14'h24 == field_data_lo_21 ? _field_data_T_40 : _GEN_3041; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3043 = 14'h25 == field_data_lo_21 ? _field_data_T_41 : _GEN_3042; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3044 = 14'h26 == field_data_lo_21 ? _field_data_T_42 : _GEN_3043; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3045 = 14'h27 == field_data_lo_21 ? _field_data_T_43 : _GEN_3044; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3046 = 14'h28 == field_data_lo_21 ? _field_data_T_44 : _GEN_3045; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3047 = 14'h29 == field_data_lo_21 ? _field_data_T_45 : _GEN_3046; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3048 = 14'h2a == field_data_lo_21 ? _field_data_T_46 : _GEN_3047; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3049 = 14'h2b == field_data_lo_21 ? _field_data_T_47 : _GEN_3048; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3050 = 14'h2c == field_data_lo_21 ? _field_data_T_48 : _GEN_3049; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3051 = 14'h2d == field_data_lo_21 ? _field_data_T_49 : _GEN_3050; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3052 = 14'h2e == field_data_lo_21 ? _field_data_T_50 : _GEN_3051; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3053 = 14'h2f == field_data_lo_21 ? _field_data_T_51 : _GEN_3052; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3054 = 14'h30 == field_data_lo_21 ? _field_data_T_52 : _GEN_3053; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3055 = 14'h31 == field_data_lo_21 ? _field_data_T_53 : _GEN_3054; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3056 = 14'h32 == field_data_lo_21 ? _field_data_T_54 : _GEN_3055; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3057 = 14'h33 == field_data_lo_21 ? _field_data_T_55 : _GEN_3056; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3058 = 14'h34 == field_data_lo_21 ? _field_data_T_56 : _GEN_3057; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3059 = 14'h35 == field_data_lo_21 ? _field_data_T_57 : _GEN_3058; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3060 = 14'h36 == field_data_lo_21 ? _field_data_T_58 : _GEN_3059; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3061 = 14'h37 == field_data_lo_21 ? _field_data_T_59 : _GEN_3060; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3062 = 14'h38 == field_data_lo_21 ? _field_data_T_60 : _GEN_3061; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3063 = 14'h39 == field_data_lo_21 ? _field_data_T_61 : _GEN_3062; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3064 = 14'h3a == field_data_lo_21 ? _field_data_T_62 : _GEN_3063; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3065 = 14'h3b == field_data_lo_21 ? _field_data_T_63 : _GEN_3064; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3066 = 14'h3c == field_data_lo_21 ? _field_data_T_64 : _GEN_3065; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3067 = 14'h3d == field_data_lo_21 ? _field_data_T_65 : _GEN_3066; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3068 = 14'h3e == field_data_lo_21 ? _field_data_T_66 : _GEN_3067; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3069 = 14'h3f == field_data_lo_21 ? _field_data_T_67 : _GEN_3068; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3070 = 14'h40 == field_data_lo_21 ? _field_data_T_68 : _GEN_3069; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3071 = 14'h41 == field_data_lo_21 ? _field_data_T_69 : _GEN_3070; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3072 = 14'h42 == field_data_lo_21 ? _field_data_T_70 : _GEN_3071; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3073 = 14'h43 == field_data_lo_21 ? _field_data_T_71 : _GEN_3072; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3074 = 14'h44 == field_data_lo_21 ? _field_data_T_72 : _GEN_3073; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3075 = 14'h45 == field_data_lo_21 ? _field_data_T_73 : _GEN_3074; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3076 = 14'h46 == field_data_lo_21 ? _field_data_T_74 : _GEN_3075; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3077 = 14'h47 == field_data_lo_21 ? _field_data_T_75 : _GEN_3076; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3078 = 14'h48 == field_data_lo_21 ? _field_data_T_76 : _GEN_3077; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3079 = 14'h49 == field_data_lo_21 ? _field_data_T_77 : _GEN_3078; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3080 = 14'h4a == field_data_lo_21 ? _field_data_T_78 : _GEN_3079; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3081 = 14'h4b == field_data_lo_21 ? _field_data_T_79 : _GEN_3080; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3082 = 14'h4c == field_data_lo_21 ? _field_data_T_80 : _GEN_3081; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3083 = 14'h4d == field_data_lo_21 ? _field_data_T_81 : _GEN_3082; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3084 = 14'h4e == field_data_lo_21 ? _field_data_T_82 : _GEN_3083; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3085 = 14'h4f == field_data_lo_21 ? _field_data_T_83 : _GEN_3084; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_54 = vliw_54[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_22 = vliw_54[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_54 = field_data_lo_22[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_54 = field_data_lo_22[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_76 = {{1'd0}, args_offset_54}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_76 = _total_offset_T_76[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3089 = 3'h1 == total_offset_76 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3090 = 3'h2 == total_offset_76 ? args_2 : _GEN_3089; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3091 = 3'h3 == total_offset_76 ? args_3 : _GEN_3090; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3092 = 3'h4 == total_offset_76 ? args_4 : _GEN_3091; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3093 = 3'h5 == total_offset_76 ? args_5 : _GEN_3092; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3094 = 3'h6 == total_offset_76 ? args_6 : _GEN_3093; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3095 = total_offset_76 < 3'h7 ? _GEN_3094 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_54_1 = 3'h0 < args_length_54 ? _GEN_3095 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_77 = args_offset_54 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3098 = 3'h1 == total_offset_77 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3099 = 3'h2 == total_offset_77 ? args_2 : _GEN_3098; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3100 = 3'h3 == total_offset_77 ? args_3 : _GEN_3099; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3101 = 3'h4 == total_offset_77 ? args_4 : _GEN_3100; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3102 = 3'h5 == total_offset_77 ? args_5 : _GEN_3101; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3103 = 3'h6 == total_offset_77 ? args_6 : _GEN_3102; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3104 = total_offset_77 < 3'h7 ? _GEN_3103 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_54_0 = 3'h1 < args_length_54 ? _GEN_3104 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1176 = {field_bytes_54_0,field_bytes_54_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_3106 = opcode_54 == 4'ha ? _field_data_T_1176 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3107 = opcode_54 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2507 = opcode_54 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_22 = field_data_lo_22[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1179 = {field_data_hi_22,field_data_lo_22}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_109 = _T_2507 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_3108 = opcode_54 == 4'h8 | opcode_54 == 4'hb ? _field_data_T_1179 : _GEN_3106; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3109 = opcode_54 == 4'h8 | opcode_54 == 4'hb ? _field_tag_T_109 : _GEN_3107; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_3110 = 14'h20 == field_data_lo_22 ? _field_data_T_36 : _GEN_3108; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3111 = 14'h21 == field_data_lo_22 ? _field_data_T_37 : _GEN_3110; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3112 = 14'h22 == field_data_lo_22 ? _field_data_T_38 : _GEN_3111; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3113 = 14'h23 == field_data_lo_22 ? _field_data_T_39 : _GEN_3112; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3114 = 14'h24 == field_data_lo_22 ? _field_data_T_40 : _GEN_3113; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3115 = 14'h25 == field_data_lo_22 ? _field_data_T_41 : _GEN_3114; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3116 = 14'h26 == field_data_lo_22 ? _field_data_T_42 : _GEN_3115; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3117 = 14'h27 == field_data_lo_22 ? _field_data_T_43 : _GEN_3116; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3118 = 14'h28 == field_data_lo_22 ? _field_data_T_44 : _GEN_3117; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3119 = 14'h29 == field_data_lo_22 ? _field_data_T_45 : _GEN_3118; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3120 = 14'h2a == field_data_lo_22 ? _field_data_T_46 : _GEN_3119; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3121 = 14'h2b == field_data_lo_22 ? _field_data_T_47 : _GEN_3120; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3122 = 14'h2c == field_data_lo_22 ? _field_data_T_48 : _GEN_3121; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3123 = 14'h2d == field_data_lo_22 ? _field_data_T_49 : _GEN_3122; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3124 = 14'h2e == field_data_lo_22 ? _field_data_T_50 : _GEN_3123; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3125 = 14'h2f == field_data_lo_22 ? _field_data_T_51 : _GEN_3124; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3126 = 14'h30 == field_data_lo_22 ? _field_data_T_52 : _GEN_3125; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3127 = 14'h31 == field_data_lo_22 ? _field_data_T_53 : _GEN_3126; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3128 = 14'h32 == field_data_lo_22 ? _field_data_T_54 : _GEN_3127; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3129 = 14'h33 == field_data_lo_22 ? _field_data_T_55 : _GEN_3128; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3130 = 14'h34 == field_data_lo_22 ? _field_data_T_56 : _GEN_3129; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3131 = 14'h35 == field_data_lo_22 ? _field_data_T_57 : _GEN_3130; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3132 = 14'h36 == field_data_lo_22 ? _field_data_T_58 : _GEN_3131; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3133 = 14'h37 == field_data_lo_22 ? _field_data_T_59 : _GEN_3132; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3134 = 14'h38 == field_data_lo_22 ? _field_data_T_60 : _GEN_3133; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3135 = 14'h39 == field_data_lo_22 ? _field_data_T_61 : _GEN_3134; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3136 = 14'h3a == field_data_lo_22 ? _field_data_T_62 : _GEN_3135; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3137 = 14'h3b == field_data_lo_22 ? _field_data_T_63 : _GEN_3136; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3138 = 14'h3c == field_data_lo_22 ? _field_data_T_64 : _GEN_3137; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3139 = 14'h3d == field_data_lo_22 ? _field_data_T_65 : _GEN_3138; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3140 = 14'h3e == field_data_lo_22 ? _field_data_T_66 : _GEN_3139; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3141 = 14'h3f == field_data_lo_22 ? _field_data_T_67 : _GEN_3140; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3142 = 14'h40 == field_data_lo_22 ? _field_data_T_68 : _GEN_3141; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3143 = 14'h41 == field_data_lo_22 ? _field_data_T_69 : _GEN_3142; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3144 = 14'h42 == field_data_lo_22 ? _field_data_T_70 : _GEN_3143; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3145 = 14'h43 == field_data_lo_22 ? _field_data_T_71 : _GEN_3144; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3146 = 14'h44 == field_data_lo_22 ? _field_data_T_72 : _GEN_3145; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3147 = 14'h45 == field_data_lo_22 ? _field_data_T_73 : _GEN_3146; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3148 = 14'h46 == field_data_lo_22 ? _field_data_T_74 : _GEN_3147; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3149 = 14'h47 == field_data_lo_22 ? _field_data_T_75 : _GEN_3148; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3150 = 14'h48 == field_data_lo_22 ? _field_data_T_76 : _GEN_3149; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3151 = 14'h49 == field_data_lo_22 ? _field_data_T_77 : _GEN_3150; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3152 = 14'h4a == field_data_lo_22 ? _field_data_T_78 : _GEN_3151; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3153 = 14'h4b == field_data_lo_22 ? _field_data_T_79 : _GEN_3152; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3154 = 14'h4c == field_data_lo_22 ? _field_data_T_80 : _GEN_3153; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3155 = 14'h4d == field_data_lo_22 ? _field_data_T_81 : _GEN_3154; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3156 = 14'h4e == field_data_lo_22 ? _field_data_T_82 : _GEN_3155; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3157 = 14'h4f == field_data_lo_22 ? _field_data_T_83 : _GEN_3156; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_55 = vliw_55[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_23 = vliw_55[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_55 = field_data_lo_23[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_55 = field_data_lo_23[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_78 = {{1'd0}, args_offset_55}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_78 = _total_offset_T_78[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3161 = 3'h1 == total_offset_78 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3162 = 3'h2 == total_offset_78 ? args_2 : _GEN_3161; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3163 = 3'h3 == total_offset_78 ? args_3 : _GEN_3162; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3164 = 3'h4 == total_offset_78 ? args_4 : _GEN_3163; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3165 = 3'h5 == total_offset_78 ? args_5 : _GEN_3164; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3166 = 3'h6 == total_offset_78 ? args_6 : _GEN_3165; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3167 = total_offset_78 < 3'h7 ? _GEN_3166 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_55_1 = 3'h0 < args_length_55 ? _GEN_3167 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_79 = args_offset_55 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3170 = 3'h1 == total_offset_79 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3171 = 3'h2 == total_offset_79 ? args_2 : _GEN_3170; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3172 = 3'h3 == total_offset_79 ? args_3 : _GEN_3171; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3173 = 3'h4 == total_offset_79 ? args_4 : _GEN_3172; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3174 = 3'h5 == total_offset_79 ? args_5 : _GEN_3173; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3175 = 3'h6 == total_offset_79 ? args_6 : _GEN_3174; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3176 = total_offset_79 < 3'h7 ? _GEN_3175 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_55_0 = 3'h1 < args_length_55 ? _GEN_3176 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1228 = {field_bytes_55_0,field_bytes_55_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_3178 = opcode_55 == 4'ha ? _field_data_T_1228 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3179 = opcode_55 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2564 = opcode_55 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_23 = field_data_lo_23[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1231 = {field_data_hi_23,field_data_lo_23}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_111 = _T_2564 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_3180 = opcode_55 == 4'h8 | opcode_55 == 4'hb ? _field_data_T_1231 : _GEN_3178; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3181 = opcode_55 == 4'h8 | opcode_55 == 4'hb ? _field_tag_T_111 : _GEN_3179; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_3182 = 14'h20 == field_data_lo_23 ? _field_data_T_36 : _GEN_3180; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3183 = 14'h21 == field_data_lo_23 ? _field_data_T_37 : _GEN_3182; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3184 = 14'h22 == field_data_lo_23 ? _field_data_T_38 : _GEN_3183; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3185 = 14'h23 == field_data_lo_23 ? _field_data_T_39 : _GEN_3184; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3186 = 14'h24 == field_data_lo_23 ? _field_data_T_40 : _GEN_3185; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3187 = 14'h25 == field_data_lo_23 ? _field_data_T_41 : _GEN_3186; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3188 = 14'h26 == field_data_lo_23 ? _field_data_T_42 : _GEN_3187; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3189 = 14'h27 == field_data_lo_23 ? _field_data_T_43 : _GEN_3188; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3190 = 14'h28 == field_data_lo_23 ? _field_data_T_44 : _GEN_3189; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3191 = 14'h29 == field_data_lo_23 ? _field_data_T_45 : _GEN_3190; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3192 = 14'h2a == field_data_lo_23 ? _field_data_T_46 : _GEN_3191; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3193 = 14'h2b == field_data_lo_23 ? _field_data_T_47 : _GEN_3192; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3194 = 14'h2c == field_data_lo_23 ? _field_data_T_48 : _GEN_3193; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3195 = 14'h2d == field_data_lo_23 ? _field_data_T_49 : _GEN_3194; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3196 = 14'h2e == field_data_lo_23 ? _field_data_T_50 : _GEN_3195; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3197 = 14'h2f == field_data_lo_23 ? _field_data_T_51 : _GEN_3196; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3198 = 14'h30 == field_data_lo_23 ? _field_data_T_52 : _GEN_3197; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3199 = 14'h31 == field_data_lo_23 ? _field_data_T_53 : _GEN_3198; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3200 = 14'h32 == field_data_lo_23 ? _field_data_T_54 : _GEN_3199; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3201 = 14'h33 == field_data_lo_23 ? _field_data_T_55 : _GEN_3200; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3202 = 14'h34 == field_data_lo_23 ? _field_data_T_56 : _GEN_3201; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3203 = 14'h35 == field_data_lo_23 ? _field_data_T_57 : _GEN_3202; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3204 = 14'h36 == field_data_lo_23 ? _field_data_T_58 : _GEN_3203; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3205 = 14'h37 == field_data_lo_23 ? _field_data_T_59 : _GEN_3204; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3206 = 14'h38 == field_data_lo_23 ? _field_data_T_60 : _GEN_3205; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3207 = 14'h39 == field_data_lo_23 ? _field_data_T_61 : _GEN_3206; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3208 = 14'h3a == field_data_lo_23 ? _field_data_T_62 : _GEN_3207; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3209 = 14'h3b == field_data_lo_23 ? _field_data_T_63 : _GEN_3208; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3210 = 14'h3c == field_data_lo_23 ? _field_data_T_64 : _GEN_3209; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3211 = 14'h3d == field_data_lo_23 ? _field_data_T_65 : _GEN_3210; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3212 = 14'h3e == field_data_lo_23 ? _field_data_T_66 : _GEN_3211; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3213 = 14'h3f == field_data_lo_23 ? _field_data_T_67 : _GEN_3212; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3214 = 14'h40 == field_data_lo_23 ? _field_data_T_68 : _GEN_3213; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3215 = 14'h41 == field_data_lo_23 ? _field_data_T_69 : _GEN_3214; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3216 = 14'h42 == field_data_lo_23 ? _field_data_T_70 : _GEN_3215; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3217 = 14'h43 == field_data_lo_23 ? _field_data_T_71 : _GEN_3216; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3218 = 14'h44 == field_data_lo_23 ? _field_data_T_72 : _GEN_3217; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3219 = 14'h45 == field_data_lo_23 ? _field_data_T_73 : _GEN_3218; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3220 = 14'h46 == field_data_lo_23 ? _field_data_T_74 : _GEN_3219; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3221 = 14'h47 == field_data_lo_23 ? _field_data_T_75 : _GEN_3220; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3222 = 14'h48 == field_data_lo_23 ? _field_data_T_76 : _GEN_3221; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3223 = 14'h49 == field_data_lo_23 ? _field_data_T_77 : _GEN_3222; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3224 = 14'h4a == field_data_lo_23 ? _field_data_T_78 : _GEN_3223; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3225 = 14'h4b == field_data_lo_23 ? _field_data_T_79 : _GEN_3224; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3226 = 14'h4c == field_data_lo_23 ? _field_data_T_80 : _GEN_3225; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3227 = 14'h4d == field_data_lo_23 ? _field_data_T_81 : _GEN_3226; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3228 = 14'h4e == field_data_lo_23 ? _field_data_T_82 : _GEN_3227; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3229 = 14'h4f == field_data_lo_23 ? _field_data_T_83 : _GEN_3228; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_56 = vliw_56[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_24 = vliw_56[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_56 = field_data_lo_24[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_56 = field_data_lo_24[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_80 = {{1'd0}, args_offset_56}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_80 = _total_offset_T_80[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3233 = 3'h1 == total_offset_80 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3234 = 3'h2 == total_offset_80 ? args_2 : _GEN_3233; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3235 = 3'h3 == total_offset_80 ? args_3 : _GEN_3234; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3236 = 3'h4 == total_offset_80 ? args_4 : _GEN_3235; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3237 = 3'h5 == total_offset_80 ? args_5 : _GEN_3236; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3238 = 3'h6 == total_offset_80 ? args_6 : _GEN_3237; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3239 = total_offset_80 < 3'h7 ? _GEN_3238 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_56_1 = 3'h0 < args_length_56 ? _GEN_3239 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_81 = args_offset_56 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3242 = 3'h1 == total_offset_81 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3243 = 3'h2 == total_offset_81 ? args_2 : _GEN_3242; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3244 = 3'h3 == total_offset_81 ? args_3 : _GEN_3243; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3245 = 3'h4 == total_offset_81 ? args_4 : _GEN_3244; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3246 = 3'h5 == total_offset_81 ? args_5 : _GEN_3245; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3247 = 3'h6 == total_offset_81 ? args_6 : _GEN_3246; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3248 = total_offset_81 < 3'h7 ? _GEN_3247 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_56_0 = 3'h1 < args_length_56 ? _GEN_3248 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1280 = {field_bytes_56_0,field_bytes_56_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_3250 = opcode_56 == 4'ha ? _field_data_T_1280 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3251 = opcode_56 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2621 = opcode_56 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_24 = field_data_lo_24[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1283 = {field_data_hi_24,field_data_lo_24}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_113 = _T_2621 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_3252 = opcode_56 == 4'h8 | opcode_56 == 4'hb ? _field_data_T_1283 : _GEN_3250; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3253 = opcode_56 == 4'h8 | opcode_56 == 4'hb ? _field_tag_T_113 : _GEN_3251; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_3254 = 14'h20 == field_data_lo_24 ? _field_data_T_36 : _GEN_3252; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3255 = 14'h21 == field_data_lo_24 ? _field_data_T_37 : _GEN_3254; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3256 = 14'h22 == field_data_lo_24 ? _field_data_T_38 : _GEN_3255; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3257 = 14'h23 == field_data_lo_24 ? _field_data_T_39 : _GEN_3256; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3258 = 14'h24 == field_data_lo_24 ? _field_data_T_40 : _GEN_3257; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3259 = 14'h25 == field_data_lo_24 ? _field_data_T_41 : _GEN_3258; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3260 = 14'h26 == field_data_lo_24 ? _field_data_T_42 : _GEN_3259; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3261 = 14'h27 == field_data_lo_24 ? _field_data_T_43 : _GEN_3260; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3262 = 14'h28 == field_data_lo_24 ? _field_data_T_44 : _GEN_3261; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3263 = 14'h29 == field_data_lo_24 ? _field_data_T_45 : _GEN_3262; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3264 = 14'h2a == field_data_lo_24 ? _field_data_T_46 : _GEN_3263; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3265 = 14'h2b == field_data_lo_24 ? _field_data_T_47 : _GEN_3264; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3266 = 14'h2c == field_data_lo_24 ? _field_data_T_48 : _GEN_3265; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3267 = 14'h2d == field_data_lo_24 ? _field_data_T_49 : _GEN_3266; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3268 = 14'h2e == field_data_lo_24 ? _field_data_T_50 : _GEN_3267; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3269 = 14'h2f == field_data_lo_24 ? _field_data_T_51 : _GEN_3268; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3270 = 14'h30 == field_data_lo_24 ? _field_data_T_52 : _GEN_3269; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3271 = 14'h31 == field_data_lo_24 ? _field_data_T_53 : _GEN_3270; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3272 = 14'h32 == field_data_lo_24 ? _field_data_T_54 : _GEN_3271; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3273 = 14'h33 == field_data_lo_24 ? _field_data_T_55 : _GEN_3272; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3274 = 14'h34 == field_data_lo_24 ? _field_data_T_56 : _GEN_3273; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3275 = 14'h35 == field_data_lo_24 ? _field_data_T_57 : _GEN_3274; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3276 = 14'h36 == field_data_lo_24 ? _field_data_T_58 : _GEN_3275; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3277 = 14'h37 == field_data_lo_24 ? _field_data_T_59 : _GEN_3276; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3278 = 14'h38 == field_data_lo_24 ? _field_data_T_60 : _GEN_3277; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3279 = 14'h39 == field_data_lo_24 ? _field_data_T_61 : _GEN_3278; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3280 = 14'h3a == field_data_lo_24 ? _field_data_T_62 : _GEN_3279; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3281 = 14'h3b == field_data_lo_24 ? _field_data_T_63 : _GEN_3280; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3282 = 14'h3c == field_data_lo_24 ? _field_data_T_64 : _GEN_3281; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3283 = 14'h3d == field_data_lo_24 ? _field_data_T_65 : _GEN_3282; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3284 = 14'h3e == field_data_lo_24 ? _field_data_T_66 : _GEN_3283; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3285 = 14'h3f == field_data_lo_24 ? _field_data_T_67 : _GEN_3284; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3286 = 14'h40 == field_data_lo_24 ? _field_data_T_68 : _GEN_3285; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3287 = 14'h41 == field_data_lo_24 ? _field_data_T_69 : _GEN_3286; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3288 = 14'h42 == field_data_lo_24 ? _field_data_T_70 : _GEN_3287; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3289 = 14'h43 == field_data_lo_24 ? _field_data_T_71 : _GEN_3288; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3290 = 14'h44 == field_data_lo_24 ? _field_data_T_72 : _GEN_3289; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3291 = 14'h45 == field_data_lo_24 ? _field_data_T_73 : _GEN_3290; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3292 = 14'h46 == field_data_lo_24 ? _field_data_T_74 : _GEN_3291; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3293 = 14'h47 == field_data_lo_24 ? _field_data_T_75 : _GEN_3292; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3294 = 14'h48 == field_data_lo_24 ? _field_data_T_76 : _GEN_3293; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3295 = 14'h49 == field_data_lo_24 ? _field_data_T_77 : _GEN_3294; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3296 = 14'h4a == field_data_lo_24 ? _field_data_T_78 : _GEN_3295; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3297 = 14'h4b == field_data_lo_24 ? _field_data_T_79 : _GEN_3296; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3298 = 14'h4c == field_data_lo_24 ? _field_data_T_80 : _GEN_3297; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3299 = 14'h4d == field_data_lo_24 ? _field_data_T_81 : _GEN_3298; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3300 = 14'h4e == field_data_lo_24 ? _field_data_T_82 : _GEN_3299; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3301 = 14'h4f == field_data_lo_24 ? _field_data_T_83 : _GEN_3300; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_57 = vliw_57[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_25 = vliw_57[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_57 = field_data_lo_25[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_57 = field_data_lo_25[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_82 = {{1'd0}, args_offset_57}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_82 = _total_offset_T_82[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3305 = 3'h1 == total_offset_82 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3306 = 3'h2 == total_offset_82 ? args_2 : _GEN_3305; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3307 = 3'h3 == total_offset_82 ? args_3 : _GEN_3306; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3308 = 3'h4 == total_offset_82 ? args_4 : _GEN_3307; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3309 = 3'h5 == total_offset_82 ? args_5 : _GEN_3308; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3310 = 3'h6 == total_offset_82 ? args_6 : _GEN_3309; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3311 = total_offset_82 < 3'h7 ? _GEN_3310 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_57_1 = 3'h0 < args_length_57 ? _GEN_3311 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_83 = args_offset_57 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3314 = 3'h1 == total_offset_83 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3315 = 3'h2 == total_offset_83 ? args_2 : _GEN_3314; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3316 = 3'h3 == total_offset_83 ? args_3 : _GEN_3315; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3317 = 3'h4 == total_offset_83 ? args_4 : _GEN_3316; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3318 = 3'h5 == total_offset_83 ? args_5 : _GEN_3317; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3319 = 3'h6 == total_offset_83 ? args_6 : _GEN_3318; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3320 = total_offset_83 < 3'h7 ? _GEN_3319 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_57_0 = 3'h1 < args_length_57 ? _GEN_3320 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1332 = {field_bytes_57_0,field_bytes_57_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_3322 = opcode_57 == 4'ha ? _field_data_T_1332 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3323 = opcode_57 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2678 = opcode_57 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_25 = field_data_lo_25[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1335 = {field_data_hi_25,field_data_lo_25}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_115 = _T_2678 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_3324 = opcode_57 == 4'h8 | opcode_57 == 4'hb ? _field_data_T_1335 : _GEN_3322; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3325 = opcode_57 == 4'h8 | opcode_57 == 4'hb ? _field_tag_T_115 : _GEN_3323; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_3326 = 14'h20 == field_data_lo_25 ? _field_data_T_36 : _GEN_3324; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3327 = 14'h21 == field_data_lo_25 ? _field_data_T_37 : _GEN_3326; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3328 = 14'h22 == field_data_lo_25 ? _field_data_T_38 : _GEN_3327; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3329 = 14'h23 == field_data_lo_25 ? _field_data_T_39 : _GEN_3328; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3330 = 14'h24 == field_data_lo_25 ? _field_data_T_40 : _GEN_3329; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3331 = 14'h25 == field_data_lo_25 ? _field_data_T_41 : _GEN_3330; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3332 = 14'h26 == field_data_lo_25 ? _field_data_T_42 : _GEN_3331; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3333 = 14'h27 == field_data_lo_25 ? _field_data_T_43 : _GEN_3332; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3334 = 14'h28 == field_data_lo_25 ? _field_data_T_44 : _GEN_3333; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3335 = 14'h29 == field_data_lo_25 ? _field_data_T_45 : _GEN_3334; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3336 = 14'h2a == field_data_lo_25 ? _field_data_T_46 : _GEN_3335; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3337 = 14'h2b == field_data_lo_25 ? _field_data_T_47 : _GEN_3336; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3338 = 14'h2c == field_data_lo_25 ? _field_data_T_48 : _GEN_3337; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3339 = 14'h2d == field_data_lo_25 ? _field_data_T_49 : _GEN_3338; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3340 = 14'h2e == field_data_lo_25 ? _field_data_T_50 : _GEN_3339; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3341 = 14'h2f == field_data_lo_25 ? _field_data_T_51 : _GEN_3340; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3342 = 14'h30 == field_data_lo_25 ? _field_data_T_52 : _GEN_3341; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3343 = 14'h31 == field_data_lo_25 ? _field_data_T_53 : _GEN_3342; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3344 = 14'h32 == field_data_lo_25 ? _field_data_T_54 : _GEN_3343; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3345 = 14'h33 == field_data_lo_25 ? _field_data_T_55 : _GEN_3344; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3346 = 14'h34 == field_data_lo_25 ? _field_data_T_56 : _GEN_3345; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3347 = 14'h35 == field_data_lo_25 ? _field_data_T_57 : _GEN_3346; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3348 = 14'h36 == field_data_lo_25 ? _field_data_T_58 : _GEN_3347; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3349 = 14'h37 == field_data_lo_25 ? _field_data_T_59 : _GEN_3348; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3350 = 14'h38 == field_data_lo_25 ? _field_data_T_60 : _GEN_3349; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3351 = 14'h39 == field_data_lo_25 ? _field_data_T_61 : _GEN_3350; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3352 = 14'h3a == field_data_lo_25 ? _field_data_T_62 : _GEN_3351; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3353 = 14'h3b == field_data_lo_25 ? _field_data_T_63 : _GEN_3352; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3354 = 14'h3c == field_data_lo_25 ? _field_data_T_64 : _GEN_3353; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3355 = 14'h3d == field_data_lo_25 ? _field_data_T_65 : _GEN_3354; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3356 = 14'h3e == field_data_lo_25 ? _field_data_T_66 : _GEN_3355; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3357 = 14'h3f == field_data_lo_25 ? _field_data_T_67 : _GEN_3356; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3358 = 14'h40 == field_data_lo_25 ? _field_data_T_68 : _GEN_3357; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3359 = 14'h41 == field_data_lo_25 ? _field_data_T_69 : _GEN_3358; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3360 = 14'h42 == field_data_lo_25 ? _field_data_T_70 : _GEN_3359; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3361 = 14'h43 == field_data_lo_25 ? _field_data_T_71 : _GEN_3360; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3362 = 14'h44 == field_data_lo_25 ? _field_data_T_72 : _GEN_3361; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3363 = 14'h45 == field_data_lo_25 ? _field_data_T_73 : _GEN_3362; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3364 = 14'h46 == field_data_lo_25 ? _field_data_T_74 : _GEN_3363; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3365 = 14'h47 == field_data_lo_25 ? _field_data_T_75 : _GEN_3364; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3366 = 14'h48 == field_data_lo_25 ? _field_data_T_76 : _GEN_3365; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3367 = 14'h49 == field_data_lo_25 ? _field_data_T_77 : _GEN_3366; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3368 = 14'h4a == field_data_lo_25 ? _field_data_T_78 : _GEN_3367; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3369 = 14'h4b == field_data_lo_25 ? _field_data_T_79 : _GEN_3368; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3370 = 14'h4c == field_data_lo_25 ? _field_data_T_80 : _GEN_3369; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3371 = 14'h4d == field_data_lo_25 ? _field_data_T_81 : _GEN_3370; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3372 = 14'h4e == field_data_lo_25 ? _field_data_T_82 : _GEN_3371; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3373 = 14'h4f == field_data_lo_25 ? _field_data_T_83 : _GEN_3372; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_58 = vliw_58[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_26 = vliw_58[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_58 = field_data_lo_26[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_58 = field_data_lo_26[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_84 = {{1'd0}, args_offset_58}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_84 = _total_offset_T_84[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3377 = 3'h1 == total_offset_84 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3378 = 3'h2 == total_offset_84 ? args_2 : _GEN_3377; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3379 = 3'h3 == total_offset_84 ? args_3 : _GEN_3378; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3380 = 3'h4 == total_offset_84 ? args_4 : _GEN_3379; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3381 = 3'h5 == total_offset_84 ? args_5 : _GEN_3380; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3382 = 3'h6 == total_offset_84 ? args_6 : _GEN_3381; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3383 = total_offset_84 < 3'h7 ? _GEN_3382 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_58_1 = 3'h0 < args_length_58 ? _GEN_3383 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_85 = args_offset_58 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3386 = 3'h1 == total_offset_85 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3387 = 3'h2 == total_offset_85 ? args_2 : _GEN_3386; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3388 = 3'h3 == total_offset_85 ? args_3 : _GEN_3387; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3389 = 3'h4 == total_offset_85 ? args_4 : _GEN_3388; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3390 = 3'h5 == total_offset_85 ? args_5 : _GEN_3389; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3391 = 3'h6 == total_offset_85 ? args_6 : _GEN_3390; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3392 = total_offset_85 < 3'h7 ? _GEN_3391 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_58_0 = 3'h1 < args_length_58 ? _GEN_3392 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1384 = {field_bytes_58_0,field_bytes_58_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_3394 = opcode_58 == 4'ha ? _field_data_T_1384 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3395 = opcode_58 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2735 = opcode_58 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_26 = field_data_lo_26[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1387 = {field_data_hi_26,field_data_lo_26}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_117 = _T_2735 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_3396 = opcode_58 == 4'h8 | opcode_58 == 4'hb ? _field_data_T_1387 : _GEN_3394; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3397 = opcode_58 == 4'h8 | opcode_58 == 4'hb ? _field_tag_T_117 : _GEN_3395; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_3398 = 14'h20 == field_data_lo_26 ? _field_data_T_36 : _GEN_3396; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3399 = 14'h21 == field_data_lo_26 ? _field_data_T_37 : _GEN_3398; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3400 = 14'h22 == field_data_lo_26 ? _field_data_T_38 : _GEN_3399; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3401 = 14'h23 == field_data_lo_26 ? _field_data_T_39 : _GEN_3400; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3402 = 14'h24 == field_data_lo_26 ? _field_data_T_40 : _GEN_3401; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3403 = 14'h25 == field_data_lo_26 ? _field_data_T_41 : _GEN_3402; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3404 = 14'h26 == field_data_lo_26 ? _field_data_T_42 : _GEN_3403; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3405 = 14'h27 == field_data_lo_26 ? _field_data_T_43 : _GEN_3404; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3406 = 14'h28 == field_data_lo_26 ? _field_data_T_44 : _GEN_3405; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3407 = 14'h29 == field_data_lo_26 ? _field_data_T_45 : _GEN_3406; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3408 = 14'h2a == field_data_lo_26 ? _field_data_T_46 : _GEN_3407; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3409 = 14'h2b == field_data_lo_26 ? _field_data_T_47 : _GEN_3408; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3410 = 14'h2c == field_data_lo_26 ? _field_data_T_48 : _GEN_3409; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3411 = 14'h2d == field_data_lo_26 ? _field_data_T_49 : _GEN_3410; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3412 = 14'h2e == field_data_lo_26 ? _field_data_T_50 : _GEN_3411; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3413 = 14'h2f == field_data_lo_26 ? _field_data_T_51 : _GEN_3412; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3414 = 14'h30 == field_data_lo_26 ? _field_data_T_52 : _GEN_3413; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3415 = 14'h31 == field_data_lo_26 ? _field_data_T_53 : _GEN_3414; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3416 = 14'h32 == field_data_lo_26 ? _field_data_T_54 : _GEN_3415; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3417 = 14'h33 == field_data_lo_26 ? _field_data_T_55 : _GEN_3416; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3418 = 14'h34 == field_data_lo_26 ? _field_data_T_56 : _GEN_3417; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3419 = 14'h35 == field_data_lo_26 ? _field_data_T_57 : _GEN_3418; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3420 = 14'h36 == field_data_lo_26 ? _field_data_T_58 : _GEN_3419; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3421 = 14'h37 == field_data_lo_26 ? _field_data_T_59 : _GEN_3420; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3422 = 14'h38 == field_data_lo_26 ? _field_data_T_60 : _GEN_3421; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3423 = 14'h39 == field_data_lo_26 ? _field_data_T_61 : _GEN_3422; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3424 = 14'h3a == field_data_lo_26 ? _field_data_T_62 : _GEN_3423; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3425 = 14'h3b == field_data_lo_26 ? _field_data_T_63 : _GEN_3424; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3426 = 14'h3c == field_data_lo_26 ? _field_data_T_64 : _GEN_3425; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3427 = 14'h3d == field_data_lo_26 ? _field_data_T_65 : _GEN_3426; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3428 = 14'h3e == field_data_lo_26 ? _field_data_T_66 : _GEN_3427; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3429 = 14'h3f == field_data_lo_26 ? _field_data_T_67 : _GEN_3428; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3430 = 14'h40 == field_data_lo_26 ? _field_data_T_68 : _GEN_3429; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3431 = 14'h41 == field_data_lo_26 ? _field_data_T_69 : _GEN_3430; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3432 = 14'h42 == field_data_lo_26 ? _field_data_T_70 : _GEN_3431; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3433 = 14'h43 == field_data_lo_26 ? _field_data_T_71 : _GEN_3432; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3434 = 14'h44 == field_data_lo_26 ? _field_data_T_72 : _GEN_3433; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3435 = 14'h45 == field_data_lo_26 ? _field_data_T_73 : _GEN_3434; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3436 = 14'h46 == field_data_lo_26 ? _field_data_T_74 : _GEN_3435; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3437 = 14'h47 == field_data_lo_26 ? _field_data_T_75 : _GEN_3436; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3438 = 14'h48 == field_data_lo_26 ? _field_data_T_76 : _GEN_3437; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3439 = 14'h49 == field_data_lo_26 ? _field_data_T_77 : _GEN_3438; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3440 = 14'h4a == field_data_lo_26 ? _field_data_T_78 : _GEN_3439; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3441 = 14'h4b == field_data_lo_26 ? _field_data_T_79 : _GEN_3440; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3442 = 14'h4c == field_data_lo_26 ? _field_data_T_80 : _GEN_3441; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3443 = 14'h4d == field_data_lo_26 ? _field_data_T_81 : _GEN_3442; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3444 = 14'h4e == field_data_lo_26 ? _field_data_T_82 : _GEN_3443; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3445 = 14'h4f == field_data_lo_26 ? _field_data_T_83 : _GEN_3444; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_59 = vliw_59[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_27 = vliw_59[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_59 = field_data_lo_27[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_59 = field_data_lo_27[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_86 = {{1'd0}, args_offset_59}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_86 = _total_offset_T_86[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3449 = 3'h1 == total_offset_86 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3450 = 3'h2 == total_offset_86 ? args_2 : _GEN_3449; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3451 = 3'h3 == total_offset_86 ? args_3 : _GEN_3450; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3452 = 3'h4 == total_offset_86 ? args_4 : _GEN_3451; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3453 = 3'h5 == total_offset_86 ? args_5 : _GEN_3452; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3454 = 3'h6 == total_offset_86 ? args_6 : _GEN_3453; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3455 = total_offset_86 < 3'h7 ? _GEN_3454 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_59_1 = 3'h0 < args_length_59 ? _GEN_3455 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_87 = args_offset_59 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3458 = 3'h1 == total_offset_87 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3459 = 3'h2 == total_offset_87 ? args_2 : _GEN_3458; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3460 = 3'h3 == total_offset_87 ? args_3 : _GEN_3459; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3461 = 3'h4 == total_offset_87 ? args_4 : _GEN_3460; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3462 = 3'h5 == total_offset_87 ? args_5 : _GEN_3461; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3463 = 3'h6 == total_offset_87 ? args_6 : _GEN_3462; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3464 = total_offset_87 < 3'h7 ? _GEN_3463 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_59_0 = 3'h1 < args_length_59 ? _GEN_3464 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1436 = {field_bytes_59_0,field_bytes_59_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_3466 = opcode_59 == 4'ha ? _field_data_T_1436 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3467 = opcode_59 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2792 = opcode_59 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_27 = field_data_lo_27[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1439 = {field_data_hi_27,field_data_lo_27}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_119 = _T_2792 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_3468 = opcode_59 == 4'h8 | opcode_59 == 4'hb ? _field_data_T_1439 : _GEN_3466; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3469 = opcode_59 == 4'h8 | opcode_59 == 4'hb ? _field_tag_T_119 : _GEN_3467; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_3470 = 14'h20 == field_data_lo_27 ? _field_data_T_36 : _GEN_3468; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3471 = 14'h21 == field_data_lo_27 ? _field_data_T_37 : _GEN_3470; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3472 = 14'h22 == field_data_lo_27 ? _field_data_T_38 : _GEN_3471; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3473 = 14'h23 == field_data_lo_27 ? _field_data_T_39 : _GEN_3472; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3474 = 14'h24 == field_data_lo_27 ? _field_data_T_40 : _GEN_3473; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3475 = 14'h25 == field_data_lo_27 ? _field_data_T_41 : _GEN_3474; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3476 = 14'h26 == field_data_lo_27 ? _field_data_T_42 : _GEN_3475; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3477 = 14'h27 == field_data_lo_27 ? _field_data_T_43 : _GEN_3476; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3478 = 14'h28 == field_data_lo_27 ? _field_data_T_44 : _GEN_3477; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3479 = 14'h29 == field_data_lo_27 ? _field_data_T_45 : _GEN_3478; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3480 = 14'h2a == field_data_lo_27 ? _field_data_T_46 : _GEN_3479; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3481 = 14'h2b == field_data_lo_27 ? _field_data_T_47 : _GEN_3480; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3482 = 14'h2c == field_data_lo_27 ? _field_data_T_48 : _GEN_3481; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3483 = 14'h2d == field_data_lo_27 ? _field_data_T_49 : _GEN_3482; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3484 = 14'h2e == field_data_lo_27 ? _field_data_T_50 : _GEN_3483; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3485 = 14'h2f == field_data_lo_27 ? _field_data_T_51 : _GEN_3484; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3486 = 14'h30 == field_data_lo_27 ? _field_data_T_52 : _GEN_3485; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3487 = 14'h31 == field_data_lo_27 ? _field_data_T_53 : _GEN_3486; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3488 = 14'h32 == field_data_lo_27 ? _field_data_T_54 : _GEN_3487; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3489 = 14'h33 == field_data_lo_27 ? _field_data_T_55 : _GEN_3488; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3490 = 14'h34 == field_data_lo_27 ? _field_data_T_56 : _GEN_3489; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3491 = 14'h35 == field_data_lo_27 ? _field_data_T_57 : _GEN_3490; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3492 = 14'h36 == field_data_lo_27 ? _field_data_T_58 : _GEN_3491; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3493 = 14'h37 == field_data_lo_27 ? _field_data_T_59 : _GEN_3492; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3494 = 14'h38 == field_data_lo_27 ? _field_data_T_60 : _GEN_3493; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3495 = 14'h39 == field_data_lo_27 ? _field_data_T_61 : _GEN_3494; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3496 = 14'h3a == field_data_lo_27 ? _field_data_T_62 : _GEN_3495; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3497 = 14'h3b == field_data_lo_27 ? _field_data_T_63 : _GEN_3496; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3498 = 14'h3c == field_data_lo_27 ? _field_data_T_64 : _GEN_3497; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3499 = 14'h3d == field_data_lo_27 ? _field_data_T_65 : _GEN_3498; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3500 = 14'h3e == field_data_lo_27 ? _field_data_T_66 : _GEN_3499; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3501 = 14'h3f == field_data_lo_27 ? _field_data_T_67 : _GEN_3500; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3502 = 14'h40 == field_data_lo_27 ? _field_data_T_68 : _GEN_3501; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3503 = 14'h41 == field_data_lo_27 ? _field_data_T_69 : _GEN_3502; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3504 = 14'h42 == field_data_lo_27 ? _field_data_T_70 : _GEN_3503; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3505 = 14'h43 == field_data_lo_27 ? _field_data_T_71 : _GEN_3504; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3506 = 14'h44 == field_data_lo_27 ? _field_data_T_72 : _GEN_3505; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3507 = 14'h45 == field_data_lo_27 ? _field_data_T_73 : _GEN_3506; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3508 = 14'h46 == field_data_lo_27 ? _field_data_T_74 : _GEN_3507; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3509 = 14'h47 == field_data_lo_27 ? _field_data_T_75 : _GEN_3508; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3510 = 14'h48 == field_data_lo_27 ? _field_data_T_76 : _GEN_3509; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3511 = 14'h49 == field_data_lo_27 ? _field_data_T_77 : _GEN_3510; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3512 = 14'h4a == field_data_lo_27 ? _field_data_T_78 : _GEN_3511; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3513 = 14'h4b == field_data_lo_27 ? _field_data_T_79 : _GEN_3512; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3514 = 14'h4c == field_data_lo_27 ? _field_data_T_80 : _GEN_3513; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3515 = 14'h4d == field_data_lo_27 ? _field_data_T_81 : _GEN_3514; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3516 = 14'h4e == field_data_lo_27 ? _field_data_T_82 : _GEN_3515; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3517 = 14'h4f == field_data_lo_27 ? _field_data_T_83 : _GEN_3516; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_60 = vliw_60[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_28 = vliw_60[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_60 = field_data_lo_28[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_60 = field_data_lo_28[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_88 = {{1'd0}, args_offset_60}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_88 = _total_offset_T_88[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3521 = 3'h1 == total_offset_88 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3522 = 3'h2 == total_offset_88 ? args_2 : _GEN_3521; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3523 = 3'h3 == total_offset_88 ? args_3 : _GEN_3522; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3524 = 3'h4 == total_offset_88 ? args_4 : _GEN_3523; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3525 = 3'h5 == total_offset_88 ? args_5 : _GEN_3524; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3526 = 3'h6 == total_offset_88 ? args_6 : _GEN_3525; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3527 = total_offset_88 < 3'h7 ? _GEN_3526 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_60_1 = 3'h0 < args_length_60 ? _GEN_3527 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_89 = args_offset_60 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3530 = 3'h1 == total_offset_89 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3531 = 3'h2 == total_offset_89 ? args_2 : _GEN_3530; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3532 = 3'h3 == total_offset_89 ? args_3 : _GEN_3531; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3533 = 3'h4 == total_offset_89 ? args_4 : _GEN_3532; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3534 = 3'h5 == total_offset_89 ? args_5 : _GEN_3533; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3535 = 3'h6 == total_offset_89 ? args_6 : _GEN_3534; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3536 = total_offset_89 < 3'h7 ? _GEN_3535 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_60_0 = 3'h1 < args_length_60 ? _GEN_3536 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1488 = {field_bytes_60_0,field_bytes_60_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_3538 = opcode_60 == 4'ha ? _field_data_T_1488 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3539 = opcode_60 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2849 = opcode_60 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_28 = field_data_lo_28[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1491 = {field_data_hi_28,field_data_lo_28}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_121 = _T_2849 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_3540 = opcode_60 == 4'h8 | opcode_60 == 4'hb ? _field_data_T_1491 : _GEN_3538; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3541 = opcode_60 == 4'h8 | opcode_60 == 4'hb ? _field_tag_T_121 : _GEN_3539; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_3542 = 14'h20 == field_data_lo_28 ? _field_data_T_36 : _GEN_3540; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3543 = 14'h21 == field_data_lo_28 ? _field_data_T_37 : _GEN_3542; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3544 = 14'h22 == field_data_lo_28 ? _field_data_T_38 : _GEN_3543; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3545 = 14'h23 == field_data_lo_28 ? _field_data_T_39 : _GEN_3544; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3546 = 14'h24 == field_data_lo_28 ? _field_data_T_40 : _GEN_3545; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3547 = 14'h25 == field_data_lo_28 ? _field_data_T_41 : _GEN_3546; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3548 = 14'h26 == field_data_lo_28 ? _field_data_T_42 : _GEN_3547; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3549 = 14'h27 == field_data_lo_28 ? _field_data_T_43 : _GEN_3548; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3550 = 14'h28 == field_data_lo_28 ? _field_data_T_44 : _GEN_3549; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3551 = 14'h29 == field_data_lo_28 ? _field_data_T_45 : _GEN_3550; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3552 = 14'h2a == field_data_lo_28 ? _field_data_T_46 : _GEN_3551; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3553 = 14'h2b == field_data_lo_28 ? _field_data_T_47 : _GEN_3552; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3554 = 14'h2c == field_data_lo_28 ? _field_data_T_48 : _GEN_3553; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3555 = 14'h2d == field_data_lo_28 ? _field_data_T_49 : _GEN_3554; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3556 = 14'h2e == field_data_lo_28 ? _field_data_T_50 : _GEN_3555; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3557 = 14'h2f == field_data_lo_28 ? _field_data_T_51 : _GEN_3556; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3558 = 14'h30 == field_data_lo_28 ? _field_data_T_52 : _GEN_3557; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3559 = 14'h31 == field_data_lo_28 ? _field_data_T_53 : _GEN_3558; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3560 = 14'h32 == field_data_lo_28 ? _field_data_T_54 : _GEN_3559; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3561 = 14'h33 == field_data_lo_28 ? _field_data_T_55 : _GEN_3560; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3562 = 14'h34 == field_data_lo_28 ? _field_data_T_56 : _GEN_3561; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3563 = 14'h35 == field_data_lo_28 ? _field_data_T_57 : _GEN_3562; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3564 = 14'h36 == field_data_lo_28 ? _field_data_T_58 : _GEN_3563; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3565 = 14'h37 == field_data_lo_28 ? _field_data_T_59 : _GEN_3564; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3566 = 14'h38 == field_data_lo_28 ? _field_data_T_60 : _GEN_3565; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3567 = 14'h39 == field_data_lo_28 ? _field_data_T_61 : _GEN_3566; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3568 = 14'h3a == field_data_lo_28 ? _field_data_T_62 : _GEN_3567; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3569 = 14'h3b == field_data_lo_28 ? _field_data_T_63 : _GEN_3568; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3570 = 14'h3c == field_data_lo_28 ? _field_data_T_64 : _GEN_3569; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3571 = 14'h3d == field_data_lo_28 ? _field_data_T_65 : _GEN_3570; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3572 = 14'h3e == field_data_lo_28 ? _field_data_T_66 : _GEN_3571; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3573 = 14'h3f == field_data_lo_28 ? _field_data_T_67 : _GEN_3572; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3574 = 14'h40 == field_data_lo_28 ? _field_data_T_68 : _GEN_3573; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3575 = 14'h41 == field_data_lo_28 ? _field_data_T_69 : _GEN_3574; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3576 = 14'h42 == field_data_lo_28 ? _field_data_T_70 : _GEN_3575; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3577 = 14'h43 == field_data_lo_28 ? _field_data_T_71 : _GEN_3576; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3578 = 14'h44 == field_data_lo_28 ? _field_data_T_72 : _GEN_3577; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3579 = 14'h45 == field_data_lo_28 ? _field_data_T_73 : _GEN_3578; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3580 = 14'h46 == field_data_lo_28 ? _field_data_T_74 : _GEN_3579; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3581 = 14'h47 == field_data_lo_28 ? _field_data_T_75 : _GEN_3580; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3582 = 14'h48 == field_data_lo_28 ? _field_data_T_76 : _GEN_3581; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3583 = 14'h49 == field_data_lo_28 ? _field_data_T_77 : _GEN_3582; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3584 = 14'h4a == field_data_lo_28 ? _field_data_T_78 : _GEN_3583; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3585 = 14'h4b == field_data_lo_28 ? _field_data_T_79 : _GEN_3584; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3586 = 14'h4c == field_data_lo_28 ? _field_data_T_80 : _GEN_3585; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3587 = 14'h4d == field_data_lo_28 ? _field_data_T_81 : _GEN_3586; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3588 = 14'h4e == field_data_lo_28 ? _field_data_T_82 : _GEN_3587; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3589 = 14'h4f == field_data_lo_28 ? _field_data_T_83 : _GEN_3588; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_61 = vliw_61[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_29 = vliw_61[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_61 = field_data_lo_29[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_61 = field_data_lo_29[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_90 = {{1'd0}, args_offset_61}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_90 = _total_offset_T_90[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3593 = 3'h1 == total_offset_90 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3594 = 3'h2 == total_offset_90 ? args_2 : _GEN_3593; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3595 = 3'h3 == total_offset_90 ? args_3 : _GEN_3594; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3596 = 3'h4 == total_offset_90 ? args_4 : _GEN_3595; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3597 = 3'h5 == total_offset_90 ? args_5 : _GEN_3596; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3598 = 3'h6 == total_offset_90 ? args_6 : _GEN_3597; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3599 = total_offset_90 < 3'h7 ? _GEN_3598 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_61_1 = 3'h0 < args_length_61 ? _GEN_3599 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_91 = args_offset_61 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3602 = 3'h1 == total_offset_91 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3603 = 3'h2 == total_offset_91 ? args_2 : _GEN_3602; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3604 = 3'h3 == total_offset_91 ? args_3 : _GEN_3603; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3605 = 3'h4 == total_offset_91 ? args_4 : _GEN_3604; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3606 = 3'h5 == total_offset_91 ? args_5 : _GEN_3605; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3607 = 3'h6 == total_offset_91 ? args_6 : _GEN_3606; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3608 = total_offset_91 < 3'h7 ? _GEN_3607 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_61_0 = 3'h1 < args_length_61 ? _GEN_3608 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1540 = {field_bytes_61_0,field_bytes_61_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_3610 = opcode_61 == 4'ha ? _field_data_T_1540 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3611 = opcode_61 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2906 = opcode_61 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_29 = field_data_lo_29[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1543 = {field_data_hi_29,field_data_lo_29}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_123 = _T_2906 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_3612 = opcode_61 == 4'h8 | opcode_61 == 4'hb ? _field_data_T_1543 : _GEN_3610; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3613 = opcode_61 == 4'h8 | opcode_61 == 4'hb ? _field_tag_T_123 : _GEN_3611; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_3614 = 14'h20 == field_data_lo_29 ? _field_data_T_36 : _GEN_3612; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3615 = 14'h21 == field_data_lo_29 ? _field_data_T_37 : _GEN_3614; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3616 = 14'h22 == field_data_lo_29 ? _field_data_T_38 : _GEN_3615; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3617 = 14'h23 == field_data_lo_29 ? _field_data_T_39 : _GEN_3616; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3618 = 14'h24 == field_data_lo_29 ? _field_data_T_40 : _GEN_3617; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3619 = 14'h25 == field_data_lo_29 ? _field_data_T_41 : _GEN_3618; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3620 = 14'h26 == field_data_lo_29 ? _field_data_T_42 : _GEN_3619; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3621 = 14'h27 == field_data_lo_29 ? _field_data_T_43 : _GEN_3620; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3622 = 14'h28 == field_data_lo_29 ? _field_data_T_44 : _GEN_3621; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3623 = 14'h29 == field_data_lo_29 ? _field_data_T_45 : _GEN_3622; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3624 = 14'h2a == field_data_lo_29 ? _field_data_T_46 : _GEN_3623; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3625 = 14'h2b == field_data_lo_29 ? _field_data_T_47 : _GEN_3624; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3626 = 14'h2c == field_data_lo_29 ? _field_data_T_48 : _GEN_3625; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3627 = 14'h2d == field_data_lo_29 ? _field_data_T_49 : _GEN_3626; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3628 = 14'h2e == field_data_lo_29 ? _field_data_T_50 : _GEN_3627; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3629 = 14'h2f == field_data_lo_29 ? _field_data_T_51 : _GEN_3628; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3630 = 14'h30 == field_data_lo_29 ? _field_data_T_52 : _GEN_3629; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3631 = 14'h31 == field_data_lo_29 ? _field_data_T_53 : _GEN_3630; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3632 = 14'h32 == field_data_lo_29 ? _field_data_T_54 : _GEN_3631; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3633 = 14'h33 == field_data_lo_29 ? _field_data_T_55 : _GEN_3632; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3634 = 14'h34 == field_data_lo_29 ? _field_data_T_56 : _GEN_3633; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3635 = 14'h35 == field_data_lo_29 ? _field_data_T_57 : _GEN_3634; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3636 = 14'h36 == field_data_lo_29 ? _field_data_T_58 : _GEN_3635; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3637 = 14'h37 == field_data_lo_29 ? _field_data_T_59 : _GEN_3636; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3638 = 14'h38 == field_data_lo_29 ? _field_data_T_60 : _GEN_3637; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3639 = 14'h39 == field_data_lo_29 ? _field_data_T_61 : _GEN_3638; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3640 = 14'h3a == field_data_lo_29 ? _field_data_T_62 : _GEN_3639; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3641 = 14'h3b == field_data_lo_29 ? _field_data_T_63 : _GEN_3640; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3642 = 14'h3c == field_data_lo_29 ? _field_data_T_64 : _GEN_3641; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3643 = 14'h3d == field_data_lo_29 ? _field_data_T_65 : _GEN_3642; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3644 = 14'h3e == field_data_lo_29 ? _field_data_T_66 : _GEN_3643; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3645 = 14'h3f == field_data_lo_29 ? _field_data_T_67 : _GEN_3644; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3646 = 14'h40 == field_data_lo_29 ? _field_data_T_68 : _GEN_3645; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3647 = 14'h41 == field_data_lo_29 ? _field_data_T_69 : _GEN_3646; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3648 = 14'h42 == field_data_lo_29 ? _field_data_T_70 : _GEN_3647; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3649 = 14'h43 == field_data_lo_29 ? _field_data_T_71 : _GEN_3648; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3650 = 14'h44 == field_data_lo_29 ? _field_data_T_72 : _GEN_3649; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3651 = 14'h45 == field_data_lo_29 ? _field_data_T_73 : _GEN_3650; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3652 = 14'h46 == field_data_lo_29 ? _field_data_T_74 : _GEN_3651; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3653 = 14'h47 == field_data_lo_29 ? _field_data_T_75 : _GEN_3652; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3654 = 14'h48 == field_data_lo_29 ? _field_data_T_76 : _GEN_3653; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3655 = 14'h49 == field_data_lo_29 ? _field_data_T_77 : _GEN_3654; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3656 = 14'h4a == field_data_lo_29 ? _field_data_T_78 : _GEN_3655; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3657 = 14'h4b == field_data_lo_29 ? _field_data_T_79 : _GEN_3656; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3658 = 14'h4c == field_data_lo_29 ? _field_data_T_80 : _GEN_3657; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3659 = 14'h4d == field_data_lo_29 ? _field_data_T_81 : _GEN_3658; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3660 = 14'h4e == field_data_lo_29 ? _field_data_T_82 : _GEN_3659; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3661 = 14'h4f == field_data_lo_29 ? _field_data_T_83 : _GEN_3660; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_62 = vliw_62[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_30 = vliw_62[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_62 = field_data_lo_30[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_62 = field_data_lo_30[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_92 = {{1'd0}, args_offset_62}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_92 = _total_offset_T_92[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3665 = 3'h1 == total_offset_92 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3666 = 3'h2 == total_offset_92 ? args_2 : _GEN_3665; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3667 = 3'h3 == total_offset_92 ? args_3 : _GEN_3666; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3668 = 3'h4 == total_offset_92 ? args_4 : _GEN_3667; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3669 = 3'h5 == total_offset_92 ? args_5 : _GEN_3668; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3670 = 3'h6 == total_offset_92 ? args_6 : _GEN_3669; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3671 = total_offset_92 < 3'h7 ? _GEN_3670 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_62_1 = 3'h0 < args_length_62 ? _GEN_3671 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_93 = args_offset_62 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3674 = 3'h1 == total_offset_93 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3675 = 3'h2 == total_offset_93 ? args_2 : _GEN_3674; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3676 = 3'h3 == total_offset_93 ? args_3 : _GEN_3675; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3677 = 3'h4 == total_offset_93 ? args_4 : _GEN_3676; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3678 = 3'h5 == total_offset_93 ? args_5 : _GEN_3677; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3679 = 3'h6 == total_offset_93 ? args_6 : _GEN_3678; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3680 = total_offset_93 < 3'h7 ? _GEN_3679 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_62_0 = 3'h1 < args_length_62 ? _GEN_3680 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1592 = {field_bytes_62_0,field_bytes_62_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_3682 = opcode_62 == 4'ha ? _field_data_T_1592 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3683 = opcode_62 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2963 = opcode_62 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_30 = field_data_lo_30[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1595 = {field_data_hi_30,field_data_lo_30}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_125 = _T_2963 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_3684 = opcode_62 == 4'h8 | opcode_62 == 4'hb ? _field_data_T_1595 : _GEN_3682; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3685 = opcode_62 == 4'h8 | opcode_62 == 4'hb ? _field_tag_T_125 : _GEN_3683; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_3686 = 14'h20 == field_data_lo_30 ? _field_data_T_36 : _GEN_3684; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3687 = 14'h21 == field_data_lo_30 ? _field_data_T_37 : _GEN_3686; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3688 = 14'h22 == field_data_lo_30 ? _field_data_T_38 : _GEN_3687; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3689 = 14'h23 == field_data_lo_30 ? _field_data_T_39 : _GEN_3688; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3690 = 14'h24 == field_data_lo_30 ? _field_data_T_40 : _GEN_3689; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3691 = 14'h25 == field_data_lo_30 ? _field_data_T_41 : _GEN_3690; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3692 = 14'h26 == field_data_lo_30 ? _field_data_T_42 : _GEN_3691; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3693 = 14'h27 == field_data_lo_30 ? _field_data_T_43 : _GEN_3692; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3694 = 14'h28 == field_data_lo_30 ? _field_data_T_44 : _GEN_3693; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3695 = 14'h29 == field_data_lo_30 ? _field_data_T_45 : _GEN_3694; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3696 = 14'h2a == field_data_lo_30 ? _field_data_T_46 : _GEN_3695; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3697 = 14'h2b == field_data_lo_30 ? _field_data_T_47 : _GEN_3696; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3698 = 14'h2c == field_data_lo_30 ? _field_data_T_48 : _GEN_3697; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3699 = 14'h2d == field_data_lo_30 ? _field_data_T_49 : _GEN_3698; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3700 = 14'h2e == field_data_lo_30 ? _field_data_T_50 : _GEN_3699; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3701 = 14'h2f == field_data_lo_30 ? _field_data_T_51 : _GEN_3700; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3702 = 14'h30 == field_data_lo_30 ? _field_data_T_52 : _GEN_3701; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3703 = 14'h31 == field_data_lo_30 ? _field_data_T_53 : _GEN_3702; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3704 = 14'h32 == field_data_lo_30 ? _field_data_T_54 : _GEN_3703; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3705 = 14'h33 == field_data_lo_30 ? _field_data_T_55 : _GEN_3704; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3706 = 14'h34 == field_data_lo_30 ? _field_data_T_56 : _GEN_3705; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3707 = 14'h35 == field_data_lo_30 ? _field_data_T_57 : _GEN_3706; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3708 = 14'h36 == field_data_lo_30 ? _field_data_T_58 : _GEN_3707; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3709 = 14'h37 == field_data_lo_30 ? _field_data_T_59 : _GEN_3708; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3710 = 14'h38 == field_data_lo_30 ? _field_data_T_60 : _GEN_3709; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3711 = 14'h39 == field_data_lo_30 ? _field_data_T_61 : _GEN_3710; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3712 = 14'h3a == field_data_lo_30 ? _field_data_T_62 : _GEN_3711; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3713 = 14'h3b == field_data_lo_30 ? _field_data_T_63 : _GEN_3712; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3714 = 14'h3c == field_data_lo_30 ? _field_data_T_64 : _GEN_3713; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3715 = 14'h3d == field_data_lo_30 ? _field_data_T_65 : _GEN_3714; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3716 = 14'h3e == field_data_lo_30 ? _field_data_T_66 : _GEN_3715; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3717 = 14'h3f == field_data_lo_30 ? _field_data_T_67 : _GEN_3716; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3718 = 14'h40 == field_data_lo_30 ? _field_data_T_68 : _GEN_3717; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3719 = 14'h41 == field_data_lo_30 ? _field_data_T_69 : _GEN_3718; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3720 = 14'h42 == field_data_lo_30 ? _field_data_T_70 : _GEN_3719; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3721 = 14'h43 == field_data_lo_30 ? _field_data_T_71 : _GEN_3720; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3722 = 14'h44 == field_data_lo_30 ? _field_data_T_72 : _GEN_3721; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3723 = 14'h45 == field_data_lo_30 ? _field_data_T_73 : _GEN_3722; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3724 = 14'h46 == field_data_lo_30 ? _field_data_T_74 : _GEN_3723; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3725 = 14'h47 == field_data_lo_30 ? _field_data_T_75 : _GEN_3724; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3726 = 14'h48 == field_data_lo_30 ? _field_data_T_76 : _GEN_3725; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3727 = 14'h49 == field_data_lo_30 ? _field_data_T_77 : _GEN_3726; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3728 = 14'h4a == field_data_lo_30 ? _field_data_T_78 : _GEN_3727; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3729 = 14'h4b == field_data_lo_30 ? _field_data_T_79 : _GEN_3728; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3730 = 14'h4c == field_data_lo_30 ? _field_data_T_80 : _GEN_3729; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3731 = 14'h4d == field_data_lo_30 ? _field_data_T_81 : _GEN_3730; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3732 = 14'h4e == field_data_lo_30 ? _field_data_T_82 : _GEN_3731; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3733 = 14'h4f == field_data_lo_30 ? _field_data_T_83 : _GEN_3732; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_63 = vliw_63[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_31 = vliw_63[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_63 = field_data_lo_31[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_63 = field_data_lo_31[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_94 = {{1'd0}, args_offset_63}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_94 = _total_offset_T_94[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3737 = 3'h1 == total_offset_94 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3738 = 3'h2 == total_offset_94 ? args_2 : _GEN_3737; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3739 = 3'h3 == total_offset_94 ? args_3 : _GEN_3738; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3740 = 3'h4 == total_offset_94 ? args_4 : _GEN_3739; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3741 = 3'h5 == total_offset_94 ? args_5 : _GEN_3740; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3742 = 3'h6 == total_offset_94 ? args_6 : _GEN_3741; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3743 = total_offset_94 < 3'h7 ? _GEN_3742 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_63_1 = 3'h0 < args_length_63 ? _GEN_3743 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_95 = args_offset_63 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3746 = 3'h1 == total_offset_95 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3747 = 3'h2 == total_offset_95 ? args_2 : _GEN_3746; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3748 = 3'h3 == total_offset_95 ? args_3 : _GEN_3747; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3749 = 3'h4 == total_offset_95 ? args_4 : _GEN_3748; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3750 = 3'h5 == total_offset_95 ? args_5 : _GEN_3749; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3751 = 3'h6 == total_offset_95 ? args_6 : _GEN_3750; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3752 = total_offset_95 < 3'h7 ? _GEN_3751 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_63_0 = 3'h1 < args_length_63 ? _GEN_3752 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1644 = {field_bytes_63_0,field_bytes_63_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_3754 = opcode_63 == 4'ha ? _field_data_T_1644 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3755 = opcode_63 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3020 = opcode_63 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_31 = field_data_lo_31[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1647 = {field_data_hi_31,field_data_lo_31}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_127 = _T_3020 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_3756 = opcode_63 == 4'h8 | opcode_63 == 4'hb ? _field_data_T_1647 : _GEN_3754; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3757 = opcode_63 == 4'h8 | opcode_63 == 4'hb ? _field_tag_T_127 : _GEN_3755; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_3758 = 14'h20 == field_data_lo_31 ? _field_data_T_36 : _GEN_3756; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3759 = 14'h21 == field_data_lo_31 ? _field_data_T_37 : _GEN_3758; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3760 = 14'h22 == field_data_lo_31 ? _field_data_T_38 : _GEN_3759; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3761 = 14'h23 == field_data_lo_31 ? _field_data_T_39 : _GEN_3760; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3762 = 14'h24 == field_data_lo_31 ? _field_data_T_40 : _GEN_3761; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3763 = 14'h25 == field_data_lo_31 ? _field_data_T_41 : _GEN_3762; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3764 = 14'h26 == field_data_lo_31 ? _field_data_T_42 : _GEN_3763; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3765 = 14'h27 == field_data_lo_31 ? _field_data_T_43 : _GEN_3764; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3766 = 14'h28 == field_data_lo_31 ? _field_data_T_44 : _GEN_3765; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3767 = 14'h29 == field_data_lo_31 ? _field_data_T_45 : _GEN_3766; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3768 = 14'h2a == field_data_lo_31 ? _field_data_T_46 : _GEN_3767; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3769 = 14'h2b == field_data_lo_31 ? _field_data_T_47 : _GEN_3768; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3770 = 14'h2c == field_data_lo_31 ? _field_data_T_48 : _GEN_3769; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3771 = 14'h2d == field_data_lo_31 ? _field_data_T_49 : _GEN_3770; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3772 = 14'h2e == field_data_lo_31 ? _field_data_T_50 : _GEN_3771; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3773 = 14'h2f == field_data_lo_31 ? _field_data_T_51 : _GEN_3772; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3774 = 14'h30 == field_data_lo_31 ? _field_data_T_52 : _GEN_3773; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3775 = 14'h31 == field_data_lo_31 ? _field_data_T_53 : _GEN_3774; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3776 = 14'h32 == field_data_lo_31 ? _field_data_T_54 : _GEN_3775; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3777 = 14'h33 == field_data_lo_31 ? _field_data_T_55 : _GEN_3776; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3778 = 14'h34 == field_data_lo_31 ? _field_data_T_56 : _GEN_3777; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3779 = 14'h35 == field_data_lo_31 ? _field_data_T_57 : _GEN_3778; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3780 = 14'h36 == field_data_lo_31 ? _field_data_T_58 : _GEN_3779; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3781 = 14'h37 == field_data_lo_31 ? _field_data_T_59 : _GEN_3780; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3782 = 14'h38 == field_data_lo_31 ? _field_data_T_60 : _GEN_3781; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3783 = 14'h39 == field_data_lo_31 ? _field_data_T_61 : _GEN_3782; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3784 = 14'h3a == field_data_lo_31 ? _field_data_T_62 : _GEN_3783; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3785 = 14'h3b == field_data_lo_31 ? _field_data_T_63 : _GEN_3784; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3786 = 14'h3c == field_data_lo_31 ? _field_data_T_64 : _GEN_3785; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3787 = 14'h3d == field_data_lo_31 ? _field_data_T_65 : _GEN_3786; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3788 = 14'h3e == field_data_lo_31 ? _field_data_T_66 : _GEN_3787; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3789 = 14'h3f == field_data_lo_31 ? _field_data_T_67 : _GEN_3788; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3790 = 14'h40 == field_data_lo_31 ? _field_data_T_68 : _GEN_3789; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3791 = 14'h41 == field_data_lo_31 ? _field_data_T_69 : _GEN_3790; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3792 = 14'h42 == field_data_lo_31 ? _field_data_T_70 : _GEN_3791; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3793 = 14'h43 == field_data_lo_31 ? _field_data_T_71 : _GEN_3792; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3794 = 14'h44 == field_data_lo_31 ? _field_data_T_72 : _GEN_3793; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3795 = 14'h45 == field_data_lo_31 ? _field_data_T_73 : _GEN_3794; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3796 = 14'h46 == field_data_lo_31 ? _field_data_T_74 : _GEN_3795; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3797 = 14'h47 == field_data_lo_31 ? _field_data_T_75 : _GEN_3796; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3798 = 14'h48 == field_data_lo_31 ? _field_data_T_76 : _GEN_3797; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3799 = 14'h49 == field_data_lo_31 ? _field_data_T_77 : _GEN_3798; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3800 = 14'h4a == field_data_lo_31 ? _field_data_T_78 : _GEN_3799; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3801 = 14'h4b == field_data_lo_31 ? _field_data_T_79 : _GEN_3800; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3802 = 14'h4c == field_data_lo_31 ? _field_data_T_80 : _GEN_3801; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3803 = 14'h4d == field_data_lo_31 ? _field_data_T_81 : _GEN_3802; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3804 = 14'h4e == field_data_lo_31 ? _field_data_T_82 : _GEN_3803; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3805 = 14'h4f == field_data_lo_31 ? _field_data_T_83 : _GEN_3804; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_64 = vliw_64[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_32 = vliw_64[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_64 = field_data_lo_32[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_64 = field_data_lo_32[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_96 = {{1'd0}, args_offset_64}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_96 = _total_offset_T_96[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3809 = 3'h1 == total_offset_96 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3810 = 3'h2 == total_offset_96 ? args_2 : _GEN_3809; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3811 = 3'h3 == total_offset_96 ? args_3 : _GEN_3810; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3812 = 3'h4 == total_offset_96 ? args_4 : _GEN_3811; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3813 = 3'h5 == total_offset_96 ? args_5 : _GEN_3812; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3814 = 3'h6 == total_offset_96 ? args_6 : _GEN_3813; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3815 = total_offset_96 < 3'h7 ? _GEN_3814 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_64_1 = 3'h0 < args_length_64 ? _GEN_3815 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_97 = args_offset_64 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3818 = 3'h1 == total_offset_97 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3819 = 3'h2 == total_offset_97 ? args_2 : _GEN_3818; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3820 = 3'h3 == total_offset_97 ? args_3 : _GEN_3819; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3821 = 3'h4 == total_offset_97 ? args_4 : _GEN_3820; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3822 = 3'h5 == total_offset_97 ? args_5 : _GEN_3821; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3823 = 3'h6 == total_offset_97 ? args_6 : _GEN_3822; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3824 = total_offset_97 < 3'h7 ? _GEN_3823 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_64_0 = 3'h1 < args_length_64 ? _GEN_3824 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1696 = {field_bytes_64_0,field_bytes_64_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_3826 = opcode_64 == 4'ha ? _field_data_T_1696 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3827 = opcode_64 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3077 = opcode_64 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_32 = field_data_lo_32[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1699 = {field_data_hi_32,field_data_lo_32}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_129 = _T_3077 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_3828 = opcode_64 == 4'h8 | opcode_64 == 4'hb ? _field_data_T_1699 : _GEN_3826; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3829 = opcode_64 == 4'h8 | opcode_64 == 4'hb ? _field_tag_T_129 : _GEN_3827; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_3830 = 14'h20 == field_data_lo_32 ? _field_data_T_36 : _GEN_3828; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3831 = 14'h21 == field_data_lo_32 ? _field_data_T_37 : _GEN_3830; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3832 = 14'h22 == field_data_lo_32 ? _field_data_T_38 : _GEN_3831; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3833 = 14'h23 == field_data_lo_32 ? _field_data_T_39 : _GEN_3832; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3834 = 14'h24 == field_data_lo_32 ? _field_data_T_40 : _GEN_3833; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3835 = 14'h25 == field_data_lo_32 ? _field_data_T_41 : _GEN_3834; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3836 = 14'h26 == field_data_lo_32 ? _field_data_T_42 : _GEN_3835; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3837 = 14'h27 == field_data_lo_32 ? _field_data_T_43 : _GEN_3836; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3838 = 14'h28 == field_data_lo_32 ? _field_data_T_44 : _GEN_3837; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3839 = 14'h29 == field_data_lo_32 ? _field_data_T_45 : _GEN_3838; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3840 = 14'h2a == field_data_lo_32 ? _field_data_T_46 : _GEN_3839; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3841 = 14'h2b == field_data_lo_32 ? _field_data_T_47 : _GEN_3840; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3842 = 14'h2c == field_data_lo_32 ? _field_data_T_48 : _GEN_3841; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3843 = 14'h2d == field_data_lo_32 ? _field_data_T_49 : _GEN_3842; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3844 = 14'h2e == field_data_lo_32 ? _field_data_T_50 : _GEN_3843; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3845 = 14'h2f == field_data_lo_32 ? _field_data_T_51 : _GEN_3844; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3846 = 14'h30 == field_data_lo_32 ? _field_data_T_52 : _GEN_3845; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3847 = 14'h31 == field_data_lo_32 ? _field_data_T_53 : _GEN_3846; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3848 = 14'h32 == field_data_lo_32 ? _field_data_T_54 : _GEN_3847; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3849 = 14'h33 == field_data_lo_32 ? _field_data_T_55 : _GEN_3848; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3850 = 14'h34 == field_data_lo_32 ? _field_data_T_56 : _GEN_3849; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3851 = 14'h35 == field_data_lo_32 ? _field_data_T_57 : _GEN_3850; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3852 = 14'h36 == field_data_lo_32 ? _field_data_T_58 : _GEN_3851; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3853 = 14'h37 == field_data_lo_32 ? _field_data_T_59 : _GEN_3852; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3854 = 14'h38 == field_data_lo_32 ? _field_data_T_60 : _GEN_3853; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3855 = 14'h39 == field_data_lo_32 ? _field_data_T_61 : _GEN_3854; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3856 = 14'h3a == field_data_lo_32 ? _field_data_T_62 : _GEN_3855; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3857 = 14'h3b == field_data_lo_32 ? _field_data_T_63 : _GEN_3856; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3858 = 14'h3c == field_data_lo_32 ? _field_data_T_64 : _GEN_3857; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3859 = 14'h3d == field_data_lo_32 ? _field_data_T_65 : _GEN_3858; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3860 = 14'h3e == field_data_lo_32 ? _field_data_T_66 : _GEN_3859; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3861 = 14'h3f == field_data_lo_32 ? _field_data_T_67 : _GEN_3860; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3862 = 14'h40 == field_data_lo_32 ? _field_data_T_68 : _GEN_3861; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3863 = 14'h41 == field_data_lo_32 ? _field_data_T_69 : _GEN_3862; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3864 = 14'h42 == field_data_lo_32 ? _field_data_T_70 : _GEN_3863; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3865 = 14'h43 == field_data_lo_32 ? _field_data_T_71 : _GEN_3864; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3866 = 14'h44 == field_data_lo_32 ? _field_data_T_72 : _GEN_3865; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3867 = 14'h45 == field_data_lo_32 ? _field_data_T_73 : _GEN_3866; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3868 = 14'h46 == field_data_lo_32 ? _field_data_T_74 : _GEN_3867; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3869 = 14'h47 == field_data_lo_32 ? _field_data_T_75 : _GEN_3868; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3870 = 14'h48 == field_data_lo_32 ? _field_data_T_76 : _GEN_3869; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3871 = 14'h49 == field_data_lo_32 ? _field_data_T_77 : _GEN_3870; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3872 = 14'h4a == field_data_lo_32 ? _field_data_T_78 : _GEN_3871; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3873 = 14'h4b == field_data_lo_32 ? _field_data_T_79 : _GEN_3872; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3874 = 14'h4c == field_data_lo_32 ? _field_data_T_80 : _GEN_3873; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3875 = 14'h4d == field_data_lo_32 ? _field_data_T_81 : _GEN_3874; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3876 = 14'h4e == field_data_lo_32 ? _field_data_T_82 : _GEN_3875; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3877 = 14'h4f == field_data_lo_32 ? _field_data_T_83 : _GEN_3876; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_65 = vliw_65[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_33 = vliw_65[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_65 = field_data_lo_33[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_65 = field_data_lo_33[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_98 = {{1'd0}, args_offset_65}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_98 = _total_offset_T_98[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3881 = 3'h1 == total_offset_98 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3882 = 3'h2 == total_offset_98 ? args_2 : _GEN_3881; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3883 = 3'h3 == total_offset_98 ? args_3 : _GEN_3882; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3884 = 3'h4 == total_offset_98 ? args_4 : _GEN_3883; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3885 = 3'h5 == total_offset_98 ? args_5 : _GEN_3884; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3886 = 3'h6 == total_offset_98 ? args_6 : _GEN_3885; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3887 = total_offset_98 < 3'h7 ? _GEN_3886 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_65_1 = 3'h0 < args_length_65 ? _GEN_3887 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_99 = args_offset_65 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3890 = 3'h1 == total_offset_99 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3891 = 3'h2 == total_offset_99 ? args_2 : _GEN_3890; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3892 = 3'h3 == total_offset_99 ? args_3 : _GEN_3891; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3893 = 3'h4 == total_offset_99 ? args_4 : _GEN_3892; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3894 = 3'h5 == total_offset_99 ? args_5 : _GEN_3893; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3895 = 3'h6 == total_offset_99 ? args_6 : _GEN_3894; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3896 = total_offset_99 < 3'h7 ? _GEN_3895 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_65_0 = 3'h1 < args_length_65 ? _GEN_3896 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1748 = {field_bytes_65_0,field_bytes_65_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_3898 = opcode_65 == 4'ha ? _field_data_T_1748 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3899 = opcode_65 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3134 = opcode_65 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_33 = field_data_lo_33[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1751 = {field_data_hi_33,field_data_lo_33}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_131 = _T_3134 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_3900 = opcode_65 == 4'h8 | opcode_65 == 4'hb ? _field_data_T_1751 : _GEN_3898; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3901 = opcode_65 == 4'h8 | opcode_65 == 4'hb ? _field_tag_T_131 : _GEN_3899; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_3902 = 14'h20 == field_data_lo_33 ? _field_data_T_36 : _GEN_3900; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3903 = 14'h21 == field_data_lo_33 ? _field_data_T_37 : _GEN_3902; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3904 = 14'h22 == field_data_lo_33 ? _field_data_T_38 : _GEN_3903; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3905 = 14'h23 == field_data_lo_33 ? _field_data_T_39 : _GEN_3904; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3906 = 14'h24 == field_data_lo_33 ? _field_data_T_40 : _GEN_3905; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3907 = 14'h25 == field_data_lo_33 ? _field_data_T_41 : _GEN_3906; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3908 = 14'h26 == field_data_lo_33 ? _field_data_T_42 : _GEN_3907; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3909 = 14'h27 == field_data_lo_33 ? _field_data_T_43 : _GEN_3908; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3910 = 14'h28 == field_data_lo_33 ? _field_data_T_44 : _GEN_3909; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3911 = 14'h29 == field_data_lo_33 ? _field_data_T_45 : _GEN_3910; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3912 = 14'h2a == field_data_lo_33 ? _field_data_T_46 : _GEN_3911; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3913 = 14'h2b == field_data_lo_33 ? _field_data_T_47 : _GEN_3912; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3914 = 14'h2c == field_data_lo_33 ? _field_data_T_48 : _GEN_3913; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3915 = 14'h2d == field_data_lo_33 ? _field_data_T_49 : _GEN_3914; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3916 = 14'h2e == field_data_lo_33 ? _field_data_T_50 : _GEN_3915; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3917 = 14'h2f == field_data_lo_33 ? _field_data_T_51 : _GEN_3916; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3918 = 14'h30 == field_data_lo_33 ? _field_data_T_52 : _GEN_3917; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3919 = 14'h31 == field_data_lo_33 ? _field_data_T_53 : _GEN_3918; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3920 = 14'h32 == field_data_lo_33 ? _field_data_T_54 : _GEN_3919; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3921 = 14'h33 == field_data_lo_33 ? _field_data_T_55 : _GEN_3920; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3922 = 14'h34 == field_data_lo_33 ? _field_data_T_56 : _GEN_3921; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3923 = 14'h35 == field_data_lo_33 ? _field_data_T_57 : _GEN_3922; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3924 = 14'h36 == field_data_lo_33 ? _field_data_T_58 : _GEN_3923; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3925 = 14'h37 == field_data_lo_33 ? _field_data_T_59 : _GEN_3924; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3926 = 14'h38 == field_data_lo_33 ? _field_data_T_60 : _GEN_3925; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3927 = 14'h39 == field_data_lo_33 ? _field_data_T_61 : _GEN_3926; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3928 = 14'h3a == field_data_lo_33 ? _field_data_T_62 : _GEN_3927; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3929 = 14'h3b == field_data_lo_33 ? _field_data_T_63 : _GEN_3928; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3930 = 14'h3c == field_data_lo_33 ? _field_data_T_64 : _GEN_3929; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3931 = 14'h3d == field_data_lo_33 ? _field_data_T_65 : _GEN_3930; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3932 = 14'h3e == field_data_lo_33 ? _field_data_T_66 : _GEN_3931; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3933 = 14'h3f == field_data_lo_33 ? _field_data_T_67 : _GEN_3932; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3934 = 14'h40 == field_data_lo_33 ? _field_data_T_68 : _GEN_3933; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3935 = 14'h41 == field_data_lo_33 ? _field_data_T_69 : _GEN_3934; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3936 = 14'h42 == field_data_lo_33 ? _field_data_T_70 : _GEN_3935; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3937 = 14'h43 == field_data_lo_33 ? _field_data_T_71 : _GEN_3936; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3938 = 14'h44 == field_data_lo_33 ? _field_data_T_72 : _GEN_3937; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3939 = 14'h45 == field_data_lo_33 ? _field_data_T_73 : _GEN_3938; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3940 = 14'h46 == field_data_lo_33 ? _field_data_T_74 : _GEN_3939; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3941 = 14'h47 == field_data_lo_33 ? _field_data_T_75 : _GEN_3940; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3942 = 14'h48 == field_data_lo_33 ? _field_data_T_76 : _GEN_3941; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3943 = 14'h49 == field_data_lo_33 ? _field_data_T_77 : _GEN_3942; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3944 = 14'h4a == field_data_lo_33 ? _field_data_T_78 : _GEN_3943; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3945 = 14'h4b == field_data_lo_33 ? _field_data_T_79 : _GEN_3944; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3946 = 14'h4c == field_data_lo_33 ? _field_data_T_80 : _GEN_3945; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3947 = 14'h4d == field_data_lo_33 ? _field_data_T_81 : _GEN_3946; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3948 = 14'h4e == field_data_lo_33 ? _field_data_T_82 : _GEN_3947; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3949 = 14'h4f == field_data_lo_33 ? _field_data_T_83 : _GEN_3948; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_66 = vliw_66[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_34 = vliw_66[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_66 = field_data_lo_34[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_66 = field_data_lo_34[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_100 = {{1'd0}, args_offset_66}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_100 = _total_offset_T_100[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3953 = 3'h1 == total_offset_100 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3954 = 3'h2 == total_offset_100 ? args_2 : _GEN_3953; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3955 = 3'h3 == total_offset_100 ? args_3 : _GEN_3954; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3956 = 3'h4 == total_offset_100 ? args_4 : _GEN_3955; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3957 = 3'h5 == total_offset_100 ? args_5 : _GEN_3956; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3958 = 3'h6 == total_offset_100 ? args_6 : _GEN_3957; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3959 = total_offset_100 < 3'h7 ? _GEN_3958 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_66_1 = 3'h0 < args_length_66 ? _GEN_3959 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_101 = args_offset_66 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3962 = 3'h1 == total_offset_101 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3963 = 3'h2 == total_offset_101 ? args_2 : _GEN_3962; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3964 = 3'h3 == total_offset_101 ? args_3 : _GEN_3963; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3965 = 3'h4 == total_offset_101 ? args_4 : _GEN_3964; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3966 = 3'h5 == total_offset_101 ? args_5 : _GEN_3965; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3967 = 3'h6 == total_offset_101 ? args_6 : _GEN_3966; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3968 = total_offset_101 < 3'h7 ? _GEN_3967 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_66_0 = 3'h1 < args_length_66 ? _GEN_3968 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1800 = {field_bytes_66_0,field_bytes_66_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_3970 = opcode_66 == 4'ha ? _field_data_T_1800 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3971 = opcode_66 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3191 = opcode_66 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_34 = field_data_lo_34[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1803 = {field_data_hi_34,field_data_lo_34}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_133 = _T_3191 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_3972 = opcode_66 == 4'h8 | opcode_66 == 4'hb ? _field_data_T_1803 : _GEN_3970; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3973 = opcode_66 == 4'h8 | opcode_66 == 4'hb ? _field_tag_T_133 : _GEN_3971; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_3974 = 14'h20 == field_data_lo_34 ? _field_data_T_36 : _GEN_3972; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3975 = 14'h21 == field_data_lo_34 ? _field_data_T_37 : _GEN_3974; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3976 = 14'h22 == field_data_lo_34 ? _field_data_T_38 : _GEN_3975; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3977 = 14'h23 == field_data_lo_34 ? _field_data_T_39 : _GEN_3976; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3978 = 14'h24 == field_data_lo_34 ? _field_data_T_40 : _GEN_3977; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3979 = 14'h25 == field_data_lo_34 ? _field_data_T_41 : _GEN_3978; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3980 = 14'h26 == field_data_lo_34 ? _field_data_T_42 : _GEN_3979; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3981 = 14'h27 == field_data_lo_34 ? _field_data_T_43 : _GEN_3980; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3982 = 14'h28 == field_data_lo_34 ? _field_data_T_44 : _GEN_3981; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3983 = 14'h29 == field_data_lo_34 ? _field_data_T_45 : _GEN_3982; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3984 = 14'h2a == field_data_lo_34 ? _field_data_T_46 : _GEN_3983; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3985 = 14'h2b == field_data_lo_34 ? _field_data_T_47 : _GEN_3984; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3986 = 14'h2c == field_data_lo_34 ? _field_data_T_48 : _GEN_3985; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3987 = 14'h2d == field_data_lo_34 ? _field_data_T_49 : _GEN_3986; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3988 = 14'h2e == field_data_lo_34 ? _field_data_T_50 : _GEN_3987; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3989 = 14'h2f == field_data_lo_34 ? _field_data_T_51 : _GEN_3988; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3990 = 14'h30 == field_data_lo_34 ? _field_data_T_52 : _GEN_3989; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3991 = 14'h31 == field_data_lo_34 ? _field_data_T_53 : _GEN_3990; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3992 = 14'h32 == field_data_lo_34 ? _field_data_T_54 : _GEN_3991; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3993 = 14'h33 == field_data_lo_34 ? _field_data_T_55 : _GEN_3992; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3994 = 14'h34 == field_data_lo_34 ? _field_data_T_56 : _GEN_3993; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3995 = 14'h35 == field_data_lo_34 ? _field_data_T_57 : _GEN_3994; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3996 = 14'h36 == field_data_lo_34 ? _field_data_T_58 : _GEN_3995; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3997 = 14'h37 == field_data_lo_34 ? _field_data_T_59 : _GEN_3996; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3998 = 14'h38 == field_data_lo_34 ? _field_data_T_60 : _GEN_3997; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_3999 = 14'h39 == field_data_lo_34 ? _field_data_T_61 : _GEN_3998; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4000 = 14'h3a == field_data_lo_34 ? _field_data_T_62 : _GEN_3999; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4001 = 14'h3b == field_data_lo_34 ? _field_data_T_63 : _GEN_4000; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4002 = 14'h3c == field_data_lo_34 ? _field_data_T_64 : _GEN_4001; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4003 = 14'h3d == field_data_lo_34 ? _field_data_T_65 : _GEN_4002; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4004 = 14'h3e == field_data_lo_34 ? _field_data_T_66 : _GEN_4003; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4005 = 14'h3f == field_data_lo_34 ? _field_data_T_67 : _GEN_4004; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4006 = 14'h40 == field_data_lo_34 ? _field_data_T_68 : _GEN_4005; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4007 = 14'h41 == field_data_lo_34 ? _field_data_T_69 : _GEN_4006; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4008 = 14'h42 == field_data_lo_34 ? _field_data_T_70 : _GEN_4007; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4009 = 14'h43 == field_data_lo_34 ? _field_data_T_71 : _GEN_4008; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4010 = 14'h44 == field_data_lo_34 ? _field_data_T_72 : _GEN_4009; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4011 = 14'h45 == field_data_lo_34 ? _field_data_T_73 : _GEN_4010; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4012 = 14'h46 == field_data_lo_34 ? _field_data_T_74 : _GEN_4011; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4013 = 14'h47 == field_data_lo_34 ? _field_data_T_75 : _GEN_4012; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4014 = 14'h48 == field_data_lo_34 ? _field_data_T_76 : _GEN_4013; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4015 = 14'h49 == field_data_lo_34 ? _field_data_T_77 : _GEN_4014; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4016 = 14'h4a == field_data_lo_34 ? _field_data_T_78 : _GEN_4015; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4017 = 14'h4b == field_data_lo_34 ? _field_data_T_79 : _GEN_4016; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4018 = 14'h4c == field_data_lo_34 ? _field_data_T_80 : _GEN_4017; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4019 = 14'h4d == field_data_lo_34 ? _field_data_T_81 : _GEN_4018; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4020 = 14'h4e == field_data_lo_34 ? _field_data_T_82 : _GEN_4019; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4021 = 14'h4f == field_data_lo_34 ? _field_data_T_83 : _GEN_4020; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_67 = vliw_67[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_35 = vliw_67[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_67 = field_data_lo_35[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_67 = field_data_lo_35[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_102 = {{1'd0}, args_offset_67}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_102 = _total_offset_T_102[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_4025 = 3'h1 == total_offset_102 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4026 = 3'h2 == total_offset_102 ? args_2 : _GEN_4025; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4027 = 3'h3 == total_offset_102 ? args_3 : _GEN_4026; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4028 = 3'h4 == total_offset_102 ? args_4 : _GEN_4027; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4029 = 3'h5 == total_offset_102 ? args_5 : _GEN_4028; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4030 = 3'h6 == total_offset_102 ? args_6 : _GEN_4029; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4031 = total_offset_102 < 3'h7 ? _GEN_4030 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_67_1 = 3'h0 < args_length_67 ? _GEN_4031 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_103 = args_offset_67 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_4034 = 3'h1 == total_offset_103 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4035 = 3'h2 == total_offset_103 ? args_2 : _GEN_4034; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4036 = 3'h3 == total_offset_103 ? args_3 : _GEN_4035; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4037 = 3'h4 == total_offset_103 ? args_4 : _GEN_4036; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4038 = 3'h5 == total_offset_103 ? args_5 : _GEN_4037; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4039 = 3'h6 == total_offset_103 ? args_6 : _GEN_4038; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4040 = total_offset_103 < 3'h7 ? _GEN_4039 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_67_0 = 3'h1 < args_length_67 ? _GEN_4040 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1852 = {field_bytes_67_0,field_bytes_67_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_4042 = opcode_67 == 4'ha ? _field_data_T_1852 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_4043 = opcode_67 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3248 = opcode_67 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_35 = field_data_lo_35[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1855 = {field_data_hi_35,field_data_lo_35}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_135 = _T_3248 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_4044 = opcode_67 == 4'h8 | opcode_67 == 4'hb ? _field_data_T_1855 : _GEN_4042; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_4045 = opcode_67 == 4'h8 | opcode_67 == 4'hb ? _field_tag_T_135 : _GEN_4043; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_4046 = 14'h20 == field_data_lo_35 ? _field_data_T_36 : _GEN_4044; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4047 = 14'h21 == field_data_lo_35 ? _field_data_T_37 : _GEN_4046; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4048 = 14'h22 == field_data_lo_35 ? _field_data_T_38 : _GEN_4047; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4049 = 14'h23 == field_data_lo_35 ? _field_data_T_39 : _GEN_4048; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4050 = 14'h24 == field_data_lo_35 ? _field_data_T_40 : _GEN_4049; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4051 = 14'h25 == field_data_lo_35 ? _field_data_T_41 : _GEN_4050; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4052 = 14'h26 == field_data_lo_35 ? _field_data_T_42 : _GEN_4051; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4053 = 14'h27 == field_data_lo_35 ? _field_data_T_43 : _GEN_4052; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4054 = 14'h28 == field_data_lo_35 ? _field_data_T_44 : _GEN_4053; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4055 = 14'h29 == field_data_lo_35 ? _field_data_T_45 : _GEN_4054; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4056 = 14'h2a == field_data_lo_35 ? _field_data_T_46 : _GEN_4055; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4057 = 14'h2b == field_data_lo_35 ? _field_data_T_47 : _GEN_4056; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4058 = 14'h2c == field_data_lo_35 ? _field_data_T_48 : _GEN_4057; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4059 = 14'h2d == field_data_lo_35 ? _field_data_T_49 : _GEN_4058; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4060 = 14'h2e == field_data_lo_35 ? _field_data_T_50 : _GEN_4059; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4061 = 14'h2f == field_data_lo_35 ? _field_data_T_51 : _GEN_4060; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4062 = 14'h30 == field_data_lo_35 ? _field_data_T_52 : _GEN_4061; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4063 = 14'h31 == field_data_lo_35 ? _field_data_T_53 : _GEN_4062; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4064 = 14'h32 == field_data_lo_35 ? _field_data_T_54 : _GEN_4063; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4065 = 14'h33 == field_data_lo_35 ? _field_data_T_55 : _GEN_4064; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4066 = 14'h34 == field_data_lo_35 ? _field_data_T_56 : _GEN_4065; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4067 = 14'h35 == field_data_lo_35 ? _field_data_T_57 : _GEN_4066; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4068 = 14'h36 == field_data_lo_35 ? _field_data_T_58 : _GEN_4067; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4069 = 14'h37 == field_data_lo_35 ? _field_data_T_59 : _GEN_4068; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4070 = 14'h38 == field_data_lo_35 ? _field_data_T_60 : _GEN_4069; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4071 = 14'h39 == field_data_lo_35 ? _field_data_T_61 : _GEN_4070; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4072 = 14'h3a == field_data_lo_35 ? _field_data_T_62 : _GEN_4071; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4073 = 14'h3b == field_data_lo_35 ? _field_data_T_63 : _GEN_4072; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4074 = 14'h3c == field_data_lo_35 ? _field_data_T_64 : _GEN_4073; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4075 = 14'h3d == field_data_lo_35 ? _field_data_T_65 : _GEN_4074; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4076 = 14'h3e == field_data_lo_35 ? _field_data_T_66 : _GEN_4075; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4077 = 14'h3f == field_data_lo_35 ? _field_data_T_67 : _GEN_4076; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4078 = 14'h40 == field_data_lo_35 ? _field_data_T_68 : _GEN_4077; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4079 = 14'h41 == field_data_lo_35 ? _field_data_T_69 : _GEN_4078; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4080 = 14'h42 == field_data_lo_35 ? _field_data_T_70 : _GEN_4079; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4081 = 14'h43 == field_data_lo_35 ? _field_data_T_71 : _GEN_4080; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4082 = 14'h44 == field_data_lo_35 ? _field_data_T_72 : _GEN_4081; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4083 = 14'h45 == field_data_lo_35 ? _field_data_T_73 : _GEN_4082; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4084 = 14'h46 == field_data_lo_35 ? _field_data_T_74 : _GEN_4083; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4085 = 14'h47 == field_data_lo_35 ? _field_data_T_75 : _GEN_4084; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4086 = 14'h48 == field_data_lo_35 ? _field_data_T_76 : _GEN_4085; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4087 = 14'h49 == field_data_lo_35 ? _field_data_T_77 : _GEN_4086; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4088 = 14'h4a == field_data_lo_35 ? _field_data_T_78 : _GEN_4087; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4089 = 14'h4b == field_data_lo_35 ? _field_data_T_79 : _GEN_4088; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4090 = 14'h4c == field_data_lo_35 ? _field_data_T_80 : _GEN_4089; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4091 = 14'h4d == field_data_lo_35 ? _field_data_T_81 : _GEN_4090; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4092 = 14'h4e == field_data_lo_35 ? _field_data_T_82 : _GEN_4091; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4093 = 14'h4f == field_data_lo_35 ? _field_data_T_83 : _GEN_4092; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_68 = vliw_68[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_36 = vliw_68[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_68 = field_data_lo_36[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_68 = field_data_lo_36[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_104 = {{1'd0}, args_offset_68}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_104 = _total_offset_T_104[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_4097 = 3'h1 == total_offset_104 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4098 = 3'h2 == total_offset_104 ? args_2 : _GEN_4097; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4099 = 3'h3 == total_offset_104 ? args_3 : _GEN_4098; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4100 = 3'h4 == total_offset_104 ? args_4 : _GEN_4099; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4101 = 3'h5 == total_offset_104 ? args_5 : _GEN_4100; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4102 = 3'h6 == total_offset_104 ? args_6 : _GEN_4101; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4103 = total_offset_104 < 3'h7 ? _GEN_4102 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_68_1 = 3'h0 < args_length_68 ? _GEN_4103 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_105 = args_offset_68 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_4106 = 3'h1 == total_offset_105 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4107 = 3'h2 == total_offset_105 ? args_2 : _GEN_4106; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4108 = 3'h3 == total_offset_105 ? args_3 : _GEN_4107; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4109 = 3'h4 == total_offset_105 ? args_4 : _GEN_4108; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4110 = 3'h5 == total_offset_105 ? args_5 : _GEN_4109; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4111 = 3'h6 == total_offset_105 ? args_6 : _GEN_4110; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4112 = total_offset_105 < 3'h7 ? _GEN_4111 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_68_0 = 3'h1 < args_length_68 ? _GEN_4112 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1904 = {field_bytes_68_0,field_bytes_68_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_4114 = opcode_68 == 4'ha ? _field_data_T_1904 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_4115 = opcode_68 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3305 = opcode_68 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_36 = field_data_lo_36[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1907 = {field_data_hi_36,field_data_lo_36}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_137 = _T_3305 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_4116 = opcode_68 == 4'h8 | opcode_68 == 4'hb ? _field_data_T_1907 : _GEN_4114; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_4117 = opcode_68 == 4'h8 | opcode_68 == 4'hb ? _field_tag_T_137 : _GEN_4115; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_4118 = 14'h20 == field_data_lo_36 ? _field_data_T_36 : _GEN_4116; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4119 = 14'h21 == field_data_lo_36 ? _field_data_T_37 : _GEN_4118; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4120 = 14'h22 == field_data_lo_36 ? _field_data_T_38 : _GEN_4119; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4121 = 14'h23 == field_data_lo_36 ? _field_data_T_39 : _GEN_4120; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4122 = 14'h24 == field_data_lo_36 ? _field_data_T_40 : _GEN_4121; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4123 = 14'h25 == field_data_lo_36 ? _field_data_T_41 : _GEN_4122; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4124 = 14'h26 == field_data_lo_36 ? _field_data_T_42 : _GEN_4123; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4125 = 14'h27 == field_data_lo_36 ? _field_data_T_43 : _GEN_4124; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4126 = 14'h28 == field_data_lo_36 ? _field_data_T_44 : _GEN_4125; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4127 = 14'h29 == field_data_lo_36 ? _field_data_T_45 : _GEN_4126; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4128 = 14'h2a == field_data_lo_36 ? _field_data_T_46 : _GEN_4127; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4129 = 14'h2b == field_data_lo_36 ? _field_data_T_47 : _GEN_4128; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4130 = 14'h2c == field_data_lo_36 ? _field_data_T_48 : _GEN_4129; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4131 = 14'h2d == field_data_lo_36 ? _field_data_T_49 : _GEN_4130; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4132 = 14'h2e == field_data_lo_36 ? _field_data_T_50 : _GEN_4131; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4133 = 14'h2f == field_data_lo_36 ? _field_data_T_51 : _GEN_4132; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4134 = 14'h30 == field_data_lo_36 ? _field_data_T_52 : _GEN_4133; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4135 = 14'h31 == field_data_lo_36 ? _field_data_T_53 : _GEN_4134; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4136 = 14'h32 == field_data_lo_36 ? _field_data_T_54 : _GEN_4135; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4137 = 14'h33 == field_data_lo_36 ? _field_data_T_55 : _GEN_4136; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4138 = 14'h34 == field_data_lo_36 ? _field_data_T_56 : _GEN_4137; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4139 = 14'h35 == field_data_lo_36 ? _field_data_T_57 : _GEN_4138; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4140 = 14'h36 == field_data_lo_36 ? _field_data_T_58 : _GEN_4139; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4141 = 14'h37 == field_data_lo_36 ? _field_data_T_59 : _GEN_4140; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4142 = 14'h38 == field_data_lo_36 ? _field_data_T_60 : _GEN_4141; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4143 = 14'h39 == field_data_lo_36 ? _field_data_T_61 : _GEN_4142; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4144 = 14'h3a == field_data_lo_36 ? _field_data_T_62 : _GEN_4143; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4145 = 14'h3b == field_data_lo_36 ? _field_data_T_63 : _GEN_4144; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4146 = 14'h3c == field_data_lo_36 ? _field_data_T_64 : _GEN_4145; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4147 = 14'h3d == field_data_lo_36 ? _field_data_T_65 : _GEN_4146; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4148 = 14'h3e == field_data_lo_36 ? _field_data_T_66 : _GEN_4147; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4149 = 14'h3f == field_data_lo_36 ? _field_data_T_67 : _GEN_4148; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4150 = 14'h40 == field_data_lo_36 ? _field_data_T_68 : _GEN_4149; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4151 = 14'h41 == field_data_lo_36 ? _field_data_T_69 : _GEN_4150; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4152 = 14'h42 == field_data_lo_36 ? _field_data_T_70 : _GEN_4151; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4153 = 14'h43 == field_data_lo_36 ? _field_data_T_71 : _GEN_4152; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4154 = 14'h44 == field_data_lo_36 ? _field_data_T_72 : _GEN_4153; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4155 = 14'h45 == field_data_lo_36 ? _field_data_T_73 : _GEN_4154; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4156 = 14'h46 == field_data_lo_36 ? _field_data_T_74 : _GEN_4155; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4157 = 14'h47 == field_data_lo_36 ? _field_data_T_75 : _GEN_4156; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4158 = 14'h48 == field_data_lo_36 ? _field_data_T_76 : _GEN_4157; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4159 = 14'h49 == field_data_lo_36 ? _field_data_T_77 : _GEN_4158; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4160 = 14'h4a == field_data_lo_36 ? _field_data_T_78 : _GEN_4159; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4161 = 14'h4b == field_data_lo_36 ? _field_data_T_79 : _GEN_4160; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4162 = 14'h4c == field_data_lo_36 ? _field_data_T_80 : _GEN_4161; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4163 = 14'h4d == field_data_lo_36 ? _field_data_T_81 : _GEN_4162; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4164 = 14'h4e == field_data_lo_36 ? _field_data_T_82 : _GEN_4163; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4165 = 14'h4f == field_data_lo_36 ? _field_data_T_83 : _GEN_4164; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_69 = vliw_69[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_37 = vliw_69[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_69 = field_data_lo_37[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_69 = field_data_lo_37[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_106 = {{1'd0}, args_offset_69}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_106 = _total_offset_T_106[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_4169 = 3'h1 == total_offset_106 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4170 = 3'h2 == total_offset_106 ? args_2 : _GEN_4169; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4171 = 3'h3 == total_offset_106 ? args_3 : _GEN_4170; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4172 = 3'h4 == total_offset_106 ? args_4 : _GEN_4171; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4173 = 3'h5 == total_offset_106 ? args_5 : _GEN_4172; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4174 = 3'h6 == total_offset_106 ? args_6 : _GEN_4173; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4175 = total_offset_106 < 3'h7 ? _GEN_4174 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_69_1 = 3'h0 < args_length_69 ? _GEN_4175 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_107 = args_offset_69 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_4178 = 3'h1 == total_offset_107 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4179 = 3'h2 == total_offset_107 ? args_2 : _GEN_4178; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4180 = 3'h3 == total_offset_107 ? args_3 : _GEN_4179; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4181 = 3'h4 == total_offset_107 ? args_4 : _GEN_4180; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4182 = 3'h5 == total_offset_107 ? args_5 : _GEN_4181; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4183 = 3'h6 == total_offset_107 ? args_6 : _GEN_4182; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4184 = total_offset_107 < 3'h7 ? _GEN_4183 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_69_0 = 3'h1 < args_length_69 ? _GEN_4184 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1956 = {field_bytes_69_0,field_bytes_69_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_4186 = opcode_69 == 4'ha ? _field_data_T_1956 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_4187 = opcode_69 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3362 = opcode_69 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_37 = field_data_lo_37[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1959 = {field_data_hi_37,field_data_lo_37}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_139 = _T_3362 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_4188 = opcode_69 == 4'h8 | opcode_69 == 4'hb ? _field_data_T_1959 : _GEN_4186; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_4189 = opcode_69 == 4'h8 | opcode_69 == 4'hb ? _field_tag_T_139 : _GEN_4187; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_4190 = 14'h20 == field_data_lo_37 ? _field_data_T_36 : _GEN_4188; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4191 = 14'h21 == field_data_lo_37 ? _field_data_T_37 : _GEN_4190; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4192 = 14'h22 == field_data_lo_37 ? _field_data_T_38 : _GEN_4191; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4193 = 14'h23 == field_data_lo_37 ? _field_data_T_39 : _GEN_4192; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4194 = 14'h24 == field_data_lo_37 ? _field_data_T_40 : _GEN_4193; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4195 = 14'h25 == field_data_lo_37 ? _field_data_T_41 : _GEN_4194; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4196 = 14'h26 == field_data_lo_37 ? _field_data_T_42 : _GEN_4195; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4197 = 14'h27 == field_data_lo_37 ? _field_data_T_43 : _GEN_4196; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4198 = 14'h28 == field_data_lo_37 ? _field_data_T_44 : _GEN_4197; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4199 = 14'h29 == field_data_lo_37 ? _field_data_T_45 : _GEN_4198; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4200 = 14'h2a == field_data_lo_37 ? _field_data_T_46 : _GEN_4199; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4201 = 14'h2b == field_data_lo_37 ? _field_data_T_47 : _GEN_4200; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4202 = 14'h2c == field_data_lo_37 ? _field_data_T_48 : _GEN_4201; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4203 = 14'h2d == field_data_lo_37 ? _field_data_T_49 : _GEN_4202; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4204 = 14'h2e == field_data_lo_37 ? _field_data_T_50 : _GEN_4203; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4205 = 14'h2f == field_data_lo_37 ? _field_data_T_51 : _GEN_4204; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4206 = 14'h30 == field_data_lo_37 ? _field_data_T_52 : _GEN_4205; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4207 = 14'h31 == field_data_lo_37 ? _field_data_T_53 : _GEN_4206; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4208 = 14'h32 == field_data_lo_37 ? _field_data_T_54 : _GEN_4207; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4209 = 14'h33 == field_data_lo_37 ? _field_data_T_55 : _GEN_4208; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4210 = 14'h34 == field_data_lo_37 ? _field_data_T_56 : _GEN_4209; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4211 = 14'h35 == field_data_lo_37 ? _field_data_T_57 : _GEN_4210; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4212 = 14'h36 == field_data_lo_37 ? _field_data_T_58 : _GEN_4211; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4213 = 14'h37 == field_data_lo_37 ? _field_data_T_59 : _GEN_4212; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4214 = 14'h38 == field_data_lo_37 ? _field_data_T_60 : _GEN_4213; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4215 = 14'h39 == field_data_lo_37 ? _field_data_T_61 : _GEN_4214; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4216 = 14'h3a == field_data_lo_37 ? _field_data_T_62 : _GEN_4215; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4217 = 14'h3b == field_data_lo_37 ? _field_data_T_63 : _GEN_4216; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4218 = 14'h3c == field_data_lo_37 ? _field_data_T_64 : _GEN_4217; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4219 = 14'h3d == field_data_lo_37 ? _field_data_T_65 : _GEN_4218; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4220 = 14'h3e == field_data_lo_37 ? _field_data_T_66 : _GEN_4219; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4221 = 14'h3f == field_data_lo_37 ? _field_data_T_67 : _GEN_4220; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4222 = 14'h40 == field_data_lo_37 ? _field_data_T_68 : _GEN_4221; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4223 = 14'h41 == field_data_lo_37 ? _field_data_T_69 : _GEN_4222; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4224 = 14'h42 == field_data_lo_37 ? _field_data_T_70 : _GEN_4223; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4225 = 14'h43 == field_data_lo_37 ? _field_data_T_71 : _GEN_4224; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4226 = 14'h44 == field_data_lo_37 ? _field_data_T_72 : _GEN_4225; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4227 = 14'h45 == field_data_lo_37 ? _field_data_T_73 : _GEN_4226; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4228 = 14'h46 == field_data_lo_37 ? _field_data_T_74 : _GEN_4227; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4229 = 14'h47 == field_data_lo_37 ? _field_data_T_75 : _GEN_4228; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4230 = 14'h48 == field_data_lo_37 ? _field_data_T_76 : _GEN_4229; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4231 = 14'h49 == field_data_lo_37 ? _field_data_T_77 : _GEN_4230; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4232 = 14'h4a == field_data_lo_37 ? _field_data_T_78 : _GEN_4231; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4233 = 14'h4b == field_data_lo_37 ? _field_data_T_79 : _GEN_4232; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4234 = 14'h4c == field_data_lo_37 ? _field_data_T_80 : _GEN_4233; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4235 = 14'h4d == field_data_lo_37 ? _field_data_T_81 : _GEN_4234; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4236 = 14'h4e == field_data_lo_37 ? _field_data_T_82 : _GEN_4235; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_4237 = 14'h4f == field_data_lo_37 ? _field_data_T_83 : _GEN_4236; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_160 = phv_data_160; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_161 = phv_data_161; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_162 = phv_data_162; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_163 = phv_data_163; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_164 = phv_data_164; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_165 = phv_data_165; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_166 = phv_data_166; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_167 = phv_data_167; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_168 = phv_data_168; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_169 = phv_data_169; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_170 = phv_data_170; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_171 = phv_data_171; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_172 = phv_data_172; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_173 = phv_data_173; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_174 = phv_data_174; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_175 = phv_data_175; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_176 = phv_data_176; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_177 = phv_data_177; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_178 = phv_data_178; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_179 = phv_data_179; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_180 = phv_data_180; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_181 = phv_data_181; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_182 = phv_data_182; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_183 = phv_data_183; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_184 = phv_data_184; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_185 = phv_data_185; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_186 = phv_data_186; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_187 = phv_data_187; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_188 = phv_data_188; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_189 = phv_data_189; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_190 = phv_data_190; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_191 = phv_data_191; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_192 = phv_data_192; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_193 = phv_data_193; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_194 = phv_data_194; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_195 = phv_data_195; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_196 = phv_data_196; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_197 = phv_data_197; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_198 = phv_data_198; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_199 = phv_data_199; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_200 = phv_data_200; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_201 = phv_data_201; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_202 = phv_data_202; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_203 = phv_data_203; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_204 = phv_data_204; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_205 = phv_data_205; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_206 = phv_data_206; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_207 = phv_data_207; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_208 = phv_data_208; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_209 = phv_data_209; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_210 = phv_data_210; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_211 = phv_data_211; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_212 = phv_data_212; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_213 = phv_data_213; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_214 = phv_data_214; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_215 = phv_data_215; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_216 = phv_data_216; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_217 = phv_data_217; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_218 = phv_data_218; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_219 = phv_data_219; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_220 = phv_data_220; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_221 = phv_data_221; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_222 = phv_data_222; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_223 = phv_data_223; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_224 = phv_data_224; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_225 = phv_data_225; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_226 = phv_data_226; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_227 = phv_data_227; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_228 = phv_data_228; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_229 = phv_data_229; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_230 = phv_data_230; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_231 = phv_data_231; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_232 = phv_data_232; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_233 = phv_data_233; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_234 = phv_data_234; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_235 = phv_data_235; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_236 = phv_data_236; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_237 = phv_data_237; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_238 = phv_data_238; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_239 = phv_data_239; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_240 = phv_data_240; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_241 = phv_data_241; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_242 = phv_data_242; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_243 = phv_data_243; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_244 = phv_data_244; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_245 = phv_data_245; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_246 = phv_data_246; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_247 = phv_data_247; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_248 = phv_data_248; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_249 = phv_data_249; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_250 = phv_data_250; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_251 = phv_data_251; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_252 = phv_data_252; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_253 = phv_data_253; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_254 = phv_data_254; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_255 = phv_data_255; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[executor_pisa.scala 163:25]
  assign io_nid_out = nid; // @[executor_pisa.scala 173:20]
  assign io_tag_out_0 = opcode == 4'h9 ? 2'h2 : _GEN_12; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_1 = opcode_1 == 4'h9 ? 2'h2 : _GEN_59; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_2 = opcode_2 == 4'h9 ? 2'h2 : _GEN_106; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_3 = opcode_3 == 4'h9 ? 2'h2 : _GEN_153; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_4 = opcode_4 == 4'h9 ? 2'h2 : _GEN_200; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_5 = opcode_5 == 4'h9 ? 2'h2 : _GEN_247; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_6 = opcode_6 == 4'h9 ? 2'h2 : _GEN_294; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_7 = opcode_7 == 4'h9 ? 2'h2 : _GEN_341; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_8 = opcode_8 == 4'h9 ? 2'h2 : _GEN_388; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_9 = opcode_9 == 4'h9 ? 2'h2 : _GEN_435; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_10 = opcode_10 == 4'h9 ? 2'h2 : _GEN_482; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_11 = opcode_11 == 4'h9 ? 2'h2 : _GEN_529; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_12 = opcode_12 == 4'h9 ? 2'h2 : _GEN_576; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_13 = opcode_13 == 4'h9 ? 2'h2 : _GEN_623; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_14 = opcode_14 == 4'h9 ? 2'h2 : _GEN_670; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_15 = opcode_15 == 4'h9 ? 2'h2 : _GEN_717; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_16 = opcode_16 == 4'h9 ? 2'h2 : _GEN_764; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_17 = opcode_17 == 4'h9 ? 2'h2 : _GEN_811; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_18 = opcode_18 == 4'h9 ? 2'h2 : _GEN_858; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_19 = opcode_19 == 4'h9 ? 2'h2 : _GEN_905; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_20 = opcode_20 == 4'h9 ? 2'h2 : _GEN_952; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_21 = opcode_21 == 4'h9 ? 2'h2 : _GEN_999; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_22 = opcode_22 == 4'h9 ? 2'h2 : _GEN_1046; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_23 = opcode_23 == 4'h9 ? 2'h2 : _GEN_1093; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_24 = opcode_24 == 4'h9 ? 2'h2 : _GEN_1140; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_25 = opcode_25 == 4'h9 ? 2'h2 : _GEN_1187; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_26 = opcode_26 == 4'h9 ? 2'h2 : _GEN_1234; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_27 = opcode_27 == 4'h9 ? 2'h2 : _GEN_1281; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_28 = opcode_28 == 4'h9 ? 2'h2 : _GEN_1328; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_29 = opcode_29 == 4'h9 ? 2'h2 : _GEN_1375; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_30 = opcode_30 == 4'h9 ? 2'h2 : _GEN_1422; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_31 = opcode_31 == 4'h9 ? 2'h2 : _GEN_1469; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_32 = opcode_32 == 4'h9 ? 2'h2 : _GEN_1525; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_33 = opcode_33 == 4'h9 ? 2'h2 : _GEN_1597; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_34 = opcode_34 == 4'h9 ? 2'h2 : _GEN_1669; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_35 = opcode_35 == 4'h9 ? 2'h2 : _GEN_1741; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_36 = opcode_36 == 4'h9 ? 2'h2 : _GEN_1813; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_37 = opcode_37 == 4'h9 ? 2'h2 : _GEN_1885; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_38 = opcode_38 == 4'h9 ? 2'h2 : _GEN_1957; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_39 = opcode_39 == 4'h9 ? 2'h2 : _GEN_2029; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_40 = opcode_40 == 4'h9 ? 2'h2 : _GEN_2101; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_41 = opcode_41 == 4'h9 ? 2'h2 : _GEN_2173; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_42 = opcode_42 == 4'h9 ? 2'h2 : _GEN_2245; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_43 = opcode_43 == 4'h9 ? 2'h2 : _GEN_2317; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_44 = opcode_44 == 4'h9 ? 2'h2 : _GEN_2389; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_45 = opcode_45 == 4'h9 ? 2'h2 : _GEN_2461; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_46 = opcode_46 == 4'h9 ? 2'h2 : _GEN_2533; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_47 = opcode_47 == 4'h9 ? 2'h2 : _GEN_2605; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_48 = opcode_48 == 4'h9 ? 2'h2 : _GEN_2677; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_49 = opcode_49 == 4'h9 ? 2'h2 : _GEN_2749; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_50 = opcode_50 == 4'h9 ? 2'h2 : _GEN_2821; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_51 = opcode_51 == 4'h9 ? 2'h2 : _GEN_2893; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_52 = opcode_52 == 4'h9 ? 2'h2 : _GEN_2965; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_53 = opcode_53 == 4'h9 ? 2'h2 : _GEN_3037; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_54 = opcode_54 == 4'h9 ? 2'h2 : _GEN_3109; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_55 = opcode_55 == 4'h9 ? 2'h2 : _GEN_3181; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_56 = opcode_56 == 4'h9 ? 2'h2 : _GEN_3253; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_57 = opcode_57 == 4'h9 ? 2'h2 : _GEN_3325; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_58 = opcode_58 == 4'h9 ? 2'h2 : _GEN_3397; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_59 = opcode_59 == 4'h9 ? 2'h2 : _GEN_3469; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_60 = opcode_60 == 4'h9 ? 2'h2 : _GEN_3541; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_61 = opcode_61 == 4'h9 ? 2'h2 : _GEN_3613; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_62 = opcode_62 == 4'h9 ? 2'h2 : _GEN_3685; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_63 = opcode_63 == 4'h9 ? 2'h2 : _GEN_3757; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_64 = opcode_64 == 4'h9 ? 2'h2 : _GEN_3829; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_65 = opcode_65 == 4'h9 ? 2'h2 : _GEN_3901; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_66 = opcode_66 == 4'h9 ? 2'h2 : _GEN_3973; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_67 = opcode_67 == 4'h9 ? 2'h2 : _GEN_4045; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_68 = opcode_68 == 4'h9 ? 2'h2 : _GEN_4117; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_69 = opcode_69 == 4'h9 ? 2'h2 : _GEN_4189; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_field_set_field8_0 = opcode == 4'h9 ? _GEN_44 : _GEN_11; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_1 = opcode_1 == 4'h9 ? _GEN_91 : _GEN_58; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_2 = opcode_2 == 4'h9 ? _GEN_138 : _GEN_105; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_3 = opcode_3 == 4'h9 ? _GEN_185 : _GEN_152; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_4 = opcode_4 == 4'h9 ? _GEN_232 : _GEN_199; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_5 = opcode_5 == 4'h9 ? _GEN_279 : _GEN_246; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_6 = opcode_6 == 4'h9 ? _GEN_326 : _GEN_293; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_7 = opcode_7 == 4'h9 ? _GEN_373 : _GEN_340; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_8 = opcode_8 == 4'h9 ? _GEN_420 : _GEN_387; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_9 = opcode_9 == 4'h9 ? _GEN_467 : _GEN_434; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_10 = opcode_10 == 4'h9 ? _GEN_514 : _GEN_481; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_11 = opcode_11 == 4'h9 ? _GEN_561 : _GEN_528; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_12 = opcode_12 == 4'h9 ? _GEN_608 : _GEN_575; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_13 = opcode_13 == 4'h9 ? _GEN_655 : _GEN_622; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_14 = opcode_14 == 4'h9 ? _GEN_702 : _GEN_669; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_15 = opcode_15 == 4'h9 ? _GEN_749 : _GEN_716; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_16 = opcode_16 == 4'h9 ? _GEN_796 : _GEN_763; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_17 = opcode_17 == 4'h9 ? _GEN_843 : _GEN_810; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_18 = opcode_18 == 4'h9 ? _GEN_890 : _GEN_857; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_19 = opcode_19 == 4'h9 ? _GEN_937 : _GEN_904; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_20 = opcode_20 == 4'h9 ? _GEN_984 : _GEN_951; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_21 = opcode_21 == 4'h9 ? _GEN_1031 : _GEN_998; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_22 = opcode_22 == 4'h9 ? _GEN_1078 : _GEN_1045; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_23 = opcode_23 == 4'h9 ? _GEN_1125 : _GEN_1092; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_24 = opcode_24 == 4'h9 ? _GEN_1172 : _GEN_1139; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_25 = opcode_25 == 4'h9 ? _GEN_1219 : _GEN_1186; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_26 = opcode_26 == 4'h9 ? _GEN_1266 : _GEN_1233; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_27 = opcode_27 == 4'h9 ? _GEN_1313 : _GEN_1280; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_28 = opcode_28 == 4'h9 ? _GEN_1360 : _GEN_1327; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_29 = opcode_29 == 4'h9 ? _GEN_1407 : _GEN_1374; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_30 = opcode_30 == 4'h9 ? _GEN_1454 : _GEN_1421; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_31 = opcode_31 == 4'h9 ? _GEN_1501 : _GEN_1468; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_0 = opcode_32 == 4'h9 ? _GEN_1573 : _GEN_1524; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_1 = opcode_33 == 4'h9 ? _GEN_1645 : _GEN_1596; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_2 = opcode_34 == 4'h9 ? _GEN_1717 : _GEN_1668; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_3 = opcode_35 == 4'h9 ? _GEN_1789 : _GEN_1740; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_4 = opcode_36 == 4'h9 ? _GEN_1861 : _GEN_1812; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_5 = opcode_37 == 4'h9 ? _GEN_1933 : _GEN_1884; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_6 = opcode_38 == 4'h9 ? _GEN_2005 : _GEN_1956; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_7 = opcode_39 == 4'h9 ? _GEN_2077 : _GEN_2028; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_8 = opcode_40 == 4'h9 ? _GEN_2149 : _GEN_2100; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_9 = opcode_41 == 4'h9 ? _GEN_2221 : _GEN_2172; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_10 = opcode_42 == 4'h9 ? _GEN_2293 : _GEN_2244; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_11 = opcode_43 == 4'h9 ? _GEN_2365 : _GEN_2316; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_12 = opcode_44 == 4'h9 ? _GEN_2437 : _GEN_2388; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_13 = opcode_45 == 4'h9 ? _GEN_2509 : _GEN_2460; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_14 = opcode_46 == 4'h9 ? _GEN_2581 : _GEN_2532; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_15 = opcode_47 == 4'h9 ? _GEN_2653 : _GEN_2604; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_16 = opcode_48 == 4'h9 ? _GEN_2725 : _GEN_2676; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_17 = opcode_49 == 4'h9 ? _GEN_2797 : _GEN_2748; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_18 = opcode_50 == 4'h9 ? _GEN_2869 : _GEN_2820; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_19 = opcode_51 == 4'h9 ? _GEN_2941 : _GEN_2892; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_20 = opcode_52 == 4'h9 ? _GEN_3013 : _GEN_2964; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_21 = opcode_53 == 4'h9 ? _GEN_3085 : _GEN_3036; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_22 = opcode_54 == 4'h9 ? _GEN_3157 : _GEN_3108; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_23 = opcode_55 == 4'h9 ? _GEN_3229 : _GEN_3180; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_24 = opcode_56 == 4'h9 ? _GEN_3301 : _GEN_3252; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_25 = opcode_57 == 4'h9 ? _GEN_3373 : _GEN_3324; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_26 = opcode_58 == 4'h9 ? _GEN_3445 : _GEN_3396; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_27 = opcode_59 == 4'h9 ? _GEN_3517 : _GEN_3468; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_28 = opcode_60 == 4'h9 ? _GEN_3589 : _GEN_3540; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_29 = opcode_61 == 4'h9 ? _GEN_3661 : _GEN_3612; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_30 = opcode_62 == 4'h9 ? _GEN_3733 : _GEN_3684; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_31 = opcode_63 == 4'h9 ? _GEN_3805 : _GEN_3756; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_32 = opcode_64 == 4'h9 ? _GEN_3877 : _GEN_3828; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_33 = opcode_65 == 4'h9 ? _GEN_3949 : _GEN_3900; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_34 = opcode_66 == 4'h9 ? _GEN_4021 : _GEN_3972; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_35 = opcode_67 == 4'h9 ? _GEN_4093 : _GEN_4044; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_36 = opcode_68 == 4'h9 ? _GEN_4165 : _GEN_4116; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_37 = opcode_69 == 4'h9 ? _GEN_4237 : _GEN_4188; // @[executor_pisa.scala 212:48]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[executor_pisa.scala 162:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[executor_pisa.scala 162:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[executor_pisa.scala 162:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[executor_pisa.scala 162:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[executor_pisa.scala 162:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[executor_pisa.scala 162:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[executor_pisa.scala 162:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[executor_pisa.scala 162:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[executor_pisa.scala 162:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[executor_pisa.scala 162:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[executor_pisa.scala 162:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[executor_pisa.scala 162:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[executor_pisa.scala 162:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[executor_pisa.scala 162:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[executor_pisa.scala 162:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[executor_pisa.scala 162:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[executor_pisa.scala 162:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[executor_pisa.scala 162:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[executor_pisa.scala 162:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[executor_pisa.scala 162:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[executor_pisa.scala 162:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[executor_pisa.scala 162:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[executor_pisa.scala 162:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[executor_pisa.scala 162:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[executor_pisa.scala 162:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[executor_pisa.scala 162:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[executor_pisa.scala 162:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[executor_pisa.scala 162:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[executor_pisa.scala 162:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[executor_pisa.scala 162:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[executor_pisa.scala 162:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[executor_pisa.scala 162:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[executor_pisa.scala 162:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[executor_pisa.scala 162:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[executor_pisa.scala 162:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[executor_pisa.scala 162:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[executor_pisa.scala 162:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[executor_pisa.scala 162:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[executor_pisa.scala 162:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[executor_pisa.scala 162:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[executor_pisa.scala 162:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[executor_pisa.scala 162:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[executor_pisa.scala 162:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[executor_pisa.scala 162:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[executor_pisa.scala 162:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[executor_pisa.scala 162:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[executor_pisa.scala 162:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[executor_pisa.scala 162:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[executor_pisa.scala 162:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[executor_pisa.scala 162:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[executor_pisa.scala 162:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[executor_pisa.scala 162:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[executor_pisa.scala 162:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[executor_pisa.scala 162:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[executor_pisa.scala 162:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[executor_pisa.scala 162:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[executor_pisa.scala 162:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[executor_pisa.scala 162:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[executor_pisa.scala 162:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[executor_pisa.scala 162:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[executor_pisa.scala 162:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[executor_pisa.scala 162:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[executor_pisa.scala 162:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[executor_pisa.scala 162:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[executor_pisa.scala 162:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[executor_pisa.scala 162:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[executor_pisa.scala 162:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[executor_pisa.scala 162:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[executor_pisa.scala 162:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[executor_pisa.scala 162:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[executor_pisa.scala 162:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[executor_pisa.scala 162:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[executor_pisa.scala 162:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[executor_pisa.scala 162:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[executor_pisa.scala 162:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[executor_pisa.scala 162:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[executor_pisa.scala 162:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[executor_pisa.scala 162:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[executor_pisa.scala 162:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[executor_pisa.scala 162:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[executor_pisa.scala 162:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[executor_pisa.scala 162:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[executor_pisa.scala 162:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[executor_pisa.scala 162:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[executor_pisa.scala 162:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[executor_pisa.scala 162:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[executor_pisa.scala 162:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[executor_pisa.scala 162:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[executor_pisa.scala 162:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[executor_pisa.scala 162:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[executor_pisa.scala 162:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[executor_pisa.scala 162:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[executor_pisa.scala 162:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[executor_pisa.scala 162:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[executor_pisa.scala 162:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[executor_pisa.scala 162:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[executor_pisa.scala 162:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[executor_pisa.scala 162:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[executor_pisa.scala 162:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[executor_pisa.scala 162:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[executor_pisa.scala 162:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[executor_pisa.scala 162:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[executor_pisa.scala 162:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[executor_pisa.scala 162:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[executor_pisa.scala 162:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[executor_pisa.scala 162:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[executor_pisa.scala 162:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[executor_pisa.scala 162:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[executor_pisa.scala 162:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[executor_pisa.scala 162:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[executor_pisa.scala 162:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[executor_pisa.scala 162:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[executor_pisa.scala 162:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[executor_pisa.scala 162:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[executor_pisa.scala 162:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[executor_pisa.scala 162:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[executor_pisa.scala 162:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[executor_pisa.scala 162:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[executor_pisa.scala 162:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[executor_pisa.scala 162:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[executor_pisa.scala 162:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[executor_pisa.scala 162:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[executor_pisa.scala 162:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[executor_pisa.scala 162:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[executor_pisa.scala 162:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[executor_pisa.scala 162:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[executor_pisa.scala 162:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[executor_pisa.scala 162:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[executor_pisa.scala 162:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[executor_pisa.scala 162:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[executor_pisa.scala 162:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[executor_pisa.scala 162:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[executor_pisa.scala 162:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[executor_pisa.scala 162:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[executor_pisa.scala 162:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[executor_pisa.scala 162:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[executor_pisa.scala 162:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[executor_pisa.scala 162:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[executor_pisa.scala 162:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[executor_pisa.scala 162:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[executor_pisa.scala 162:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[executor_pisa.scala 162:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[executor_pisa.scala 162:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[executor_pisa.scala 162:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[executor_pisa.scala 162:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[executor_pisa.scala 162:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[executor_pisa.scala 162:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[executor_pisa.scala 162:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[executor_pisa.scala 162:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[executor_pisa.scala 162:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[executor_pisa.scala 162:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[executor_pisa.scala 162:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[executor_pisa.scala 162:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[executor_pisa.scala 162:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[executor_pisa.scala 162:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[executor_pisa.scala 162:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[executor_pisa.scala 162:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[executor_pisa.scala 162:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[executor_pisa.scala 162:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[executor_pisa.scala 162:13]
    phv_data_160 <= io_pipe_phv_in_data_160; // @[executor_pisa.scala 162:13]
    phv_data_161 <= io_pipe_phv_in_data_161; // @[executor_pisa.scala 162:13]
    phv_data_162 <= io_pipe_phv_in_data_162; // @[executor_pisa.scala 162:13]
    phv_data_163 <= io_pipe_phv_in_data_163; // @[executor_pisa.scala 162:13]
    phv_data_164 <= io_pipe_phv_in_data_164; // @[executor_pisa.scala 162:13]
    phv_data_165 <= io_pipe_phv_in_data_165; // @[executor_pisa.scala 162:13]
    phv_data_166 <= io_pipe_phv_in_data_166; // @[executor_pisa.scala 162:13]
    phv_data_167 <= io_pipe_phv_in_data_167; // @[executor_pisa.scala 162:13]
    phv_data_168 <= io_pipe_phv_in_data_168; // @[executor_pisa.scala 162:13]
    phv_data_169 <= io_pipe_phv_in_data_169; // @[executor_pisa.scala 162:13]
    phv_data_170 <= io_pipe_phv_in_data_170; // @[executor_pisa.scala 162:13]
    phv_data_171 <= io_pipe_phv_in_data_171; // @[executor_pisa.scala 162:13]
    phv_data_172 <= io_pipe_phv_in_data_172; // @[executor_pisa.scala 162:13]
    phv_data_173 <= io_pipe_phv_in_data_173; // @[executor_pisa.scala 162:13]
    phv_data_174 <= io_pipe_phv_in_data_174; // @[executor_pisa.scala 162:13]
    phv_data_175 <= io_pipe_phv_in_data_175; // @[executor_pisa.scala 162:13]
    phv_data_176 <= io_pipe_phv_in_data_176; // @[executor_pisa.scala 162:13]
    phv_data_177 <= io_pipe_phv_in_data_177; // @[executor_pisa.scala 162:13]
    phv_data_178 <= io_pipe_phv_in_data_178; // @[executor_pisa.scala 162:13]
    phv_data_179 <= io_pipe_phv_in_data_179; // @[executor_pisa.scala 162:13]
    phv_data_180 <= io_pipe_phv_in_data_180; // @[executor_pisa.scala 162:13]
    phv_data_181 <= io_pipe_phv_in_data_181; // @[executor_pisa.scala 162:13]
    phv_data_182 <= io_pipe_phv_in_data_182; // @[executor_pisa.scala 162:13]
    phv_data_183 <= io_pipe_phv_in_data_183; // @[executor_pisa.scala 162:13]
    phv_data_184 <= io_pipe_phv_in_data_184; // @[executor_pisa.scala 162:13]
    phv_data_185 <= io_pipe_phv_in_data_185; // @[executor_pisa.scala 162:13]
    phv_data_186 <= io_pipe_phv_in_data_186; // @[executor_pisa.scala 162:13]
    phv_data_187 <= io_pipe_phv_in_data_187; // @[executor_pisa.scala 162:13]
    phv_data_188 <= io_pipe_phv_in_data_188; // @[executor_pisa.scala 162:13]
    phv_data_189 <= io_pipe_phv_in_data_189; // @[executor_pisa.scala 162:13]
    phv_data_190 <= io_pipe_phv_in_data_190; // @[executor_pisa.scala 162:13]
    phv_data_191 <= io_pipe_phv_in_data_191; // @[executor_pisa.scala 162:13]
    phv_data_192 <= io_pipe_phv_in_data_192; // @[executor_pisa.scala 162:13]
    phv_data_193 <= io_pipe_phv_in_data_193; // @[executor_pisa.scala 162:13]
    phv_data_194 <= io_pipe_phv_in_data_194; // @[executor_pisa.scala 162:13]
    phv_data_195 <= io_pipe_phv_in_data_195; // @[executor_pisa.scala 162:13]
    phv_data_196 <= io_pipe_phv_in_data_196; // @[executor_pisa.scala 162:13]
    phv_data_197 <= io_pipe_phv_in_data_197; // @[executor_pisa.scala 162:13]
    phv_data_198 <= io_pipe_phv_in_data_198; // @[executor_pisa.scala 162:13]
    phv_data_199 <= io_pipe_phv_in_data_199; // @[executor_pisa.scala 162:13]
    phv_data_200 <= io_pipe_phv_in_data_200; // @[executor_pisa.scala 162:13]
    phv_data_201 <= io_pipe_phv_in_data_201; // @[executor_pisa.scala 162:13]
    phv_data_202 <= io_pipe_phv_in_data_202; // @[executor_pisa.scala 162:13]
    phv_data_203 <= io_pipe_phv_in_data_203; // @[executor_pisa.scala 162:13]
    phv_data_204 <= io_pipe_phv_in_data_204; // @[executor_pisa.scala 162:13]
    phv_data_205 <= io_pipe_phv_in_data_205; // @[executor_pisa.scala 162:13]
    phv_data_206 <= io_pipe_phv_in_data_206; // @[executor_pisa.scala 162:13]
    phv_data_207 <= io_pipe_phv_in_data_207; // @[executor_pisa.scala 162:13]
    phv_data_208 <= io_pipe_phv_in_data_208; // @[executor_pisa.scala 162:13]
    phv_data_209 <= io_pipe_phv_in_data_209; // @[executor_pisa.scala 162:13]
    phv_data_210 <= io_pipe_phv_in_data_210; // @[executor_pisa.scala 162:13]
    phv_data_211 <= io_pipe_phv_in_data_211; // @[executor_pisa.scala 162:13]
    phv_data_212 <= io_pipe_phv_in_data_212; // @[executor_pisa.scala 162:13]
    phv_data_213 <= io_pipe_phv_in_data_213; // @[executor_pisa.scala 162:13]
    phv_data_214 <= io_pipe_phv_in_data_214; // @[executor_pisa.scala 162:13]
    phv_data_215 <= io_pipe_phv_in_data_215; // @[executor_pisa.scala 162:13]
    phv_data_216 <= io_pipe_phv_in_data_216; // @[executor_pisa.scala 162:13]
    phv_data_217 <= io_pipe_phv_in_data_217; // @[executor_pisa.scala 162:13]
    phv_data_218 <= io_pipe_phv_in_data_218; // @[executor_pisa.scala 162:13]
    phv_data_219 <= io_pipe_phv_in_data_219; // @[executor_pisa.scala 162:13]
    phv_data_220 <= io_pipe_phv_in_data_220; // @[executor_pisa.scala 162:13]
    phv_data_221 <= io_pipe_phv_in_data_221; // @[executor_pisa.scala 162:13]
    phv_data_222 <= io_pipe_phv_in_data_222; // @[executor_pisa.scala 162:13]
    phv_data_223 <= io_pipe_phv_in_data_223; // @[executor_pisa.scala 162:13]
    phv_data_224 <= io_pipe_phv_in_data_224; // @[executor_pisa.scala 162:13]
    phv_data_225 <= io_pipe_phv_in_data_225; // @[executor_pisa.scala 162:13]
    phv_data_226 <= io_pipe_phv_in_data_226; // @[executor_pisa.scala 162:13]
    phv_data_227 <= io_pipe_phv_in_data_227; // @[executor_pisa.scala 162:13]
    phv_data_228 <= io_pipe_phv_in_data_228; // @[executor_pisa.scala 162:13]
    phv_data_229 <= io_pipe_phv_in_data_229; // @[executor_pisa.scala 162:13]
    phv_data_230 <= io_pipe_phv_in_data_230; // @[executor_pisa.scala 162:13]
    phv_data_231 <= io_pipe_phv_in_data_231; // @[executor_pisa.scala 162:13]
    phv_data_232 <= io_pipe_phv_in_data_232; // @[executor_pisa.scala 162:13]
    phv_data_233 <= io_pipe_phv_in_data_233; // @[executor_pisa.scala 162:13]
    phv_data_234 <= io_pipe_phv_in_data_234; // @[executor_pisa.scala 162:13]
    phv_data_235 <= io_pipe_phv_in_data_235; // @[executor_pisa.scala 162:13]
    phv_data_236 <= io_pipe_phv_in_data_236; // @[executor_pisa.scala 162:13]
    phv_data_237 <= io_pipe_phv_in_data_237; // @[executor_pisa.scala 162:13]
    phv_data_238 <= io_pipe_phv_in_data_238; // @[executor_pisa.scala 162:13]
    phv_data_239 <= io_pipe_phv_in_data_239; // @[executor_pisa.scala 162:13]
    phv_data_240 <= io_pipe_phv_in_data_240; // @[executor_pisa.scala 162:13]
    phv_data_241 <= io_pipe_phv_in_data_241; // @[executor_pisa.scala 162:13]
    phv_data_242 <= io_pipe_phv_in_data_242; // @[executor_pisa.scala 162:13]
    phv_data_243 <= io_pipe_phv_in_data_243; // @[executor_pisa.scala 162:13]
    phv_data_244 <= io_pipe_phv_in_data_244; // @[executor_pisa.scala 162:13]
    phv_data_245 <= io_pipe_phv_in_data_245; // @[executor_pisa.scala 162:13]
    phv_data_246 <= io_pipe_phv_in_data_246; // @[executor_pisa.scala 162:13]
    phv_data_247 <= io_pipe_phv_in_data_247; // @[executor_pisa.scala 162:13]
    phv_data_248 <= io_pipe_phv_in_data_248; // @[executor_pisa.scala 162:13]
    phv_data_249 <= io_pipe_phv_in_data_249; // @[executor_pisa.scala 162:13]
    phv_data_250 <= io_pipe_phv_in_data_250; // @[executor_pisa.scala 162:13]
    phv_data_251 <= io_pipe_phv_in_data_251; // @[executor_pisa.scala 162:13]
    phv_data_252 <= io_pipe_phv_in_data_252; // @[executor_pisa.scala 162:13]
    phv_data_253 <= io_pipe_phv_in_data_253; // @[executor_pisa.scala 162:13]
    phv_data_254 <= io_pipe_phv_in_data_254; // @[executor_pisa.scala 162:13]
    phv_data_255 <= io_pipe_phv_in_data_255; // @[executor_pisa.scala 162:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[executor_pisa.scala 162:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[executor_pisa.scala 162:13]
    args_0 <= io_args_in_0; // @[executor_pisa.scala 166:14]
    args_1 <= io_args_in_1; // @[executor_pisa.scala 166:14]
    args_2 <= io_args_in_2; // @[executor_pisa.scala 166:14]
    args_3 <= io_args_in_3; // @[executor_pisa.scala 166:14]
    args_4 <= io_args_in_4; // @[executor_pisa.scala 166:14]
    args_5 <= io_args_in_5; // @[executor_pisa.scala 166:14]
    args_6 <= io_args_in_6; // @[executor_pisa.scala 166:14]
    vliw_0 <= io_vliw_in_0; // @[executor_pisa.scala 169:14]
    vliw_1 <= io_vliw_in_1; // @[executor_pisa.scala 169:14]
    vliw_2 <= io_vliw_in_2; // @[executor_pisa.scala 169:14]
    vliw_3 <= io_vliw_in_3; // @[executor_pisa.scala 169:14]
    vliw_4 <= io_vliw_in_4; // @[executor_pisa.scala 169:14]
    vliw_5 <= io_vliw_in_5; // @[executor_pisa.scala 169:14]
    vliw_6 <= io_vliw_in_6; // @[executor_pisa.scala 169:14]
    vliw_7 <= io_vliw_in_7; // @[executor_pisa.scala 169:14]
    vliw_8 <= io_vliw_in_8; // @[executor_pisa.scala 169:14]
    vliw_9 <= io_vliw_in_9; // @[executor_pisa.scala 169:14]
    vliw_10 <= io_vliw_in_10; // @[executor_pisa.scala 169:14]
    vliw_11 <= io_vliw_in_11; // @[executor_pisa.scala 169:14]
    vliw_12 <= io_vliw_in_12; // @[executor_pisa.scala 169:14]
    vliw_13 <= io_vliw_in_13; // @[executor_pisa.scala 169:14]
    vliw_14 <= io_vliw_in_14; // @[executor_pisa.scala 169:14]
    vliw_15 <= io_vliw_in_15; // @[executor_pisa.scala 169:14]
    vliw_16 <= io_vliw_in_16; // @[executor_pisa.scala 169:14]
    vliw_17 <= io_vliw_in_17; // @[executor_pisa.scala 169:14]
    vliw_18 <= io_vliw_in_18; // @[executor_pisa.scala 169:14]
    vliw_19 <= io_vliw_in_19; // @[executor_pisa.scala 169:14]
    vliw_20 <= io_vliw_in_20; // @[executor_pisa.scala 169:14]
    vliw_21 <= io_vliw_in_21; // @[executor_pisa.scala 169:14]
    vliw_22 <= io_vliw_in_22; // @[executor_pisa.scala 169:14]
    vliw_23 <= io_vliw_in_23; // @[executor_pisa.scala 169:14]
    vliw_24 <= io_vliw_in_24; // @[executor_pisa.scala 169:14]
    vliw_25 <= io_vliw_in_25; // @[executor_pisa.scala 169:14]
    vliw_26 <= io_vliw_in_26; // @[executor_pisa.scala 169:14]
    vliw_27 <= io_vliw_in_27; // @[executor_pisa.scala 169:14]
    vliw_28 <= io_vliw_in_28; // @[executor_pisa.scala 169:14]
    vliw_29 <= io_vliw_in_29; // @[executor_pisa.scala 169:14]
    vliw_30 <= io_vliw_in_30; // @[executor_pisa.scala 169:14]
    vliw_31 <= io_vliw_in_31; // @[executor_pisa.scala 169:14]
    vliw_32 <= io_vliw_in_32; // @[executor_pisa.scala 169:14]
    vliw_33 <= io_vliw_in_33; // @[executor_pisa.scala 169:14]
    vliw_34 <= io_vliw_in_34; // @[executor_pisa.scala 169:14]
    vliw_35 <= io_vliw_in_35; // @[executor_pisa.scala 169:14]
    vliw_36 <= io_vliw_in_36; // @[executor_pisa.scala 169:14]
    vliw_37 <= io_vliw_in_37; // @[executor_pisa.scala 169:14]
    vliw_38 <= io_vliw_in_38; // @[executor_pisa.scala 169:14]
    vliw_39 <= io_vliw_in_39; // @[executor_pisa.scala 169:14]
    vliw_40 <= io_vliw_in_40; // @[executor_pisa.scala 169:14]
    vliw_41 <= io_vliw_in_41; // @[executor_pisa.scala 169:14]
    vliw_42 <= io_vliw_in_42; // @[executor_pisa.scala 169:14]
    vliw_43 <= io_vliw_in_43; // @[executor_pisa.scala 169:14]
    vliw_44 <= io_vliw_in_44; // @[executor_pisa.scala 169:14]
    vliw_45 <= io_vliw_in_45; // @[executor_pisa.scala 169:14]
    vliw_46 <= io_vliw_in_46; // @[executor_pisa.scala 169:14]
    vliw_47 <= io_vliw_in_47; // @[executor_pisa.scala 169:14]
    vliw_48 <= io_vliw_in_48; // @[executor_pisa.scala 169:14]
    vliw_49 <= io_vliw_in_49; // @[executor_pisa.scala 169:14]
    vliw_50 <= io_vliw_in_50; // @[executor_pisa.scala 169:14]
    vliw_51 <= io_vliw_in_51; // @[executor_pisa.scala 169:14]
    vliw_52 <= io_vliw_in_52; // @[executor_pisa.scala 169:14]
    vliw_53 <= io_vliw_in_53; // @[executor_pisa.scala 169:14]
    vliw_54 <= io_vliw_in_54; // @[executor_pisa.scala 169:14]
    vliw_55 <= io_vliw_in_55; // @[executor_pisa.scala 169:14]
    vliw_56 <= io_vliw_in_56; // @[executor_pisa.scala 169:14]
    vliw_57 <= io_vliw_in_57; // @[executor_pisa.scala 169:14]
    vliw_58 <= io_vliw_in_58; // @[executor_pisa.scala 169:14]
    vliw_59 <= io_vliw_in_59; // @[executor_pisa.scala 169:14]
    vliw_60 <= io_vliw_in_60; // @[executor_pisa.scala 169:14]
    vliw_61 <= io_vliw_in_61; // @[executor_pisa.scala 169:14]
    vliw_62 <= io_vliw_in_62; // @[executor_pisa.scala 169:14]
    vliw_63 <= io_vliw_in_63; // @[executor_pisa.scala 169:14]
    vliw_64 <= io_vliw_in_64; // @[executor_pisa.scala 169:14]
    vliw_65 <= io_vliw_in_65; // @[executor_pisa.scala 169:14]
    vliw_66 <= io_vliw_in_66; // @[executor_pisa.scala 169:14]
    vliw_67 <= io_vliw_in_67; // @[executor_pisa.scala 169:14]
    vliw_68 <= io_vliw_in_68; // @[executor_pisa.scala 169:14]
    vliw_69 <= io_vliw_in_69; // @[executor_pisa.scala 169:14]
    nid <= io_nid_in; // @[executor_pisa.scala 172:13]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_data_160 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  phv_data_161 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  phv_data_162 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  phv_data_163 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  phv_data_164 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  phv_data_165 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  phv_data_166 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  phv_data_167 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  phv_data_168 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  phv_data_169 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  phv_data_170 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  phv_data_171 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  phv_data_172 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  phv_data_173 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  phv_data_174 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  phv_data_175 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  phv_data_176 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_data_177 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_data_178 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  phv_data_179 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  phv_data_180 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  phv_data_181 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  phv_data_182 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  phv_data_183 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  phv_data_184 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  phv_data_185 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  phv_data_186 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  phv_data_187 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  phv_data_188 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  phv_data_189 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  phv_data_190 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  phv_data_191 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  phv_data_192 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  phv_data_193 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  phv_data_194 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  phv_data_195 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  phv_data_196 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  phv_data_197 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  phv_data_198 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  phv_data_199 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  phv_data_200 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  phv_data_201 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  phv_data_202 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  phv_data_203 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  phv_data_204 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  phv_data_205 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  phv_data_206 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  phv_data_207 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  phv_data_208 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  phv_data_209 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  phv_data_210 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  phv_data_211 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  phv_data_212 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  phv_data_213 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  phv_data_214 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  phv_data_215 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  phv_data_216 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  phv_data_217 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  phv_data_218 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  phv_data_219 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  phv_data_220 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  phv_data_221 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  phv_data_222 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  phv_data_223 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  phv_data_224 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  phv_data_225 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  phv_data_226 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  phv_data_227 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  phv_data_228 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  phv_data_229 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  phv_data_230 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  phv_data_231 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  phv_data_232 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  phv_data_233 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  phv_data_234 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  phv_data_235 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  phv_data_236 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  phv_data_237 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  phv_data_238 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  phv_data_239 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  phv_data_240 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  phv_data_241 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  phv_data_242 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  phv_data_243 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  phv_data_244 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  phv_data_245 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  phv_data_246 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  phv_data_247 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  phv_data_248 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  phv_data_249 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  phv_data_250 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  phv_data_251 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  phv_data_252 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  phv_data_253 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  phv_data_254 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  phv_data_255 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_256[3:0];
  _RAND_257 = {1{`RANDOM}};
  phv_next_config_id = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  args_0 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  args_1 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  args_2 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  args_3 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  args_4 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  args_5 = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  args_6 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  vliw_0 = _RAND_265[17:0];
  _RAND_266 = {1{`RANDOM}};
  vliw_1 = _RAND_266[17:0];
  _RAND_267 = {1{`RANDOM}};
  vliw_2 = _RAND_267[17:0];
  _RAND_268 = {1{`RANDOM}};
  vliw_3 = _RAND_268[17:0];
  _RAND_269 = {1{`RANDOM}};
  vliw_4 = _RAND_269[17:0];
  _RAND_270 = {1{`RANDOM}};
  vliw_5 = _RAND_270[17:0];
  _RAND_271 = {1{`RANDOM}};
  vliw_6 = _RAND_271[17:0];
  _RAND_272 = {1{`RANDOM}};
  vliw_7 = _RAND_272[17:0];
  _RAND_273 = {1{`RANDOM}};
  vliw_8 = _RAND_273[17:0];
  _RAND_274 = {1{`RANDOM}};
  vliw_9 = _RAND_274[17:0];
  _RAND_275 = {1{`RANDOM}};
  vliw_10 = _RAND_275[17:0];
  _RAND_276 = {1{`RANDOM}};
  vliw_11 = _RAND_276[17:0];
  _RAND_277 = {1{`RANDOM}};
  vliw_12 = _RAND_277[17:0];
  _RAND_278 = {1{`RANDOM}};
  vliw_13 = _RAND_278[17:0];
  _RAND_279 = {1{`RANDOM}};
  vliw_14 = _RAND_279[17:0];
  _RAND_280 = {1{`RANDOM}};
  vliw_15 = _RAND_280[17:0];
  _RAND_281 = {1{`RANDOM}};
  vliw_16 = _RAND_281[17:0];
  _RAND_282 = {1{`RANDOM}};
  vliw_17 = _RAND_282[17:0];
  _RAND_283 = {1{`RANDOM}};
  vliw_18 = _RAND_283[17:0];
  _RAND_284 = {1{`RANDOM}};
  vliw_19 = _RAND_284[17:0];
  _RAND_285 = {1{`RANDOM}};
  vliw_20 = _RAND_285[17:0];
  _RAND_286 = {1{`RANDOM}};
  vliw_21 = _RAND_286[17:0];
  _RAND_287 = {1{`RANDOM}};
  vliw_22 = _RAND_287[17:0];
  _RAND_288 = {1{`RANDOM}};
  vliw_23 = _RAND_288[17:0];
  _RAND_289 = {1{`RANDOM}};
  vliw_24 = _RAND_289[17:0];
  _RAND_290 = {1{`RANDOM}};
  vliw_25 = _RAND_290[17:0];
  _RAND_291 = {1{`RANDOM}};
  vliw_26 = _RAND_291[17:0];
  _RAND_292 = {1{`RANDOM}};
  vliw_27 = _RAND_292[17:0];
  _RAND_293 = {1{`RANDOM}};
  vliw_28 = _RAND_293[17:0];
  _RAND_294 = {1{`RANDOM}};
  vliw_29 = _RAND_294[17:0];
  _RAND_295 = {1{`RANDOM}};
  vliw_30 = _RAND_295[17:0];
  _RAND_296 = {1{`RANDOM}};
  vliw_31 = _RAND_296[17:0];
  _RAND_297 = {1{`RANDOM}};
  vliw_32 = _RAND_297[17:0];
  _RAND_298 = {1{`RANDOM}};
  vliw_33 = _RAND_298[17:0];
  _RAND_299 = {1{`RANDOM}};
  vliw_34 = _RAND_299[17:0];
  _RAND_300 = {1{`RANDOM}};
  vliw_35 = _RAND_300[17:0];
  _RAND_301 = {1{`RANDOM}};
  vliw_36 = _RAND_301[17:0];
  _RAND_302 = {1{`RANDOM}};
  vliw_37 = _RAND_302[17:0];
  _RAND_303 = {1{`RANDOM}};
  vliw_38 = _RAND_303[17:0];
  _RAND_304 = {1{`RANDOM}};
  vliw_39 = _RAND_304[17:0];
  _RAND_305 = {1{`RANDOM}};
  vliw_40 = _RAND_305[17:0];
  _RAND_306 = {1{`RANDOM}};
  vliw_41 = _RAND_306[17:0];
  _RAND_307 = {1{`RANDOM}};
  vliw_42 = _RAND_307[17:0];
  _RAND_308 = {1{`RANDOM}};
  vliw_43 = _RAND_308[17:0];
  _RAND_309 = {1{`RANDOM}};
  vliw_44 = _RAND_309[17:0];
  _RAND_310 = {1{`RANDOM}};
  vliw_45 = _RAND_310[17:0];
  _RAND_311 = {1{`RANDOM}};
  vliw_46 = _RAND_311[17:0];
  _RAND_312 = {1{`RANDOM}};
  vliw_47 = _RAND_312[17:0];
  _RAND_313 = {1{`RANDOM}};
  vliw_48 = _RAND_313[17:0];
  _RAND_314 = {1{`RANDOM}};
  vliw_49 = _RAND_314[17:0];
  _RAND_315 = {1{`RANDOM}};
  vliw_50 = _RAND_315[17:0];
  _RAND_316 = {1{`RANDOM}};
  vliw_51 = _RAND_316[17:0];
  _RAND_317 = {1{`RANDOM}};
  vliw_52 = _RAND_317[17:0];
  _RAND_318 = {1{`RANDOM}};
  vliw_53 = _RAND_318[17:0];
  _RAND_319 = {1{`RANDOM}};
  vliw_54 = _RAND_319[17:0];
  _RAND_320 = {1{`RANDOM}};
  vliw_55 = _RAND_320[17:0];
  _RAND_321 = {1{`RANDOM}};
  vliw_56 = _RAND_321[17:0];
  _RAND_322 = {1{`RANDOM}};
  vliw_57 = _RAND_322[17:0];
  _RAND_323 = {1{`RANDOM}};
  vliw_58 = _RAND_323[17:0];
  _RAND_324 = {1{`RANDOM}};
  vliw_59 = _RAND_324[17:0];
  _RAND_325 = {1{`RANDOM}};
  vliw_60 = _RAND_325[17:0];
  _RAND_326 = {1{`RANDOM}};
  vliw_61 = _RAND_326[17:0];
  _RAND_327 = {1{`RANDOM}};
  vliw_62 = _RAND_327[17:0];
  _RAND_328 = {1{`RANDOM}};
  vliw_63 = _RAND_328[17:0];
  _RAND_329 = {1{`RANDOM}};
  vliw_64 = _RAND_329[17:0];
  _RAND_330 = {1{`RANDOM}};
  vliw_65 = _RAND_330[17:0];
  _RAND_331 = {1{`RANDOM}};
  vliw_66 = _RAND_331[17:0];
  _RAND_332 = {1{`RANDOM}};
  vliw_67 = _RAND_332[17:0];
  _RAND_333 = {1{`RANDOM}};
  vliw_68 = _RAND_333[17:0];
  _RAND_334 = {1{`RANDOM}};
  vliw_69 = _RAND_334[17:0];
  _RAND_335 = {1{`RANDOM}};
  nid = _RAND_335[14:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
