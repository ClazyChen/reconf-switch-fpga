module ParserPISA(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_valid,
  input         io_mod_en,
  input         io_mod_last_mau_id_mod,
  input  [3:0]  io_mod_last_mau_id,
  input  [2:0]  io_mod_cs,
  input         io_mod_module_mod_state_id_mod,
  input  [7:0]  io_mod_module_mod_state_id,
  input         io_mod_module_mod_sram_w_cs,
  input         io_mod_module_mod_sram_w_en,
  input  [7:0]  io_mod_module_mod_sram_w_addr,
  input  [63:0] io_mod_module_mod_sram_w_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  mau_0_clock; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_159; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_in_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_in_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_0_io_pipe_phv_in_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_0_io_pipe_phv_in_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_0_io_pipe_phv_in_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_0_io_pipe_phv_in_valid; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_159; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_0_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_0_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_0_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_0_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_0_io_pipe_phv_out_valid; // @[parser_pisa.scala 31:25]
  wire  mau_0_io_mod_state_id_mod; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_mod_state_id; // @[parser_pisa.scala 31:25]
  wire  mau_0_io_mod_sram_w_cs; // @[parser_pisa.scala 31:25]
  wire  mau_0_io_mod_sram_w_en; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_0_io_mod_sram_w_addr; // @[parser_pisa.scala 31:25]
  wire [63:0] mau_0_io_mod_sram_w_data; // @[parser_pisa.scala 31:25]
  wire  mau_1_clock; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_159; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_in_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_in_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_1_io_pipe_phv_in_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_1_io_pipe_phv_in_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_1_io_pipe_phv_in_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_1_io_pipe_phv_in_valid; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_159; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_1_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_1_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_1_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_1_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_1_io_pipe_phv_out_valid; // @[parser_pisa.scala 31:25]
  wire  mau_1_io_mod_state_id_mod; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_mod_state_id; // @[parser_pisa.scala 31:25]
  wire  mau_1_io_mod_sram_w_cs; // @[parser_pisa.scala 31:25]
  wire  mau_1_io_mod_sram_w_en; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_1_io_mod_sram_w_addr; // @[parser_pisa.scala 31:25]
  wire [63:0] mau_1_io_mod_sram_w_data; // @[parser_pisa.scala 31:25]
  wire  mau_2_clock; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_159; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_in_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_in_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_2_io_pipe_phv_in_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_2_io_pipe_phv_in_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_2_io_pipe_phv_in_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_2_io_pipe_phv_in_valid; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_159; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_2_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_2_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_2_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_2_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_2_io_pipe_phv_out_valid; // @[parser_pisa.scala 31:25]
  wire  mau_2_io_mod_state_id_mod; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_mod_state_id; // @[parser_pisa.scala 31:25]
  wire  mau_2_io_mod_sram_w_cs; // @[parser_pisa.scala 31:25]
  wire  mau_2_io_mod_sram_w_en; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_2_io_mod_sram_w_addr; // @[parser_pisa.scala 31:25]
  wire [63:0] mau_2_io_mod_sram_w_data; // @[parser_pisa.scala 31:25]
  wire  mau_3_clock; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_159; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_in_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_in_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_3_io_pipe_phv_in_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_3_io_pipe_phv_in_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_3_io_pipe_phv_in_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_3_io_pipe_phv_in_valid; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_159; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_3_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_3_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_3_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_3_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_3_io_pipe_phv_out_valid; // @[parser_pisa.scala 31:25]
  wire  mau_3_io_mod_state_id_mod; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_mod_state_id; // @[parser_pisa.scala 31:25]
  wire  mau_3_io_mod_sram_w_cs; // @[parser_pisa.scala 31:25]
  wire  mau_3_io_mod_sram_w_en; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_3_io_mod_sram_w_addr; // @[parser_pisa.scala 31:25]
  wire [63:0] mau_3_io_mod_sram_w_data; // @[parser_pisa.scala 31:25]
  wire  mau_4_clock; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_data_159; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_in_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_in_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_4_io_pipe_phv_in_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_4_io_pipe_phv_in_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_4_io_pipe_phv_in_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_4_io_pipe_phv_in_valid; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_data_159; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_4_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_4_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_4_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_4_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_4_io_pipe_phv_out_valid; // @[parser_pisa.scala 31:25]
  wire  mau_4_io_mod_state_id_mod; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_mod_state_id; // @[parser_pisa.scala 31:25]
  wire  mau_4_io_mod_sram_w_cs; // @[parser_pisa.scala 31:25]
  wire  mau_4_io_mod_sram_w_en; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_4_io_mod_sram_w_addr; // @[parser_pisa.scala 31:25]
  wire [63:0] mau_4_io_mod_sram_w_data; // @[parser_pisa.scala 31:25]
  wire  mau_5_clock; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_data_159; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_in_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_in_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_5_io_pipe_phv_in_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_5_io_pipe_phv_in_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_5_io_pipe_phv_in_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_5_io_pipe_phv_in_valid; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_data_159; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_5_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_5_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_5_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_5_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_5_io_pipe_phv_out_valid; // @[parser_pisa.scala 31:25]
  wire  mau_5_io_mod_state_id_mod; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_mod_state_id; // @[parser_pisa.scala 31:25]
  wire  mau_5_io_mod_sram_w_cs; // @[parser_pisa.scala 31:25]
  wire  mau_5_io_mod_sram_w_en; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_5_io_mod_sram_w_addr; // @[parser_pisa.scala 31:25]
  wire [63:0] mau_5_io_mod_sram_w_data; // @[parser_pisa.scala 31:25]
  wire  mau_6_clock; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_data_159; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_in_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_in_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_6_io_pipe_phv_in_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_6_io_pipe_phv_in_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_6_io_pipe_phv_in_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_6_io_pipe_phv_in_valid; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_data_159; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_6_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_6_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_6_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_6_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_6_io_pipe_phv_out_valid; // @[parser_pisa.scala 31:25]
  wire  mau_6_io_mod_state_id_mod; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_mod_state_id; // @[parser_pisa.scala 31:25]
  wire  mau_6_io_mod_sram_w_cs; // @[parser_pisa.scala 31:25]
  wire  mau_6_io_mod_sram_w_en; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_6_io_mod_sram_w_addr; // @[parser_pisa.scala 31:25]
  wire [63:0] mau_6_io_mod_sram_w_data; // @[parser_pisa.scala 31:25]
  wire  mau_7_clock; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_data_159; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_in_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_in_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_7_io_pipe_phv_in_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_7_io_pipe_phv_in_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_7_io_pipe_phv_in_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_7_io_pipe_phv_in_valid; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_0; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_1; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_2; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_3; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_4; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_5; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_6; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_7; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_8; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_9; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_10; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_11; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_12; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_13; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_14; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_16; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_17; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_18; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_19; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_20; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_21; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_22; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_23; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_24; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_25; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_26; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_27; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_28; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_29; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_30; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_31; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_32; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_33; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_34; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_35; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_36; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_37; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_38; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_39; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_40; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_41; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_42; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_43; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_44; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_45; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_46; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_47; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_48; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_49; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_50; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_51; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_52; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_53; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_54; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_55; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_56; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_57; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_58; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_59; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_60; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_61; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_62; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_63; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_64; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_65; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_66; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_67; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_68; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_69; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_70; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_71; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_72; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_73; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_74; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_75; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_76; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_77; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_78; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_79; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_80; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_81; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_82; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_83; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_84; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_85; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_86; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_87; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_88; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_89; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_90; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_91; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_92; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_93; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_94; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_95; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_96; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_97; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_98; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_99; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_100; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_101; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_102; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_103; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_104; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_105; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_106; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_107; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_108; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_109; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_110; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_111; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_112; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_113; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_114; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_115; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_116; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_117; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_118; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_119; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_120; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_121; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_122; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_123; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_124; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_125; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_126; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_127; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_128; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_129; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_130; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_131; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_132; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_133; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_134; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_135; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_136; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_137; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_138; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_139; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_140; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_141; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_142; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_143; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_144; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_145; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_146; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_147; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_148; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_149; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_150; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_151; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_152; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_153; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_154; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_155; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_156; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_157; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_158; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_data_159; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_0; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_1; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_2; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_3; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_4; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_5; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_6; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_7; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_8; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_9; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_10; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_11; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_12; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_13; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_14; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_header_15; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 31:25]
  wire [15:0] mau_7_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 31:25]
  wire [3:0] mau_7_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 31:25]
  wire  mau_7_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 31:25]
  wire  mau_7_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 31:25]
  wire  mau_7_io_pipe_phv_out_valid; // @[parser_pisa.scala 31:25]
  wire  mau_7_io_mod_state_id_mod; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_mod_state_id; // @[parser_pisa.scala 31:25]
  wire  mau_7_io_mod_sram_w_cs; // @[parser_pisa.scala 31:25]
  wire  mau_7_io_mod_sram_w_en; // @[parser_pisa.scala 31:25]
  wire [7:0] mau_7_io_mod_sram_w_addr; // @[parser_pisa.scala 31:25]
  wire [63:0] mau_7_io_mod_sram_w_data; // @[parser_pisa.scala 31:25]
  reg [3:0] last_mau_id; // @[parser_pisa.scala 24:26]
  wire  _GEN_0 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_valid : 1'h1; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire  _GEN_2 = 4'h1 == last_mau_id & mau_1_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [3:0] _GEN_3 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_next_processor_id : 4'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_23 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_0 : io_pipe_phv_in_data_0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_24 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_1 : io_pipe_phv_in_data_1; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_25 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_2 : io_pipe_phv_in_data_2; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_26 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_3 : io_pipe_phv_in_data_3; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_27 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_4 : io_pipe_phv_in_data_4; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_28 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_5 : io_pipe_phv_in_data_5; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_29 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_6 : io_pipe_phv_in_data_6; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_30 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_7 : io_pipe_phv_in_data_7; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_31 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_8 : io_pipe_phv_in_data_8; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_32 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_9 : io_pipe_phv_in_data_9; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_33 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_10 : io_pipe_phv_in_data_10; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_34 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_11 : io_pipe_phv_in_data_11; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_35 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_12 : io_pipe_phv_in_data_12; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_36 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_13 : io_pipe_phv_in_data_13; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_37 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_14 : io_pipe_phv_in_data_14; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_38 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_15 : io_pipe_phv_in_data_15; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_39 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_16 : io_pipe_phv_in_data_16; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_40 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_17 : io_pipe_phv_in_data_17; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_41 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_18 : io_pipe_phv_in_data_18; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_42 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_19 : io_pipe_phv_in_data_19; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_43 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_20 : io_pipe_phv_in_data_20; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_44 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_21 : io_pipe_phv_in_data_21; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_45 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_22 : io_pipe_phv_in_data_22; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_46 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_23 : io_pipe_phv_in_data_23; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_47 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_24 : io_pipe_phv_in_data_24; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_48 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_25 : io_pipe_phv_in_data_25; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_49 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_26 : io_pipe_phv_in_data_26; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_50 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_27 : io_pipe_phv_in_data_27; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_51 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_28 : io_pipe_phv_in_data_28; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_52 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_29 : io_pipe_phv_in_data_29; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_53 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_30 : io_pipe_phv_in_data_30; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_54 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_31 : io_pipe_phv_in_data_31; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_55 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_32 : io_pipe_phv_in_data_32; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_56 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_33 : io_pipe_phv_in_data_33; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_57 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_34 : io_pipe_phv_in_data_34; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_58 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_35 : io_pipe_phv_in_data_35; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_59 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_36 : io_pipe_phv_in_data_36; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_60 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_37 : io_pipe_phv_in_data_37; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_61 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_38 : io_pipe_phv_in_data_38; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_62 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_39 : io_pipe_phv_in_data_39; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_63 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_40 : io_pipe_phv_in_data_40; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_64 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_41 : io_pipe_phv_in_data_41; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_65 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_42 : io_pipe_phv_in_data_42; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_66 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_43 : io_pipe_phv_in_data_43; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_67 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_44 : io_pipe_phv_in_data_44; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_68 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_45 : io_pipe_phv_in_data_45; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_69 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_46 : io_pipe_phv_in_data_46; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_70 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_47 : io_pipe_phv_in_data_47; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_71 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_48 : io_pipe_phv_in_data_48; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_72 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_49 : io_pipe_phv_in_data_49; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_73 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_50 : io_pipe_phv_in_data_50; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_74 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_51 : io_pipe_phv_in_data_51; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_75 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_52 : io_pipe_phv_in_data_52; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_76 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_53 : io_pipe_phv_in_data_53; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_77 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_54 : io_pipe_phv_in_data_54; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_78 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_55 : io_pipe_phv_in_data_55; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_79 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_56 : io_pipe_phv_in_data_56; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_80 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_57 : io_pipe_phv_in_data_57; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_81 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_58 : io_pipe_phv_in_data_58; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_82 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_59 : io_pipe_phv_in_data_59; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_83 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_60 : io_pipe_phv_in_data_60; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_84 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_61 : io_pipe_phv_in_data_61; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_85 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_62 : io_pipe_phv_in_data_62; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_86 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_63 : io_pipe_phv_in_data_63; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_87 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_64 : io_pipe_phv_in_data_64; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_88 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_65 : io_pipe_phv_in_data_65; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_89 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_66 : io_pipe_phv_in_data_66; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_90 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_67 : io_pipe_phv_in_data_67; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_91 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_68 : io_pipe_phv_in_data_68; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_92 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_69 : io_pipe_phv_in_data_69; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_93 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_70 : io_pipe_phv_in_data_70; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_94 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_71 : io_pipe_phv_in_data_71; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_95 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_72 : io_pipe_phv_in_data_72; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_96 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_73 : io_pipe_phv_in_data_73; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_97 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_74 : io_pipe_phv_in_data_74; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_98 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_75 : io_pipe_phv_in_data_75; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_99 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_76 : io_pipe_phv_in_data_76; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_100 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_77 : io_pipe_phv_in_data_77; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_101 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_78 : io_pipe_phv_in_data_78; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_102 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_79 : io_pipe_phv_in_data_79; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_103 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_80 : io_pipe_phv_in_data_80; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_104 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_81 : io_pipe_phv_in_data_81; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_105 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_82 : io_pipe_phv_in_data_82; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_106 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_83 : io_pipe_phv_in_data_83; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_107 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_84 : io_pipe_phv_in_data_84; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_108 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_85 : io_pipe_phv_in_data_85; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_109 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_86 : io_pipe_phv_in_data_86; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_110 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_87 : io_pipe_phv_in_data_87; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_111 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_88 : io_pipe_phv_in_data_88; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_112 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_89 : io_pipe_phv_in_data_89; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_113 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_90 : io_pipe_phv_in_data_90; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_114 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_91 : io_pipe_phv_in_data_91; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_115 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_92 : io_pipe_phv_in_data_92; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_116 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_93 : io_pipe_phv_in_data_93; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_117 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_94 : io_pipe_phv_in_data_94; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_118 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_95 : io_pipe_phv_in_data_95; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_119 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_96 : io_pipe_phv_in_data_96; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_120 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_97 : io_pipe_phv_in_data_97; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_121 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_98 : io_pipe_phv_in_data_98; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_122 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_99 : io_pipe_phv_in_data_99; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_123 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_100 : io_pipe_phv_in_data_100; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_124 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_101 : io_pipe_phv_in_data_101; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_125 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_102 : io_pipe_phv_in_data_102; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_126 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_103 : io_pipe_phv_in_data_103; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_127 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_104 : io_pipe_phv_in_data_104; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_128 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_105 : io_pipe_phv_in_data_105; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_129 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_106 : io_pipe_phv_in_data_106; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_130 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_107 : io_pipe_phv_in_data_107; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_131 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_108 : io_pipe_phv_in_data_108; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_132 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_109 : io_pipe_phv_in_data_109; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_133 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_110 : io_pipe_phv_in_data_110; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_134 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_111 : io_pipe_phv_in_data_111; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_135 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_112 : io_pipe_phv_in_data_112; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_136 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_113 : io_pipe_phv_in_data_113; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_137 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_114 : io_pipe_phv_in_data_114; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_138 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_115 : io_pipe_phv_in_data_115; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_139 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_116 : io_pipe_phv_in_data_116; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_140 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_117 : io_pipe_phv_in_data_117; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_141 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_118 : io_pipe_phv_in_data_118; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_142 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_119 : io_pipe_phv_in_data_119; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_143 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_120 : io_pipe_phv_in_data_120; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_144 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_121 : io_pipe_phv_in_data_121; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_145 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_122 : io_pipe_phv_in_data_122; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_146 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_123 : io_pipe_phv_in_data_123; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_147 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_124 : io_pipe_phv_in_data_124; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_148 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_125 : io_pipe_phv_in_data_125; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_149 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_126 : io_pipe_phv_in_data_126; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_150 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_127 : io_pipe_phv_in_data_127; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_151 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_128 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_152 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_129 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_153 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_130 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_154 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_131 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_155 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_132 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_156 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_133 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_157 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_134 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_158 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_135 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_159 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_136 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_160 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_137 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_161 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_138 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_162 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_139 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_163 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_140 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_164 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_141 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_165 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_142 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_166 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_143 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_167 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_144 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_168 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_145 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_169 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_146 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_170 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_147 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_171 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_148 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_172 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_149 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_173 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_150 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_174 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_151 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_175 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_152 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_176 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_153 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_177 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_154 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_178 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_155 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_179 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_156 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_180 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_157 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_181 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_158 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire [7:0] _GEN_182 = 4'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_159 : 8'h0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35 parser_pisa.scala 36:21]
  wire  _GEN_183 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_valid : _GEN_0; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire  _GEN_185 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_next_config_id : _GEN_2; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [3:0] _GEN_186 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_next_processor_id : _GEN_3; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_206 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_0 : _GEN_23; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_207 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_1 : _GEN_24; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_208 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_2 : _GEN_25; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_209 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_3 : _GEN_26; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_210 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_4 : _GEN_27; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_211 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_5 : _GEN_28; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_212 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_6 : _GEN_29; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_213 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_7 : _GEN_30; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_214 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_8 : _GEN_31; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_215 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_9 : _GEN_32; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_216 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_10 : _GEN_33; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_217 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_11 : _GEN_34; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_218 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_12 : _GEN_35; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_219 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_13 : _GEN_36; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_220 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_14 : _GEN_37; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_221 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_15 : _GEN_38; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_222 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_16 : _GEN_39; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_223 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_17 : _GEN_40; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_224 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_18 : _GEN_41; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_225 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_19 : _GEN_42; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_226 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_20 : _GEN_43; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_227 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_21 : _GEN_44; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_228 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_22 : _GEN_45; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_229 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_23 : _GEN_46; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_230 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_24 : _GEN_47; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_231 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_25 : _GEN_48; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_232 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_26 : _GEN_49; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_233 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_27 : _GEN_50; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_234 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_28 : _GEN_51; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_235 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_29 : _GEN_52; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_236 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_30 : _GEN_53; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_237 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_31 : _GEN_54; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_238 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_32 : _GEN_55; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_239 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_33 : _GEN_56; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_240 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_34 : _GEN_57; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_241 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_35 : _GEN_58; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_242 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_36 : _GEN_59; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_243 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_37 : _GEN_60; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_244 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_38 : _GEN_61; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_245 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_39 : _GEN_62; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_246 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_40 : _GEN_63; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_247 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_41 : _GEN_64; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_248 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_42 : _GEN_65; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_249 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_43 : _GEN_66; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_250 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_44 : _GEN_67; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_251 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_45 : _GEN_68; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_252 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_46 : _GEN_69; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_253 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_47 : _GEN_70; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_254 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_48 : _GEN_71; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_255 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_49 : _GEN_72; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_256 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_50 : _GEN_73; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_257 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_51 : _GEN_74; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_258 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_52 : _GEN_75; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_259 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_53 : _GEN_76; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_260 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_54 : _GEN_77; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_261 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_55 : _GEN_78; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_262 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_56 : _GEN_79; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_263 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_57 : _GEN_80; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_264 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_58 : _GEN_81; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_265 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_59 : _GEN_82; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_266 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_60 : _GEN_83; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_267 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_61 : _GEN_84; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_268 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_62 : _GEN_85; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_269 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_63 : _GEN_86; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_270 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_64 : _GEN_87; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_271 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_65 : _GEN_88; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_272 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_66 : _GEN_89; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_273 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_67 : _GEN_90; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_274 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_68 : _GEN_91; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_275 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_69 : _GEN_92; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_276 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_70 : _GEN_93; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_277 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_71 : _GEN_94; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_278 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_72 : _GEN_95; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_279 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_73 : _GEN_96; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_280 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_74 : _GEN_97; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_281 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_75 : _GEN_98; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_282 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_76 : _GEN_99; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_283 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_77 : _GEN_100; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_284 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_78 : _GEN_101; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_285 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_79 : _GEN_102; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_286 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_80 : _GEN_103; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_287 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_81 : _GEN_104; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_288 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_82 : _GEN_105; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_289 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_83 : _GEN_106; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_290 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_84 : _GEN_107; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_291 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_85 : _GEN_108; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_292 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_86 : _GEN_109; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_293 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_87 : _GEN_110; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_294 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_88 : _GEN_111; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_295 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_89 : _GEN_112; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_296 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_90 : _GEN_113; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_297 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_91 : _GEN_114; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_298 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_92 : _GEN_115; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_299 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_93 : _GEN_116; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_300 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_94 : _GEN_117; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_301 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_95 : _GEN_118; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_302 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_96 : _GEN_119; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_303 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_97 : _GEN_120; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_304 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_98 : _GEN_121; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_305 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_99 : _GEN_122; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_306 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_100 : _GEN_123; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_307 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_101 : _GEN_124; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_308 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_102 : _GEN_125; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_309 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_103 : _GEN_126; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_310 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_104 : _GEN_127; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_311 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_105 : _GEN_128; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_312 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_106 : _GEN_129; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_313 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_107 : _GEN_130; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_314 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_108 : _GEN_131; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_315 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_109 : _GEN_132; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_316 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_110 : _GEN_133; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_317 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_111 : _GEN_134; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_318 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_112 : _GEN_135; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_319 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_113 : _GEN_136; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_320 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_114 : _GEN_137; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_321 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_115 : _GEN_138; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_322 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_116 : _GEN_139; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_323 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_117 : _GEN_140; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_324 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_118 : _GEN_141; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_325 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_119 : _GEN_142; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_326 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_120 : _GEN_143; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_327 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_121 : _GEN_144; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_328 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_122 : _GEN_145; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_329 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_123 : _GEN_146; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_330 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_124 : _GEN_147; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_331 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_125 : _GEN_148; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_332 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_126 : _GEN_149; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_333 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_127 : _GEN_150; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_334 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_128 : _GEN_151; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_335 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_129 : _GEN_152; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_336 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_130 : _GEN_153; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_337 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_131 : _GEN_154; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_338 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_132 : _GEN_155; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_339 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_133 : _GEN_156; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_340 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_134 : _GEN_157; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_341 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_135 : _GEN_158; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_342 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_136 : _GEN_159; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_343 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_137 : _GEN_160; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_344 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_138 : _GEN_161; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_345 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_139 : _GEN_162; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_346 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_140 : _GEN_163; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_347 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_141 : _GEN_164; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_348 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_142 : _GEN_165; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_349 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_143 : _GEN_166; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_350 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_144 : _GEN_167; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_351 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_145 : _GEN_168; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_352 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_146 : _GEN_169; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_353 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_147 : _GEN_170; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_354 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_148 : _GEN_171; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_355 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_149 : _GEN_172; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_356 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_150 : _GEN_173; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_357 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_151 : _GEN_174; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_358 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_152 : _GEN_175; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_359 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_153 : _GEN_176; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_360 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_154 : _GEN_177; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_361 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_155 : _GEN_178; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_362 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_156 : _GEN_179; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_363 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_157 : _GEN_180; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_364 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_158 : _GEN_181; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_365 = 4'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_159 : _GEN_182; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire  _GEN_366 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_valid : _GEN_183; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire  _GEN_368 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_next_config_id : _GEN_185; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [3:0] _GEN_369 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_next_processor_id : _GEN_186; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_389 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_0 : _GEN_206; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_390 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_1 : _GEN_207; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_391 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_2 : _GEN_208; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_392 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_3 : _GEN_209; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_393 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_4 : _GEN_210; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_394 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_5 : _GEN_211; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_395 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_6 : _GEN_212; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_396 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_7 : _GEN_213; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_397 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_8 : _GEN_214; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_398 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_9 : _GEN_215; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_399 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_10 : _GEN_216; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_400 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_11 : _GEN_217; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_401 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_12 : _GEN_218; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_402 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_13 : _GEN_219; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_403 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_14 : _GEN_220; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_404 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_15 : _GEN_221; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_405 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_16 : _GEN_222; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_406 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_17 : _GEN_223; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_407 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_18 : _GEN_224; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_408 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_19 : _GEN_225; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_409 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_20 : _GEN_226; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_410 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_21 : _GEN_227; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_411 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_22 : _GEN_228; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_412 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_23 : _GEN_229; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_413 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_24 : _GEN_230; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_414 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_25 : _GEN_231; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_415 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_26 : _GEN_232; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_416 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_27 : _GEN_233; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_417 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_28 : _GEN_234; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_418 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_29 : _GEN_235; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_419 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_30 : _GEN_236; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_420 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_31 : _GEN_237; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_421 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_32 : _GEN_238; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_422 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_33 : _GEN_239; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_423 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_34 : _GEN_240; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_424 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_35 : _GEN_241; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_425 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_36 : _GEN_242; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_426 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_37 : _GEN_243; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_427 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_38 : _GEN_244; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_428 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_39 : _GEN_245; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_429 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_40 : _GEN_246; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_430 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_41 : _GEN_247; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_431 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_42 : _GEN_248; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_432 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_43 : _GEN_249; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_433 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_44 : _GEN_250; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_434 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_45 : _GEN_251; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_435 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_46 : _GEN_252; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_436 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_47 : _GEN_253; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_437 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_48 : _GEN_254; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_438 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_49 : _GEN_255; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_439 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_50 : _GEN_256; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_440 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_51 : _GEN_257; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_441 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_52 : _GEN_258; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_442 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_53 : _GEN_259; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_443 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_54 : _GEN_260; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_444 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_55 : _GEN_261; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_445 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_56 : _GEN_262; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_446 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_57 : _GEN_263; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_447 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_58 : _GEN_264; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_448 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_59 : _GEN_265; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_449 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_60 : _GEN_266; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_450 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_61 : _GEN_267; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_451 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_62 : _GEN_268; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_452 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_63 : _GEN_269; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_453 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_64 : _GEN_270; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_454 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_65 : _GEN_271; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_455 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_66 : _GEN_272; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_456 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_67 : _GEN_273; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_457 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_68 : _GEN_274; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_458 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_69 : _GEN_275; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_459 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_70 : _GEN_276; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_460 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_71 : _GEN_277; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_461 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_72 : _GEN_278; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_462 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_73 : _GEN_279; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_463 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_74 : _GEN_280; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_464 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_75 : _GEN_281; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_465 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_76 : _GEN_282; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_466 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_77 : _GEN_283; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_467 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_78 : _GEN_284; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_468 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_79 : _GEN_285; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_469 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_80 : _GEN_286; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_470 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_81 : _GEN_287; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_471 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_82 : _GEN_288; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_472 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_83 : _GEN_289; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_473 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_84 : _GEN_290; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_474 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_85 : _GEN_291; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_475 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_86 : _GEN_292; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_476 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_87 : _GEN_293; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_477 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_88 : _GEN_294; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_478 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_89 : _GEN_295; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_479 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_90 : _GEN_296; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_480 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_91 : _GEN_297; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_481 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_92 : _GEN_298; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_482 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_93 : _GEN_299; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_483 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_94 : _GEN_300; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_484 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_95 : _GEN_301; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_485 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_96 : _GEN_302; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_486 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_97 : _GEN_303; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_487 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_98 : _GEN_304; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_488 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_99 : _GEN_305; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_489 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_100 : _GEN_306; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_490 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_101 : _GEN_307; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_491 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_102 : _GEN_308; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_492 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_103 : _GEN_309; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_493 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_104 : _GEN_310; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_494 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_105 : _GEN_311; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_495 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_106 : _GEN_312; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_496 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_107 : _GEN_313; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_497 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_108 : _GEN_314; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_498 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_109 : _GEN_315; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_499 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_110 : _GEN_316; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_500 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_111 : _GEN_317; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_501 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_112 : _GEN_318; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_502 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_113 : _GEN_319; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_503 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_114 : _GEN_320; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_504 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_115 : _GEN_321; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_505 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_116 : _GEN_322; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_506 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_117 : _GEN_323; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_507 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_118 : _GEN_324; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_508 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_119 : _GEN_325; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_509 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_120 : _GEN_326; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_510 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_121 : _GEN_327; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_511 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_122 : _GEN_328; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_512 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_123 : _GEN_329; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_513 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_124 : _GEN_330; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_514 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_125 : _GEN_331; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_515 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_126 : _GEN_332; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_516 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_127 : _GEN_333; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_517 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_128 : _GEN_334; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_518 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_129 : _GEN_335; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_519 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_130 : _GEN_336; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_520 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_131 : _GEN_337; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_521 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_132 : _GEN_338; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_522 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_133 : _GEN_339; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_523 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_134 : _GEN_340; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_524 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_135 : _GEN_341; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_525 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_136 : _GEN_342; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_526 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_137 : _GEN_343; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_527 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_138 : _GEN_344; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_528 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_139 : _GEN_345; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_529 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_140 : _GEN_346; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_530 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_141 : _GEN_347; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_531 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_142 : _GEN_348; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_532 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_143 : _GEN_349; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_533 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_144 : _GEN_350; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_534 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_145 : _GEN_351; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_535 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_146 : _GEN_352; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_536 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_147 : _GEN_353; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_537 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_148 : _GEN_354; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_538 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_149 : _GEN_355; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_539 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_150 : _GEN_356; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_540 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_151 : _GEN_357; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_541 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_152 : _GEN_358; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_542 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_153 : _GEN_359; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_543 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_154 : _GEN_360; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_544 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_155 : _GEN_361; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_545 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_156 : _GEN_362; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_546 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_157 : _GEN_363; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_547 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_158 : _GEN_364; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_548 = 4'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_159 : _GEN_365; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire  _GEN_549 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_valid : _GEN_366; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire  _GEN_551 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_next_config_id : _GEN_368; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [3:0] _GEN_552 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_next_processor_id : _GEN_369; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_572 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_0 : _GEN_389; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_573 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_1 : _GEN_390; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_574 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_2 : _GEN_391; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_575 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_3 : _GEN_392; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_576 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_4 : _GEN_393; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_577 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_5 : _GEN_394; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_578 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_6 : _GEN_395; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_579 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_7 : _GEN_396; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_580 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_8 : _GEN_397; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_581 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_9 : _GEN_398; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_582 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_10 : _GEN_399; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_583 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_11 : _GEN_400; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_584 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_12 : _GEN_401; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_585 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_13 : _GEN_402; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_586 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_14 : _GEN_403; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_587 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_15 : _GEN_404; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_588 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_16 : _GEN_405; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_589 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_17 : _GEN_406; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_590 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_18 : _GEN_407; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_591 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_19 : _GEN_408; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_592 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_20 : _GEN_409; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_593 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_21 : _GEN_410; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_594 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_22 : _GEN_411; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_595 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_23 : _GEN_412; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_596 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_24 : _GEN_413; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_597 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_25 : _GEN_414; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_598 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_26 : _GEN_415; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_599 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_27 : _GEN_416; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_600 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_28 : _GEN_417; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_601 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_29 : _GEN_418; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_602 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_30 : _GEN_419; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_603 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_31 : _GEN_420; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_604 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_32 : _GEN_421; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_605 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_33 : _GEN_422; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_606 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_34 : _GEN_423; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_607 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_35 : _GEN_424; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_608 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_36 : _GEN_425; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_609 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_37 : _GEN_426; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_610 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_38 : _GEN_427; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_611 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_39 : _GEN_428; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_612 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_40 : _GEN_429; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_613 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_41 : _GEN_430; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_614 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_42 : _GEN_431; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_615 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_43 : _GEN_432; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_616 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_44 : _GEN_433; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_617 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_45 : _GEN_434; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_618 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_46 : _GEN_435; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_619 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_47 : _GEN_436; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_620 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_48 : _GEN_437; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_621 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_49 : _GEN_438; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_622 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_50 : _GEN_439; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_623 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_51 : _GEN_440; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_624 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_52 : _GEN_441; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_625 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_53 : _GEN_442; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_626 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_54 : _GEN_443; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_627 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_55 : _GEN_444; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_628 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_56 : _GEN_445; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_629 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_57 : _GEN_446; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_630 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_58 : _GEN_447; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_631 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_59 : _GEN_448; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_632 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_60 : _GEN_449; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_633 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_61 : _GEN_450; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_634 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_62 : _GEN_451; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_635 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_63 : _GEN_452; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_636 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_64 : _GEN_453; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_637 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_65 : _GEN_454; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_638 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_66 : _GEN_455; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_639 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_67 : _GEN_456; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_640 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_68 : _GEN_457; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_641 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_69 : _GEN_458; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_642 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_70 : _GEN_459; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_643 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_71 : _GEN_460; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_644 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_72 : _GEN_461; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_645 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_73 : _GEN_462; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_646 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_74 : _GEN_463; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_647 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_75 : _GEN_464; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_648 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_76 : _GEN_465; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_649 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_77 : _GEN_466; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_650 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_78 : _GEN_467; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_651 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_79 : _GEN_468; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_652 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_80 : _GEN_469; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_653 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_81 : _GEN_470; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_654 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_82 : _GEN_471; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_655 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_83 : _GEN_472; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_656 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_84 : _GEN_473; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_657 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_85 : _GEN_474; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_658 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_86 : _GEN_475; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_659 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_87 : _GEN_476; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_660 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_88 : _GEN_477; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_661 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_89 : _GEN_478; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_662 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_90 : _GEN_479; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_663 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_91 : _GEN_480; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_664 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_92 : _GEN_481; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_665 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_93 : _GEN_482; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_666 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_94 : _GEN_483; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_667 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_95 : _GEN_484; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_668 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_96 : _GEN_485; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_669 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_97 : _GEN_486; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_670 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_98 : _GEN_487; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_671 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_99 : _GEN_488; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_672 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_100 : _GEN_489; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_673 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_101 : _GEN_490; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_674 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_102 : _GEN_491; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_675 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_103 : _GEN_492; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_676 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_104 : _GEN_493; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_677 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_105 : _GEN_494; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_678 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_106 : _GEN_495; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_679 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_107 : _GEN_496; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_680 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_108 : _GEN_497; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_681 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_109 : _GEN_498; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_682 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_110 : _GEN_499; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_683 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_111 : _GEN_500; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_684 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_112 : _GEN_501; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_685 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_113 : _GEN_502; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_686 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_114 : _GEN_503; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_687 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_115 : _GEN_504; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_688 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_116 : _GEN_505; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_689 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_117 : _GEN_506; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_690 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_118 : _GEN_507; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_691 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_119 : _GEN_508; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_692 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_120 : _GEN_509; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_693 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_121 : _GEN_510; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_694 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_122 : _GEN_511; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_695 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_123 : _GEN_512; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_696 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_124 : _GEN_513; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_697 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_125 : _GEN_514; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_698 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_126 : _GEN_515; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_699 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_127 : _GEN_516; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_700 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_128 : _GEN_517; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_701 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_129 : _GEN_518; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_702 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_130 : _GEN_519; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_703 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_131 : _GEN_520; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_704 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_132 : _GEN_521; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_705 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_133 : _GEN_522; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_706 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_134 : _GEN_523; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_707 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_135 : _GEN_524; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_708 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_136 : _GEN_525; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_709 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_137 : _GEN_526; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_710 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_138 : _GEN_527; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_711 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_139 : _GEN_528; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_712 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_140 : _GEN_529; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_713 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_141 : _GEN_530; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_714 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_142 : _GEN_531; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_715 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_143 : _GEN_532; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_716 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_144 : _GEN_533; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_717 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_145 : _GEN_534; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_718 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_146 : _GEN_535; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_719 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_147 : _GEN_536; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_720 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_148 : _GEN_537; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_721 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_149 : _GEN_538; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_722 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_150 : _GEN_539; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_723 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_151 : _GEN_540; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_724 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_152 : _GEN_541; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_725 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_153 : _GEN_542; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_726 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_154 : _GEN_543; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_727 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_155 : _GEN_544; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_728 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_156 : _GEN_545; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_729 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_157 : _GEN_546; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_730 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_158 : _GEN_547; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_731 = 4'h4 == last_mau_id ? mau_4_io_pipe_phv_out_data_159 : _GEN_548; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire  _GEN_732 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_valid : _GEN_549; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire  _GEN_734 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_next_config_id : _GEN_551; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [3:0] _GEN_735 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_next_processor_id : _GEN_552; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_755 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_0 : _GEN_572; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_756 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_1 : _GEN_573; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_757 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_2 : _GEN_574; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_758 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_3 : _GEN_575; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_759 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_4 : _GEN_576; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_760 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_5 : _GEN_577; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_761 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_6 : _GEN_578; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_762 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_7 : _GEN_579; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_763 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_8 : _GEN_580; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_764 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_9 : _GEN_581; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_765 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_10 : _GEN_582; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_766 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_11 : _GEN_583; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_767 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_12 : _GEN_584; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_768 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_13 : _GEN_585; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_769 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_14 : _GEN_586; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_770 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_15 : _GEN_587; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_771 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_16 : _GEN_588; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_772 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_17 : _GEN_589; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_773 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_18 : _GEN_590; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_774 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_19 : _GEN_591; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_775 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_20 : _GEN_592; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_776 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_21 : _GEN_593; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_777 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_22 : _GEN_594; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_778 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_23 : _GEN_595; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_779 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_24 : _GEN_596; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_780 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_25 : _GEN_597; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_781 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_26 : _GEN_598; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_782 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_27 : _GEN_599; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_783 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_28 : _GEN_600; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_784 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_29 : _GEN_601; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_785 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_30 : _GEN_602; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_786 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_31 : _GEN_603; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_787 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_32 : _GEN_604; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_788 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_33 : _GEN_605; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_789 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_34 : _GEN_606; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_790 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_35 : _GEN_607; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_791 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_36 : _GEN_608; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_792 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_37 : _GEN_609; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_793 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_38 : _GEN_610; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_794 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_39 : _GEN_611; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_795 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_40 : _GEN_612; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_796 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_41 : _GEN_613; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_797 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_42 : _GEN_614; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_798 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_43 : _GEN_615; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_799 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_44 : _GEN_616; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_800 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_45 : _GEN_617; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_801 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_46 : _GEN_618; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_802 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_47 : _GEN_619; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_803 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_48 : _GEN_620; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_804 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_49 : _GEN_621; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_805 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_50 : _GEN_622; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_806 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_51 : _GEN_623; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_807 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_52 : _GEN_624; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_808 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_53 : _GEN_625; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_809 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_54 : _GEN_626; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_810 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_55 : _GEN_627; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_811 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_56 : _GEN_628; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_812 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_57 : _GEN_629; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_813 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_58 : _GEN_630; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_814 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_59 : _GEN_631; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_815 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_60 : _GEN_632; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_816 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_61 : _GEN_633; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_817 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_62 : _GEN_634; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_818 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_63 : _GEN_635; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_819 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_64 : _GEN_636; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_820 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_65 : _GEN_637; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_821 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_66 : _GEN_638; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_822 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_67 : _GEN_639; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_823 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_68 : _GEN_640; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_824 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_69 : _GEN_641; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_825 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_70 : _GEN_642; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_826 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_71 : _GEN_643; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_827 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_72 : _GEN_644; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_828 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_73 : _GEN_645; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_829 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_74 : _GEN_646; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_830 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_75 : _GEN_647; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_831 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_76 : _GEN_648; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_832 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_77 : _GEN_649; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_833 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_78 : _GEN_650; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_834 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_79 : _GEN_651; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_835 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_80 : _GEN_652; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_836 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_81 : _GEN_653; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_837 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_82 : _GEN_654; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_838 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_83 : _GEN_655; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_839 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_84 : _GEN_656; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_840 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_85 : _GEN_657; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_841 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_86 : _GEN_658; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_842 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_87 : _GEN_659; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_843 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_88 : _GEN_660; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_844 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_89 : _GEN_661; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_845 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_90 : _GEN_662; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_846 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_91 : _GEN_663; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_847 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_92 : _GEN_664; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_848 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_93 : _GEN_665; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_849 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_94 : _GEN_666; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_850 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_95 : _GEN_667; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_851 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_96 : _GEN_668; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_852 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_97 : _GEN_669; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_853 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_98 : _GEN_670; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_854 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_99 : _GEN_671; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_855 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_100 : _GEN_672; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_856 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_101 : _GEN_673; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_857 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_102 : _GEN_674; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_858 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_103 : _GEN_675; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_859 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_104 : _GEN_676; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_860 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_105 : _GEN_677; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_861 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_106 : _GEN_678; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_862 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_107 : _GEN_679; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_863 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_108 : _GEN_680; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_864 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_109 : _GEN_681; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_865 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_110 : _GEN_682; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_866 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_111 : _GEN_683; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_867 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_112 : _GEN_684; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_868 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_113 : _GEN_685; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_869 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_114 : _GEN_686; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_870 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_115 : _GEN_687; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_871 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_116 : _GEN_688; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_872 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_117 : _GEN_689; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_873 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_118 : _GEN_690; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_874 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_119 : _GEN_691; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_875 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_120 : _GEN_692; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_876 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_121 : _GEN_693; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_877 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_122 : _GEN_694; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_878 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_123 : _GEN_695; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_879 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_124 : _GEN_696; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_880 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_125 : _GEN_697; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_881 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_126 : _GEN_698; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_882 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_127 : _GEN_699; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_883 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_128 : _GEN_700; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_884 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_129 : _GEN_701; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_885 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_130 : _GEN_702; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_886 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_131 : _GEN_703; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_887 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_132 : _GEN_704; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_888 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_133 : _GEN_705; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_889 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_134 : _GEN_706; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_890 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_135 : _GEN_707; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_891 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_136 : _GEN_708; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_892 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_137 : _GEN_709; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_893 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_138 : _GEN_710; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_894 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_139 : _GEN_711; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_895 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_140 : _GEN_712; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_896 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_141 : _GEN_713; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_897 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_142 : _GEN_714; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_898 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_143 : _GEN_715; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_899 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_144 : _GEN_716; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_900 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_145 : _GEN_717; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_901 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_146 : _GEN_718; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_902 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_147 : _GEN_719; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_903 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_148 : _GEN_720; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_904 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_149 : _GEN_721; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_905 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_150 : _GEN_722; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_906 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_151 : _GEN_723; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_907 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_152 : _GEN_724; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_908 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_153 : _GEN_725; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_909 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_154 : _GEN_726; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_910 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_155 : _GEN_727; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_911 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_156 : _GEN_728; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_912 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_157 : _GEN_729; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_913 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_158 : _GEN_730; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_914 = 4'h5 == last_mau_id ? mau_5_io_pipe_phv_out_data_159 : _GEN_731; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire  _GEN_915 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_valid : _GEN_732; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire  _GEN_917 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_next_config_id : _GEN_734; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [3:0] _GEN_918 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_next_processor_id : _GEN_735; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_938 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_0 : _GEN_755; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_939 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_1 : _GEN_756; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_940 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_2 : _GEN_757; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_941 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_3 : _GEN_758; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_942 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_4 : _GEN_759; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_943 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_5 : _GEN_760; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_944 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_6 : _GEN_761; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_945 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_7 : _GEN_762; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_946 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_8 : _GEN_763; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_947 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_9 : _GEN_764; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_948 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_10 : _GEN_765; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_949 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_11 : _GEN_766; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_950 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_12 : _GEN_767; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_951 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_13 : _GEN_768; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_952 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_14 : _GEN_769; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_953 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_15 : _GEN_770; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_954 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_16 : _GEN_771; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_955 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_17 : _GEN_772; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_956 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_18 : _GEN_773; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_957 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_19 : _GEN_774; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_958 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_20 : _GEN_775; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_959 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_21 : _GEN_776; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_960 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_22 : _GEN_777; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_961 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_23 : _GEN_778; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_962 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_24 : _GEN_779; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_963 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_25 : _GEN_780; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_964 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_26 : _GEN_781; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_965 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_27 : _GEN_782; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_966 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_28 : _GEN_783; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_967 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_29 : _GEN_784; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_968 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_30 : _GEN_785; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_969 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_31 : _GEN_786; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_970 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_32 : _GEN_787; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_971 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_33 : _GEN_788; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_972 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_34 : _GEN_789; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_973 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_35 : _GEN_790; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_974 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_36 : _GEN_791; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_975 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_37 : _GEN_792; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_976 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_38 : _GEN_793; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_977 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_39 : _GEN_794; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_978 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_40 : _GEN_795; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_979 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_41 : _GEN_796; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_980 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_42 : _GEN_797; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_981 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_43 : _GEN_798; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_982 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_44 : _GEN_799; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_983 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_45 : _GEN_800; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_984 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_46 : _GEN_801; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_985 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_47 : _GEN_802; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_986 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_48 : _GEN_803; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_987 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_49 : _GEN_804; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_988 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_50 : _GEN_805; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_989 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_51 : _GEN_806; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_990 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_52 : _GEN_807; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_991 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_53 : _GEN_808; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_992 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_54 : _GEN_809; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_993 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_55 : _GEN_810; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_994 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_56 : _GEN_811; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_995 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_57 : _GEN_812; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_996 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_58 : _GEN_813; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_997 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_59 : _GEN_814; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_998 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_60 : _GEN_815; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_999 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_61 : _GEN_816; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1000 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_62 : _GEN_817; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1001 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_63 : _GEN_818; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1002 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_64 : _GEN_819; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1003 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_65 : _GEN_820; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1004 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_66 : _GEN_821; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1005 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_67 : _GEN_822; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1006 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_68 : _GEN_823; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1007 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_69 : _GEN_824; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1008 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_70 : _GEN_825; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1009 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_71 : _GEN_826; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1010 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_72 : _GEN_827; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1011 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_73 : _GEN_828; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1012 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_74 : _GEN_829; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1013 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_75 : _GEN_830; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1014 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_76 : _GEN_831; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1015 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_77 : _GEN_832; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1016 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_78 : _GEN_833; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1017 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_79 : _GEN_834; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1018 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_80 : _GEN_835; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1019 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_81 : _GEN_836; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1020 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_82 : _GEN_837; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1021 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_83 : _GEN_838; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1022 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_84 : _GEN_839; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1023 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_85 : _GEN_840; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1024 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_86 : _GEN_841; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1025 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_87 : _GEN_842; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1026 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_88 : _GEN_843; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1027 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_89 : _GEN_844; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1028 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_90 : _GEN_845; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1029 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_91 : _GEN_846; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1030 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_92 : _GEN_847; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1031 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_93 : _GEN_848; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1032 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_94 : _GEN_849; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1033 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_95 : _GEN_850; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1034 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_96 : _GEN_851; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1035 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_97 : _GEN_852; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1036 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_98 : _GEN_853; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1037 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_99 : _GEN_854; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1038 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_100 : _GEN_855; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1039 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_101 : _GEN_856; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1040 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_102 : _GEN_857; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1041 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_103 : _GEN_858; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1042 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_104 : _GEN_859; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1043 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_105 : _GEN_860; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1044 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_106 : _GEN_861; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1045 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_107 : _GEN_862; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1046 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_108 : _GEN_863; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1047 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_109 : _GEN_864; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1048 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_110 : _GEN_865; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1049 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_111 : _GEN_866; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1050 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_112 : _GEN_867; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1051 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_113 : _GEN_868; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1052 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_114 : _GEN_869; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1053 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_115 : _GEN_870; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1054 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_116 : _GEN_871; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1055 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_117 : _GEN_872; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1056 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_118 : _GEN_873; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1057 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_119 : _GEN_874; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1058 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_120 : _GEN_875; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1059 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_121 : _GEN_876; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1060 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_122 : _GEN_877; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1061 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_123 : _GEN_878; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1062 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_124 : _GEN_879; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1063 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_125 : _GEN_880; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1064 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_126 : _GEN_881; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1065 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_127 : _GEN_882; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1066 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_128 : _GEN_883; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1067 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_129 : _GEN_884; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1068 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_130 : _GEN_885; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1069 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_131 : _GEN_886; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1070 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_132 : _GEN_887; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1071 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_133 : _GEN_888; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1072 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_134 : _GEN_889; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1073 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_135 : _GEN_890; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1074 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_136 : _GEN_891; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1075 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_137 : _GEN_892; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1076 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_138 : _GEN_893; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1077 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_139 : _GEN_894; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1078 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_140 : _GEN_895; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1079 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_141 : _GEN_896; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1080 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_142 : _GEN_897; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1081 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_143 : _GEN_898; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1082 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_144 : _GEN_899; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1083 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_145 : _GEN_900; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1084 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_146 : _GEN_901; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1085 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_147 : _GEN_902; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1086 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_148 : _GEN_903; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1087 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_149 : _GEN_904; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1088 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_150 : _GEN_905; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1089 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_151 : _GEN_906; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1090 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_152 : _GEN_907; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1091 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_153 : _GEN_908; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1092 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_154 : _GEN_909; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1093 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_155 : _GEN_910; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1094 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_156 : _GEN_911; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1095 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_157 : _GEN_912; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1096 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_158 : _GEN_913; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire [7:0] _GEN_1097 = 4'h6 == last_mau_id ? mau_6_io_pipe_phv_out_data_159 : _GEN_914; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  wire  mod_j = io_mod_cs == 3'h0; // @[parser_pisa.scala 56:35]
  wire  mod_j_1 = io_mod_cs == 3'h1; // @[parser_pisa.scala 56:35]
  wire  mod_j_2 = io_mod_cs == 3'h2; // @[parser_pisa.scala 56:35]
  wire  mod_j_3 = io_mod_cs == 3'h3; // @[parser_pisa.scala 56:35]
  wire  mod_j_4 = io_mod_cs == 3'h4; // @[parser_pisa.scala 56:35]
  wire  mod_j_5 = io_mod_cs == 3'h5; // @[parser_pisa.scala 56:35]
  wire  mod_j_6 = io_mod_cs == 3'h6; // @[parser_pisa.scala 56:35]
  wire  mod_j_7 = io_mod_cs == 3'h7; // @[parser_pisa.scala 56:35]
  ParseModule mau_0 ( // @[parser_pisa.scala 31:25]
    .clock(mau_0_clock),
    .io_pipe_phv_in_data_0(mau_0_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_0_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_0_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_0_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_0_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_0_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_0_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_0_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_0_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_0_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_0_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_0_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_0_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_0_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_0_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_0_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_0_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_0_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_0_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_0_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_0_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_0_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_0_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_0_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_0_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_0_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_0_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_0_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_0_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_0_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_0_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_0_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_0_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_0_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_0_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_0_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_0_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_0_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_0_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_0_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_0_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_0_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_0_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_0_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_0_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_0_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_0_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_0_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_0_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_0_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_0_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_0_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_0_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_0_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_0_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_0_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_0_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_0_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_0_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_0_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_0_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_0_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_0_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_0_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_0_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_0_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_0_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_0_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_0_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_0_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_0_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_0_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_0_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_0_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_0_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_0_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_0_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_0_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_0_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_0_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_0_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_0_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_0_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_0_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_0_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_0_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_0_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_0_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_0_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_0_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_0_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_0_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_0_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_0_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_0_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_0_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_0_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_0_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_0_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_0_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_0_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_0_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_0_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_0_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_0_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_0_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_0_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_0_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_0_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_0_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_0_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_0_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_0_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_0_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_0_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_0_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_0_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_0_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_0_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_0_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_0_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_0_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_0_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_0_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_0_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_0_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_0_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_0_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_0_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_0_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_0_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_0_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_0_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_0_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_0_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_0_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_0_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_0_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_0_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_0_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_0_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_0_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_0_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_0_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_0_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_0_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_0_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_0_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_0_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_0_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_0_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_0_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_0_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_0_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_0_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_0_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_0_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_0_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_0_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_0_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(mau_0_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_0_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_0_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_0_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_0_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_0_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_0_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_0_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_0_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_0_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_0_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_0_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_0_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_0_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_0_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_0_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_0_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_0_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_0_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_0_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_0_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_0_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(mau_0_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(mau_0_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_0_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_0_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_0_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_0_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_0_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_0_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_0_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_0_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_0_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_0_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_0_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_0_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_0_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_0_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_0_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_0_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_0_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_0_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_0_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_0_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_0_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_0_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_0_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_0_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_0_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_0_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_0_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_0_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_0_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_0_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_0_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_0_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_0_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_0_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_0_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_0_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_0_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_0_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_0_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_0_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_0_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_0_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_0_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_0_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_0_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_0_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_0_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_0_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_0_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_0_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_0_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_0_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_0_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_0_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_0_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_0_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_0_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_0_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_0_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_0_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_0_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_0_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_0_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_0_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_0_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_0_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_0_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_0_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_0_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_0_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_0_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_0_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_0_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_0_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_0_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_0_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_0_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_0_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_0_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_0_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_0_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_0_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_0_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_0_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_0_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_0_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_0_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_0_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_0_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_0_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_0_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_0_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_0_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_0_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_0_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_0_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_0_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_0_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_0_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_0_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_0_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_0_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_0_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_0_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_0_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_0_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_0_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_0_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_0_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_0_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_0_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_0_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_0_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_0_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_0_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_0_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_0_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_0_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_0_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_0_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_0_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_0_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_0_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_0_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_0_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_0_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_0_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_0_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_0_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_0_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_0_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_0_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_0_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_0_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_0_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_0_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_0_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_0_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_0_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_0_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_0_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_0_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_0_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_0_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_0_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_0_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_0_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_0_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_0_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_0_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_0_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_0_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_0_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_0_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_0_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_0_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_0_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_0_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_0_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(mau_0_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_0_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_0_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_0_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_0_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_0_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_0_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_0_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_0_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_0_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_0_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_0_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_0_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_0_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_0_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_0_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_0_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_0_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_0_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_0_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_0_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_0_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(mau_0_io_pipe_phv_out_valid),
    .io_mod_state_id_mod(mau_0_io_mod_state_id_mod),
    .io_mod_state_id(mau_0_io_mod_state_id),
    .io_mod_sram_w_cs(mau_0_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_0_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_0_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_0_io_mod_sram_w_data)
  );
  ParseModule mau_1 ( // @[parser_pisa.scala 31:25]
    .clock(mau_1_clock),
    .io_pipe_phv_in_data_0(mau_1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(mau_1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(mau_1_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(mau_1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(mau_1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_1_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(mau_1_io_pipe_phv_out_valid),
    .io_mod_state_id_mod(mau_1_io_mod_state_id_mod),
    .io_mod_state_id(mau_1_io_mod_state_id),
    .io_mod_sram_w_cs(mau_1_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_1_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_1_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_1_io_mod_sram_w_data)
  );
  ParseModule mau_2 ( // @[parser_pisa.scala 31:25]
    .clock(mau_2_clock),
    .io_pipe_phv_in_data_0(mau_2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(mau_2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(mau_2_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(mau_2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(mau_2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_2_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(mau_2_io_pipe_phv_out_valid),
    .io_mod_state_id_mod(mau_2_io_mod_state_id_mod),
    .io_mod_state_id(mau_2_io_mod_state_id),
    .io_mod_sram_w_cs(mau_2_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_2_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_2_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_2_io_mod_sram_w_data)
  );
  ParseModule mau_3 ( // @[parser_pisa.scala 31:25]
    .clock(mau_3_clock),
    .io_pipe_phv_in_data_0(mau_3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_3_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_3_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_3_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_3_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_3_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_3_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_3_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_3_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_3_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_3_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_3_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_3_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_3_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_3_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_3_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_3_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_3_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_3_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_3_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_3_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_3_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_3_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_3_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_3_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_3_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_3_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_3_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_3_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_3_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_3_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_3_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_3_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_3_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_3_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_3_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_3_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_3_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_3_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_3_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_3_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_3_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_3_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_3_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_3_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_3_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_3_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_3_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_3_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_3_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_3_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_3_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_3_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_3_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_3_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_3_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_3_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_3_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_3_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_3_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_3_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_3_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_3_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_3_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_3_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(mau_3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(mau_3_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(mau_3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_3_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_3_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_3_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_3_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_3_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_3_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_3_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_3_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_3_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_3_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_3_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_3_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_3_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_3_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_3_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_3_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_3_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_3_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_3_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_3_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_3_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_3_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_3_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_3_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_3_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_3_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_3_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_3_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_3_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_3_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_3_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_3_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_3_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_3_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_3_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_3_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_3_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_3_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_3_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_3_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_3_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_3_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_3_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_3_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_3_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_3_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_3_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_3_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_3_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_3_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_3_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_3_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_3_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_3_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_3_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_3_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_3_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_3_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_3_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_3_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_3_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_3_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_3_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_3_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(mau_3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_3_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(mau_3_io_pipe_phv_out_valid),
    .io_mod_state_id_mod(mau_3_io_mod_state_id_mod),
    .io_mod_state_id(mau_3_io_mod_state_id),
    .io_mod_sram_w_cs(mau_3_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_3_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_3_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_3_io_mod_sram_w_data)
  );
  ParseModule mau_4 ( // @[parser_pisa.scala 31:25]
    .clock(mau_4_clock),
    .io_pipe_phv_in_data_0(mau_4_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_4_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_4_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_4_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_4_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_4_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_4_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_4_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_4_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_4_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_4_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_4_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_4_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_4_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_4_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_4_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_4_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_4_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_4_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_4_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_4_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_4_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_4_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_4_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_4_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_4_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_4_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_4_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_4_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_4_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_4_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_4_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_4_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_4_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_4_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_4_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_4_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_4_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_4_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_4_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_4_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_4_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_4_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_4_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_4_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_4_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_4_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_4_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_4_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_4_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_4_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_4_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_4_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_4_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_4_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_4_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_4_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_4_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_4_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_4_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_4_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_4_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_4_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_4_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_4_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_4_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_4_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_4_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_4_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_4_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_4_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_4_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_4_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_4_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_4_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_4_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_4_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_4_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_4_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_4_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_4_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_4_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_4_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_4_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_4_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_4_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_4_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_4_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_4_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_4_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_4_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_4_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_4_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_4_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_4_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_4_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_4_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_4_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_4_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_4_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_4_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_4_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_4_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_4_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_4_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_4_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_4_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_4_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_4_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_4_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_4_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_4_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_4_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_4_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_4_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_4_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_4_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_4_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_4_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_4_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_4_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_4_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_4_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_4_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_4_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_4_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_4_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_4_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_4_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_4_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_4_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_4_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_4_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_4_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_4_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_4_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_4_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_4_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_4_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_4_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_4_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_4_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_4_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_4_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_4_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_4_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_4_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_4_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_4_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_4_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_4_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_4_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_4_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_4_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_4_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_4_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_4_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_4_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_4_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_4_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(mau_4_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_4_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_4_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_4_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_4_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_4_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_4_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_4_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_4_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_4_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_4_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_4_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_4_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_4_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_4_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_4_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_4_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_4_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_4_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_4_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_4_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_4_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(mau_4_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(mau_4_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_4_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_4_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_4_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_4_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_4_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_4_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_4_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_4_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_4_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_4_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_4_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_4_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_4_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_4_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_4_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_4_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_4_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_4_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_4_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_4_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_4_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_4_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_4_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_4_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_4_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_4_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_4_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_4_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_4_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_4_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_4_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_4_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_4_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_4_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_4_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_4_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_4_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_4_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_4_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_4_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_4_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_4_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_4_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_4_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_4_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_4_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_4_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_4_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_4_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_4_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_4_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_4_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_4_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_4_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_4_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_4_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_4_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_4_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_4_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_4_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_4_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_4_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_4_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_4_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_4_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_4_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_4_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_4_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_4_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_4_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_4_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_4_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_4_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_4_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_4_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_4_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_4_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_4_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_4_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_4_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_4_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_4_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_4_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_4_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_4_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_4_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_4_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_4_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_4_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_4_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_4_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_4_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_4_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_4_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_4_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_4_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_4_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_4_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_4_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_4_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_4_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_4_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_4_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_4_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_4_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_4_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_4_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_4_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_4_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_4_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_4_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_4_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_4_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_4_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_4_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_4_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_4_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_4_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_4_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_4_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_4_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_4_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_4_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_4_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_4_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_4_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_4_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_4_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_4_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_4_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_4_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_4_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_4_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_4_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_4_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_4_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_4_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_4_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_4_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_4_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_4_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_4_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_4_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_4_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_4_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_4_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_4_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_4_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_4_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_4_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_4_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_4_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_4_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_4_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_4_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_4_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_4_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_4_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_4_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(mau_4_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_4_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_4_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_4_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_4_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_4_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_4_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_4_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_4_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_4_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_4_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_4_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_4_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_4_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_4_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_4_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_4_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_4_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_4_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_4_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_4_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_4_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(mau_4_io_pipe_phv_out_valid),
    .io_mod_state_id_mod(mau_4_io_mod_state_id_mod),
    .io_mod_state_id(mau_4_io_mod_state_id),
    .io_mod_sram_w_cs(mau_4_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_4_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_4_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_4_io_mod_sram_w_data)
  );
  ParseModule mau_5 ( // @[parser_pisa.scala 31:25]
    .clock(mau_5_clock),
    .io_pipe_phv_in_data_0(mau_5_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_5_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_5_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_5_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_5_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_5_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_5_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_5_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_5_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_5_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_5_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_5_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_5_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_5_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_5_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_5_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_5_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_5_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_5_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_5_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_5_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_5_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_5_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_5_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_5_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_5_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_5_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_5_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_5_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_5_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_5_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_5_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_5_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_5_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_5_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_5_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_5_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_5_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_5_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_5_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_5_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_5_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_5_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_5_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_5_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_5_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_5_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_5_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_5_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_5_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_5_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_5_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_5_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_5_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_5_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_5_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_5_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_5_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_5_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_5_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_5_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_5_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_5_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_5_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_5_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_5_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_5_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_5_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_5_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_5_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_5_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_5_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_5_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_5_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_5_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_5_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_5_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_5_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_5_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_5_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_5_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_5_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_5_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_5_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_5_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_5_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_5_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_5_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_5_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_5_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_5_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_5_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_5_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_5_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_5_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_5_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_5_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_5_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_5_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_5_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_5_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_5_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_5_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_5_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_5_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_5_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_5_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_5_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_5_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_5_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_5_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_5_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_5_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_5_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_5_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_5_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_5_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_5_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_5_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_5_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_5_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_5_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_5_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_5_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_5_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_5_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_5_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_5_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_5_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_5_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_5_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_5_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_5_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_5_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_5_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_5_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_5_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_5_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_5_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_5_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_5_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_5_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_5_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_5_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_5_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_5_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_5_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_5_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_5_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_5_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_5_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_5_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_5_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_5_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_5_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_5_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_5_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_5_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_5_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_5_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(mau_5_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_5_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_5_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_5_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_5_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_5_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_5_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_5_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_5_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_5_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_5_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_5_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_5_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_5_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_5_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_5_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_5_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_5_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_5_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_5_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_5_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_5_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(mau_5_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(mau_5_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_5_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_5_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_5_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_5_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_5_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_5_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_5_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_5_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_5_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_5_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_5_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_5_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_5_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_5_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_5_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_5_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_5_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_5_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_5_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_5_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_5_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_5_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_5_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_5_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_5_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_5_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_5_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_5_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_5_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_5_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_5_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_5_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_5_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_5_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_5_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_5_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_5_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_5_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_5_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_5_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_5_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_5_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_5_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_5_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_5_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_5_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_5_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_5_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_5_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_5_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_5_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_5_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_5_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_5_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_5_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_5_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_5_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_5_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_5_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_5_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_5_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_5_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_5_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_5_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_5_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_5_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_5_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_5_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_5_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_5_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_5_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_5_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_5_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_5_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_5_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_5_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_5_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_5_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_5_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_5_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_5_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_5_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_5_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_5_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_5_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_5_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_5_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_5_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_5_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_5_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_5_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_5_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_5_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_5_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_5_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_5_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_5_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_5_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_5_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_5_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_5_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_5_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_5_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_5_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_5_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_5_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_5_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_5_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_5_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_5_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_5_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_5_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_5_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_5_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_5_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_5_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_5_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_5_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_5_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_5_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_5_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_5_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_5_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_5_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_5_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_5_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_5_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_5_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_5_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_5_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_5_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_5_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_5_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_5_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_5_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_5_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_5_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_5_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_5_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_5_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_5_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_5_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_5_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_5_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_5_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_5_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_5_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_5_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_5_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_5_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_5_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_5_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_5_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_5_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_5_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_5_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_5_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_5_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_5_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(mau_5_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_5_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_5_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_5_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_5_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_5_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_5_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_5_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_5_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_5_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_5_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_5_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_5_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_5_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_5_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_5_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_5_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_5_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_5_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_5_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_5_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_5_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(mau_5_io_pipe_phv_out_valid),
    .io_mod_state_id_mod(mau_5_io_mod_state_id_mod),
    .io_mod_state_id(mau_5_io_mod_state_id),
    .io_mod_sram_w_cs(mau_5_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_5_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_5_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_5_io_mod_sram_w_data)
  );
  ParseModule mau_6 ( // @[parser_pisa.scala 31:25]
    .clock(mau_6_clock),
    .io_pipe_phv_in_data_0(mau_6_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_6_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_6_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_6_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_6_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_6_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_6_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_6_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_6_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_6_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_6_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_6_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_6_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_6_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_6_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_6_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_6_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_6_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_6_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_6_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_6_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_6_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_6_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_6_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_6_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_6_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_6_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_6_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_6_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_6_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_6_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_6_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_6_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_6_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_6_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_6_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_6_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_6_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_6_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_6_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_6_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_6_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_6_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_6_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_6_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_6_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_6_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_6_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_6_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_6_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_6_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_6_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_6_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_6_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_6_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_6_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_6_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_6_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_6_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_6_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_6_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_6_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_6_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_6_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_6_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_6_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_6_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_6_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_6_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_6_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_6_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_6_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_6_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_6_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_6_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_6_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_6_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_6_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_6_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_6_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_6_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_6_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_6_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_6_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_6_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_6_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_6_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_6_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_6_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_6_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_6_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_6_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_6_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_6_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_6_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_6_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_6_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_6_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_6_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_6_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_6_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_6_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_6_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_6_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_6_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_6_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_6_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_6_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_6_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_6_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_6_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_6_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_6_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_6_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_6_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_6_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_6_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_6_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_6_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_6_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_6_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_6_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_6_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_6_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_6_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_6_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_6_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_6_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_6_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_6_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_6_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_6_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_6_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_6_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_6_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_6_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_6_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_6_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_6_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_6_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_6_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_6_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_6_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_6_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_6_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_6_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_6_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_6_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_6_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_6_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_6_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_6_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_6_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_6_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_6_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_6_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_6_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_6_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_6_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_6_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(mau_6_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_6_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_6_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_6_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_6_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_6_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_6_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_6_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_6_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_6_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_6_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_6_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_6_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_6_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_6_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_6_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_6_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_6_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_6_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_6_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_6_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_6_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(mau_6_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(mau_6_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_6_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_6_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_6_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_6_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_6_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_6_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_6_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_6_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_6_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_6_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_6_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_6_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_6_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_6_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_6_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_6_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_6_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_6_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_6_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_6_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_6_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_6_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_6_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_6_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_6_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_6_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_6_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_6_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_6_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_6_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_6_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_6_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_6_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_6_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_6_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_6_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_6_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_6_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_6_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_6_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_6_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_6_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_6_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_6_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_6_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_6_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_6_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_6_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_6_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_6_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_6_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_6_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_6_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_6_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_6_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_6_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_6_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_6_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_6_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_6_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_6_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_6_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_6_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_6_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_6_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_6_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_6_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_6_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_6_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_6_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_6_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_6_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_6_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_6_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_6_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_6_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_6_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_6_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_6_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_6_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_6_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_6_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_6_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_6_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_6_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_6_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_6_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_6_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_6_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_6_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_6_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_6_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_6_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_6_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_6_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_6_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_6_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_6_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_6_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_6_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_6_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_6_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_6_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_6_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_6_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_6_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_6_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_6_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_6_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_6_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_6_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_6_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_6_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_6_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_6_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_6_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_6_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_6_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_6_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_6_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_6_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_6_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_6_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_6_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_6_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_6_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_6_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_6_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_6_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_6_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_6_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_6_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_6_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_6_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_6_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_6_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_6_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_6_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_6_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_6_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_6_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_6_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_6_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_6_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_6_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_6_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_6_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_6_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_6_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_6_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_6_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_6_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_6_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_6_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_6_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_6_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_6_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_6_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_6_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(mau_6_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_6_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_6_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_6_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_6_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_6_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_6_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_6_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_6_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_6_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_6_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_6_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_6_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_6_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_6_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_6_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_6_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_6_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_6_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_6_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_6_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_6_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(mau_6_io_pipe_phv_out_valid),
    .io_mod_state_id_mod(mau_6_io_mod_state_id_mod),
    .io_mod_state_id(mau_6_io_mod_state_id),
    .io_mod_sram_w_cs(mau_6_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_6_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_6_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_6_io_mod_sram_w_data)
  );
  ParseModule mau_7 ( // @[parser_pisa.scala 31:25]
    .clock(mau_7_clock),
    .io_pipe_phv_in_data_0(mau_7_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_7_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_7_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_7_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_7_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_7_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_7_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_7_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_7_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_7_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_7_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_7_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_7_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_7_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_7_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_7_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_7_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_7_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_7_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_7_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_7_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_7_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_7_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_7_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_7_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_7_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_7_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_7_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_7_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_7_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_7_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_7_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_7_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_7_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_7_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_7_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_7_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_7_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_7_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_7_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_7_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_7_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_7_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_7_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_7_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_7_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_7_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_7_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_7_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_7_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_7_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_7_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_7_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_7_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_7_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_7_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_7_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_7_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_7_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_7_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_7_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_7_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_7_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_7_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_7_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_7_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_7_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_7_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_7_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_7_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_7_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_7_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_7_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_7_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_7_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_7_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_7_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_7_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_7_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_7_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_7_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_7_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_7_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_7_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_7_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_7_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_7_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_7_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_7_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_7_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_7_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_7_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_7_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_7_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_7_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_7_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_7_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_7_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_7_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_7_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_7_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_7_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_7_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_7_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_7_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_7_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_7_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_7_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_7_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_7_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_7_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_7_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_7_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_7_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_7_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_7_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_7_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_7_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_7_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_7_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_7_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_7_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_7_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_7_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_7_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_7_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_7_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_7_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_7_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_7_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_7_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_7_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_7_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_7_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_7_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_7_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_7_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_7_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_7_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_7_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_7_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_7_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_7_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_7_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_7_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_7_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_7_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_7_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_7_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_7_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_7_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_7_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_7_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_7_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_7_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_7_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_7_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_7_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_7_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_7_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(mau_7_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_7_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_7_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_7_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_7_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_7_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_7_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_7_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_7_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_7_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_7_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_7_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_7_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_7_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_7_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_7_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_7_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_7_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_7_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_7_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_7_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_7_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(mau_7_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(mau_7_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_7_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_7_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_7_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_7_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_7_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_7_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_7_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_7_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_7_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_7_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_7_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_7_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_7_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_7_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_7_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_7_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_7_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_7_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_7_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_7_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_7_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_7_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_7_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_7_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_7_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_7_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_7_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_7_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_7_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_7_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_7_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_7_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_7_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_7_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_7_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_7_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_7_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_7_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_7_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_7_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_7_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_7_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_7_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_7_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_7_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_7_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_7_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_7_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_7_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_7_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_7_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_7_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_7_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_7_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_7_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_7_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_7_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_7_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_7_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_7_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_7_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_7_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_7_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_7_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_7_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_7_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_7_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_7_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_7_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_7_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_7_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_7_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_7_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_7_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_7_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_7_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_7_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_7_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_7_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_7_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_7_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_7_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_7_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_7_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_7_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_7_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_7_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_7_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_7_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_7_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_7_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_7_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_7_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_7_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_7_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_7_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_7_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_7_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_7_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_7_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_7_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_7_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_7_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_7_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_7_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_7_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_7_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_7_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_7_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_7_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_7_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_7_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_7_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_7_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_7_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_7_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_7_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_7_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_7_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_7_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_7_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_7_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_7_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_7_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_7_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_7_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_7_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_7_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_7_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_7_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_7_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_7_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_7_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_7_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_7_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_7_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_7_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_7_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_7_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_7_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_7_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_7_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_7_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_7_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_7_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_7_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_7_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_7_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_7_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_7_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_7_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_7_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_7_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_7_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_7_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_7_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_7_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_7_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_7_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(mau_7_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_7_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_7_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_7_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_7_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_7_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_7_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_7_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_7_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_7_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_7_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_7_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_7_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_7_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_7_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_7_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_7_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_7_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_7_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_7_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_7_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_7_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(mau_7_io_pipe_phv_out_valid),
    .io_mod_state_id_mod(mau_7_io_mod_state_id_mod),
    .io_mod_state_id(mau_7_io_mod_state_id),
    .io_mod_sram_w_cs(mau_7_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_7_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_7_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_7_io_mod_sram_w_data)
  );
  assign io_pipe_phv_out_data_0 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_0 : _GEN_938; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_1 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_1 : _GEN_939; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_2 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_2 : _GEN_940; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_3 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_3 : _GEN_941; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_4 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_4 : _GEN_942; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_5 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_5 : _GEN_943; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_6 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_6 : _GEN_944; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_7 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_7 : _GEN_945; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_8 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_8 : _GEN_946; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_9 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_9 : _GEN_947; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_10 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_10 : _GEN_948; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_11 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_11 : _GEN_949; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_12 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_12 : _GEN_950; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_13 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_13 : _GEN_951; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_14 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_14 : _GEN_952; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_15 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_15 : _GEN_953; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_16 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_16 : _GEN_954; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_17 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_17 : _GEN_955; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_18 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_18 : _GEN_956; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_19 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_19 : _GEN_957; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_20 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_20 : _GEN_958; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_21 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_21 : _GEN_959; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_22 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_22 : _GEN_960; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_23 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_23 : _GEN_961; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_24 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_24 : _GEN_962; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_25 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_25 : _GEN_963; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_26 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_26 : _GEN_964; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_27 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_27 : _GEN_965; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_28 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_28 : _GEN_966; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_29 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_29 : _GEN_967; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_30 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_30 : _GEN_968; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_31 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_31 : _GEN_969; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_32 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_32 : _GEN_970; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_33 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_33 : _GEN_971; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_34 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_34 : _GEN_972; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_35 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_35 : _GEN_973; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_36 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_36 : _GEN_974; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_37 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_37 : _GEN_975; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_38 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_38 : _GEN_976; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_39 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_39 : _GEN_977; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_40 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_40 : _GEN_978; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_41 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_41 : _GEN_979; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_42 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_42 : _GEN_980; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_43 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_43 : _GEN_981; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_44 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_44 : _GEN_982; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_45 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_45 : _GEN_983; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_46 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_46 : _GEN_984; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_47 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_47 : _GEN_985; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_48 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_48 : _GEN_986; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_49 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_49 : _GEN_987; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_50 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_50 : _GEN_988; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_51 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_51 : _GEN_989; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_52 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_52 : _GEN_990; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_53 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_53 : _GEN_991; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_54 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_54 : _GEN_992; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_55 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_55 : _GEN_993; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_56 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_56 : _GEN_994; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_57 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_57 : _GEN_995; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_58 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_58 : _GEN_996; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_59 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_59 : _GEN_997; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_60 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_60 : _GEN_998; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_61 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_61 : _GEN_999; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_62 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_62 : _GEN_1000; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_63 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_63 : _GEN_1001; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_64 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_64 : _GEN_1002; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_65 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_65 : _GEN_1003; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_66 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_66 : _GEN_1004; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_67 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_67 : _GEN_1005; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_68 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_68 : _GEN_1006; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_69 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_69 : _GEN_1007; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_70 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_70 : _GEN_1008; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_71 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_71 : _GEN_1009; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_72 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_72 : _GEN_1010; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_73 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_73 : _GEN_1011; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_74 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_74 : _GEN_1012; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_75 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_75 : _GEN_1013; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_76 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_76 : _GEN_1014; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_77 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_77 : _GEN_1015; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_78 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_78 : _GEN_1016; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_79 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_79 : _GEN_1017; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_80 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_80 : _GEN_1018; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_81 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_81 : _GEN_1019; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_82 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_82 : _GEN_1020; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_83 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_83 : _GEN_1021; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_84 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_84 : _GEN_1022; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_85 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_85 : _GEN_1023; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_86 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_86 : _GEN_1024; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_87 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_87 : _GEN_1025; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_88 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_88 : _GEN_1026; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_89 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_89 : _GEN_1027; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_90 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_90 : _GEN_1028; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_91 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_91 : _GEN_1029; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_92 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_92 : _GEN_1030; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_93 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_93 : _GEN_1031; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_94 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_94 : _GEN_1032; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_95 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_95 : _GEN_1033; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_96 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_96 : _GEN_1034; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_97 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_97 : _GEN_1035; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_98 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_98 : _GEN_1036; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_99 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_99 : _GEN_1037; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_100 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_100 : _GEN_1038; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_101 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_101 : _GEN_1039; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_102 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_102 : _GEN_1040; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_103 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_103 : _GEN_1041; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_104 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_104 : _GEN_1042; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_105 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_105 : _GEN_1043; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_106 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_106 : _GEN_1044; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_107 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_107 : _GEN_1045; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_108 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_108 : _GEN_1046; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_109 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_109 : _GEN_1047; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_110 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_110 : _GEN_1048; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_111 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_111 : _GEN_1049; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_112 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_112 : _GEN_1050; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_113 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_113 : _GEN_1051; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_114 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_114 : _GEN_1052; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_115 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_115 : _GEN_1053; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_116 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_116 : _GEN_1054; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_117 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_117 : _GEN_1055; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_118 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_118 : _GEN_1056; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_119 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_119 : _GEN_1057; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_120 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_120 : _GEN_1058; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_121 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_121 : _GEN_1059; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_122 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_122 : _GEN_1060; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_123 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_123 : _GEN_1061; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_124 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_124 : _GEN_1062; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_125 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_125 : _GEN_1063; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_126 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_126 : _GEN_1064; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_127 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_127 : _GEN_1065; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_128 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_128 : _GEN_1066; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_129 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_129 : _GEN_1067; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_130 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_130 : _GEN_1068; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_131 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_131 : _GEN_1069; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_132 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_132 : _GEN_1070; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_133 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_133 : _GEN_1071; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_134 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_134 : _GEN_1072; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_135 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_135 : _GEN_1073; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_136 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_136 : _GEN_1074; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_137 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_137 : _GEN_1075; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_138 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_138 : _GEN_1076; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_139 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_139 : _GEN_1077; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_140 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_140 : _GEN_1078; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_141 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_141 : _GEN_1079; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_142 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_142 : _GEN_1080; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_143 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_143 : _GEN_1081; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_144 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_144 : _GEN_1082; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_145 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_145 : _GEN_1083; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_146 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_146 : _GEN_1084; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_147 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_147 : _GEN_1085; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_148 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_148 : _GEN_1086; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_149 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_149 : _GEN_1087; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_150 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_150 : _GEN_1088; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_151 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_151 : _GEN_1089; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_152 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_152 : _GEN_1090; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_153 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_153 : _GEN_1091; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_154 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_154 : _GEN_1092; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_155 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_155 : _GEN_1093; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_156 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_156 : _GEN_1094; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_157 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_157 : _GEN_1095; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_158 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_158 : _GEN_1096; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_data_159 = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_data_159 : _GEN_1097; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_next_processor_id = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_next_processor_id : _GEN_918; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_next_config_id = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_next_config_id : _GEN_917; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign io_pipe_phv_out_valid = 4'h7 == last_mau_id ? mau_7_io_pipe_phv_out_valid : _GEN_915; // @[parser_pisa.scala 43:45 parser_pisa.scala 44:35]
  assign mau_0_clock = clock;
  assign mau_0_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_128 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_129 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_130 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_131 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_132 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_133 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_134 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_135 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_136 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_137 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_138 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_139 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_140 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_141 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_142 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_143 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_144 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_145 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_146 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_147 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_148 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_149 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_150 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_151 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_152 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_153 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_154 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_155 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_156 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_157 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_158 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_data_159 = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_0 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_1 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_2 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_3 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_4 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_5 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_6 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_7 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_8 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_9 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_10 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_11 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_12 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_13 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_14 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_header_15 = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_parse_current_state = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_parse_current_offset = 8'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_parse_transition_field = 16'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_next_processor_id = 4'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_next_config_id = 1'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_is_valid_processor = 1'h0; // @[parser_pisa.scala 40:35]
  assign mau_0_io_pipe_phv_in_valid = 1'h1; // @[parser_pisa.scala 40:35]
  assign mau_0_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j : io_mod_module_mod_state_id_mod
    ; // @[parser_pisa.scala 51:22 parser_pisa.scala 58:40 parser_pisa.scala 47:23]
  assign mau_0_io_mod_state_id = io_mod_module_mod_state_id; // @[parser_pisa.scala 47:23]
  assign mau_0_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser_pisa.scala 47:23]
  assign mau_0_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j : io_mod_module_mod_sram_w_en; // @[parser_pisa.scala 51:22 parser_pisa.scala 57:40 parser_pisa.scala 47:23]
  assign mau_0_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser_pisa.scala 47:23]
  assign mau_0_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser_pisa.scala 47:23]
  assign mau_1_clock = clock;
  assign mau_1_io_pipe_phv_in_data_0 = mau_0_io_pipe_phv_out_data_0; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_1 = mau_0_io_pipe_phv_out_data_1; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_2 = mau_0_io_pipe_phv_out_data_2; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_3 = mau_0_io_pipe_phv_out_data_3; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_4 = mau_0_io_pipe_phv_out_data_4; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_5 = mau_0_io_pipe_phv_out_data_5; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_6 = mau_0_io_pipe_phv_out_data_6; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_7 = mau_0_io_pipe_phv_out_data_7; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_8 = mau_0_io_pipe_phv_out_data_8; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_9 = mau_0_io_pipe_phv_out_data_9; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_10 = mau_0_io_pipe_phv_out_data_10; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_11 = mau_0_io_pipe_phv_out_data_11; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_12 = mau_0_io_pipe_phv_out_data_12; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_13 = mau_0_io_pipe_phv_out_data_13; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_14 = mau_0_io_pipe_phv_out_data_14; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_15 = mau_0_io_pipe_phv_out_data_15; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_16 = mau_0_io_pipe_phv_out_data_16; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_17 = mau_0_io_pipe_phv_out_data_17; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_18 = mau_0_io_pipe_phv_out_data_18; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_19 = mau_0_io_pipe_phv_out_data_19; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_20 = mau_0_io_pipe_phv_out_data_20; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_21 = mau_0_io_pipe_phv_out_data_21; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_22 = mau_0_io_pipe_phv_out_data_22; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_23 = mau_0_io_pipe_phv_out_data_23; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_24 = mau_0_io_pipe_phv_out_data_24; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_25 = mau_0_io_pipe_phv_out_data_25; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_26 = mau_0_io_pipe_phv_out_data_26; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_27 = mau_0_io_pipe_phv_out_data_27; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_28 = mau_0_io_pipe_phv_out_data_28; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_29 = mau_0_io_pipe_phv_out_data_29; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_30 = mau_0_io_pipe_phv_out_data_30; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_31 = mau_0_io_pipe_phv_out_data_31; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_32 = mau_0_io_pipe_phv_out_data_32; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_33 = mau_0_io_pipe_phv_out_data_33; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_34 = mau_0_io_pipe_phv_out_data_34; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_35 = mau_0_io_pipe_phv_out_data_35; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_36 = mau_0_io_pipe_phv_out_data_36; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_37 = mau_0_io_pipe_phv_out_data_37; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_38 = mau_0_io_pipe_phv_out_data_38; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_39 = mau_0_io_pipe_phv_out_data_39; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_40 = mau_0_io_pipe_phv_out_data_40; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_41 = mau_0_io_pipe_phv_out_data_41; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_42 = mau_0_io_pipe_phv_out_data_42; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_43 = mau_0_io_pipe_phv_out_data_43; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_44 = mau_0_io_pipe_phv_out_data_44; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_45 = mau_0_io_pipe_phv_out_data_45; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_46 = mau_0_io_pipe_phv_out_data_46; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_47 = mau_0_io_pipe_phv_out_data_47; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_48 = mau_0_io_pipe_phv_out_data_48; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_49 = mau_0_io_pipe_phv_out_data_49; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_50 = mau_0_io_pipe_phv_out_data_50; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_51 = mau_0_io_pipe_phv_out_data_51; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_52 = mau_0_io_pipe_phv_out_data_52; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_53 = mau_0_io_pipe_phv_out_data_53; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_54 = mau_0_io_pipe_phv_out_data_54; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_55 = mau_0_io_pipe_phv_out_data_55; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_56 = mau_0_io_pipe_phv_out_data_56; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_57 = mau_0_io_pipe_phv_out_data_57; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_58 = mau_0_io_pipe_phv_out_data_58; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_59 = mau_0_io_pipe_phv_out_data_59; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_60 = mau_0_io_pipe_phv_out_data_60; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_61 = mau_0_io_pipe_phv_out_data_61; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_62 = mau_0_io_pipe_phv_out_data_62; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_63 = mau_0_io_pipe_phv_out_data_63; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_64 = mau_0_io_pipe_phv_out_data_64; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_65 = mau_0_io_pipe_phv_out_data_65; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_66 = mau_0_io_pipe_phv_out_data_66; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_67 = mau_0_io_pipe_phv_out_data_67; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_68 = mau_0_io_pipe_phv_out_data_68; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_69 = mau_0_io_pipe_phv_out_data_69; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_70 = mau_0_io_pipe_phv_out_data_70; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_71 = mau_0_io_pipe_phv_out_data_71; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_72 = mau_0_io_pipe_phv_out_data_72; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_73 = mau_0_io_pipe_phv_out_data_73; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_74 = mau_0_io_pipe_phv_out_data_74; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_75 = mau_0_io_pipe_phv_out_data_75; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_76 = mau_0_io_pipe_phv_out_data_76; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_77 = mau_0_io_pipe_phv_out_data_77; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_78 = mau_0_io_pipe_phv_out_data_78; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_79 = mau_0_io_pipe_phv_out_data_79; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_80 = mau_0_io_pipe_phv_out_data_80; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_81 = mau_0_io_pipe_phv_out_data_81; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_82 = mau_0_io_pipe_phv_out_data_82; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_83 = mau_0_io_pipe_phv_out_data_83; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_84 = mau_0_io_pipe_phv_out_data_84; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_85 = mau_0_io_pipe_phv_out_data_85; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_86 = mau_0_io_pipe_phv_out_data_86; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_87 = mau_0_io_pipe_phv_out_data_87; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_88 = mau_0_io_pipe_phv_out_data_88; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_89 = mau_0_io_pipe_phv_out_data_89; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_90 = mau_0_io_pipe_phv_out_data_90; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_91 = mau_0_io_pipe_phv_out_data_91; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_92 = mau_0_io_pipe_phv_out_data_92; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_93 = mau_0_io_pipe_phv_out_data_93; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_94 = mau_0_io_pipe_phv_out_data_94; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_95 = mau_0_io_pipe_phv_out_data_95; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_96 = mau_0_io_pipe_phv_out_data_96; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_97 = mau_0_io_pipe_phv_out_data_97; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_98 = mau_0_io_pipe_phv_out_data_98; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_99 = mau_0_io_pipe_phv_out_data_99; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_100 = mau_0_io_pipe_phv_out_data_100; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_101 = mau_0_io_pipe_phv_out_data_101; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_102 = mau_0_io_pipe_phv_out_data_102; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_103 = mau_0_io_pipe_phv_out_data_103; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_104 = mau_0_io_pipe_phv_out_data_104; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_105 = mau_0_io_pipe_phv_out_data_105; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_106 = mau_0_io_pipe_phv_out_data_106; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_107 = mau_0_io_pipe_phv_out_data_107; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_108 = mau_0_io_pipe_phv_out_data_108; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_109 = mau_0_io_pipe_phv_out_data_109; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_110 = mau_0_io_pipe_phv_out_data_110; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_111 = mau_0_io_pipe_phv_out_data_111; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_112 = mau_0_io_pipe_phv_out_data_112; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_113 = mau_0_io_pipe_phv_out_data_113; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_114 = mau_0_io_pipe_phv_out_data_114; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_115 = mau_0_io_pipe_phv_out_data_115; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_116 = mau_0_io_pipe_phv_out_data_116; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_117 = mau_0_io_pipe_phv_out_data_117; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_118 = mau_0_io_pipe_phv_out_data_118; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_119 = mau_0_io_pipe_phv_out_data_119; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_120 = mau_0_io_pipe_phv_out_data_120; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_121 = mau_0_io_pipe_phv_out_data_121; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_122 = mau_0_io_pipe_phv_out_data_122; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_123 = mau_0_io_pipe_phv_out_data_123; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_124 = mau_0_io_pipe_phv_out_data_124; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_125 = mau_0_io_pipe_phv_out_data_125; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_126 = mau_0_io_pipe_phv_out_data_126; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_127 = mau_0_io_pipe_phv_out_data_127; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_128 = mau_0_io_pipe_phv_out_data_128; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_129 = mau_0_io_pipe_phv_out_data_129; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_130 = mau_0_io_pipe_phv_out_data_130; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_131 = mau_0_io_pipe_phv_out_data_131; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_132 = mau_0_io_pipe_phv_out_data_132; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_133 = mau_0_io_pipe_phv_out_data_133; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_134 = mau_0_io_pipe_phv_out_data_134; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_135 = mau_0_io_pipe_phv_out_data_135; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_136 = mau_0_io_pipe_phv_out_data_136; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_137 = mau_0_io_pipe_phv_out_data_137; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_138 = mau_0_io_pipe_phv_out_data_138; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_139 = mau_0_io_pipe_phv_out_data_139; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_140 = mau_0_io_pipe_phv_out_data_140; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_141 = mau_0_io_pipe_phv_out_data_141; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_142 = mau_0_io_pipe_phv_out_data_142; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_143 = mau_0_io_pipe_phv_out_data_143; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_144 = mau_0_io_pipe_phv_out_data_144; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_145 = mau_0_io_pipe_phv_out_data_145; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_146 = mau_0_io_pipe_phv_out_data_146; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_147 = mau_0_io_pipe_phv_out_data_147; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_148 = mau_0_io_pipe_phv_out_data_148; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_149 = mau_0_io_pipe_phv_out_data_149; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_150 = mau_0_io_pipe_phv_out_data_150; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_151 = mau_0_io_pipe_phv_out_data_151; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_152 = mau_0_io_pipe_phv_out_data_152; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_153 = mau_0_io_pipe_phv_out_data_153; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_154 = mau_0_io_pipe_phv_out_data_154; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_155 = mau_0_io_pipe_phv_out_data_155; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_156 = mau_0_io_pipe_phv_out_data_156; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_157 = mau_0_io_pipe_phv_out_data_157; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_158 = mau_0_io_pipe_phv_out_data_158; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_data_159 = mau_0_io_pipe_phv_out_data_159; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_0 = mau_0_io_pipe_phv_out_header_0; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_1 = mau_0_io_pipe_phv_out_header_1; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_2 = mau_0_io_pipe_phv_out_header_2; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_3 = mau_0_io_pipe_phv_out_header_3; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_4 = mau_0_io_pipe_phv_out_header_4; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_5 = mau_0_io_pipe_phv_out_header_5; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_6 = mau_0_io_pipe_phv_out_header_6; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_7 = mau_0_io_pipe_phv_out_header_7; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_8 = mau_0_io_pipe_phv_out_header_8; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_9 = mau_0_io_pipe_phv_out_header_9; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_10 = mau_0_io_pipe_phv_out_header_10; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_11 = mau_0_io_pipe_phv_out_header_11; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_12 = mau_0_io_pipe_phv_out_header_12; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_13 = mau_0_io_pipe_phv_out_header_13; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_14 = mau_0_io_pipe_phv_out_header_14; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_header_15 = mau_0_io_pipe_phv_out_header_15; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_parse_current_state = mau_0_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_parse_current_offset = mau_0_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_parse_transition_field = mau_0_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_next_processor_id = mau_0_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_next_config_id = mau_0_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_is_valid_processor = mau_0_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 42:35]
  assign mau_1_io_pipe_phv_in_valid = mau_0_io_pipe_phv_out_valid; // @[parser_pisa.scala 42:35]
  assign mau_1_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_1 :
    io_mod_module_mod_state_id_mod; // @[parser_pisa.scala 51:22 parser_pisa.scala 58:40 parser_pisa.scala 47:23]
  assign mau_1_io_mod_state_id = io_mod_module_mod_state_id; // @[parser_pisa.scala 47:23]
  assign mau_1_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser_pisa.scala 47:23]
  assign mau_1_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_1 : io_mod_module_mod_sram_w_en; // @[parser_pisa.scala 51:22 parser_pisa.scala 57:40 parser_pisa.scala 47:23]
  assign mau_1_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser_pisa.scala 47:23]
  assign mau_1_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser_pisa.scala 47:23]
  assign mau_2_clock = clock;
  assign mau_2_io_pipe_phv_in_data_0 = mau_1_io_pipe_phv_out_data_0; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_1 = mau_1_io_pipe_phv_out_data_1; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_2 = mau_1_io_pipe_phv_out_data_2; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_3 = mau_1_io_pipe_phv_out_data_3; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_4 = mau_1_io_pipe_phv_out_data_4; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_5 = mau_1_io_pipe_phv_out_data_5; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_6 = mau_1_io_pipe_phv_out_data_6; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_7 = mau_1_io_pipe_phv_out_data_7; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_8 = mau_1_io_pipe_phv_out_data_8; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_9 = mau_1_io_pipe_phv_out_data_9; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_10 = mau_1_io_pipe_phv_out_data_10; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_11 = mau_1_io_pipe_phv_out_data_11; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_12 = mau_1_io_pipe_phv_out_data_12; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_13 = mau_1_io_pipe_phv_out_data_13; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_14 = mau_1_io_pipe_phv_out_data_14; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_15 = mau_1_io_pipe_phv_out_data_15; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_16 = mau_1_io_pipe_phv_out_data_16; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_17 = mau_1_io_pipe_phv_out_data_17; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_18 = mau_1_io_pipe_phv_out_data_18; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_19 = mau_1_io_pipe_phv_out_data_19; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_20 = mau_1_io_pipe_phv_out_data_20; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_21 = mau_1_io_pipe_phv_out_data_21; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_22 = mau_1_io_pipe_phv_out_data_22; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_23 = mau_1_io_pipe_phv_out_data_23; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_24 = mau_1_io_pipe_phv_out_data_24; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_25 = mau_1_io_pipe_phv_out_data_25; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_26 = mau_1_io_pipe_phv_out_data_26; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_27 = mau_1_io_pipe_phv_out_data_27; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_28 = mau_1_io_pipe_phv_out_data_28; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_29 = mau_1_io_pipe_phv_out_data_29; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_30 = mau_1_io_pipe_phv_out_data_30; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_31 = mau_1_io_pipe_phv_out_data_31; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_32 = mau_1_io_pipe_phv_out_data_32; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_33 = mau_1_io_pipe_phv_out_data_33; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_34 = mau_1_io_pipe_phv_out_data_34; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_35 = mau_1_io_pipe_phv_out_data_35; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_36 = mau_1_io_pipe_phv_out_data_36; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_37 = mau_1_io_pipe_phv_out_data_37; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_38 = mau_1_io_pipe_phv_out_data_38; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_39 = mau_1_io_pipe_phv_out_data_39; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_40 = mau_1_io_pipe_phv_out_data_40; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_41 = mau_1_io_pipe_phv_out_data_41; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_42 = mau_1_io_pipe_phv_out_data_42; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_43 = mau_1_io_pipe_phv_out_data_43; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_44 = mau_1_io_pipe_phv_out_data_44; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_45 = mau_1_io_pipe_phv_out_data_45; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_46 = mau_1_io_pipe_phv_out_data_46; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_47 = mau_1_io_pipe_phv_out_data_47; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_48 = mau_1_io_pipe_phv_out_data_48; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_49 = mau_1_io_pipe_phv_out_data_49; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_50 = mau_1_io_pipe_phv_out_data_50; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_51 = mau_1_io_pipe_phv_out_data_51; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_52 = mau_1_io_pipe_phv_out_data_52; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_53 = mau_1_io_pipe_phv_out_data_53; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_54 = mau_1_io_pipe_phv_out_data_54; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_55 = mau_1_io_pipe_phv_out_data_55; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_56 = mau_1_io_pipe_phv_out_data_56; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_57 = mau_1_io_pipe_phv_out_data_57; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_58 = mau_1_io_pipe_phv_out_data_58; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_59 = mau_1_io_pipe_phv_out_data_59; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_60 = mau_1_io_pipe_phv_out_data_60; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_61 = mau_1_io_pipe_phv_out_data_61; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_62 = mau_1_io_pipe_phv_out_data_62; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_63 = mau_1_io_pipe_phv_out_data_63; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_64 = mau_1_io_pipe_phv_out_data_64; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_65 = mau_1_io_pipe_phv_out_data_65; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_66 = mau_1_io_pipe_phv_out_data_66; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_67 = mau_1_io_pipe_phv_out_data_67; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_68 = mau_1_io_pipe_phv_out_data_68; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_69 = mau_1_io_pipe_phv_out_data_69; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_70 = mau_1_io_pipe_phv_out_data_70; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_71 = mau_1_io_pipe_phv_out_data_71; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_72 = mau_1_io_pipe_phv_out_data_72; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_73 = mau_1_io_pipe_phv_out_data_73; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_74 = mau_1_io_pipe_phv_out_data_74; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_75 = mau_1_io_pipe_phv_out_data_75; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_76 = mau_1_io_pipe_phv_out_data_76; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_77 = mau_1_io_pipe_phv_out_data_77; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_78 = mau_1_io_pipe_phv_out_data_78; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_79 = mau_1_io_pipe_phv_out_data_79; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_80 = mau_1_io_pipe_phv_out_data_80; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_81 = mau_1_io_pipe_phv_out_data_81; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_82 = mau_1_io_pipe_phv_out_data_82; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_83 = mau_1_io_pipe_phv_out_data_83; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_84 = mau_1_io_pipe_phv_out_data_84; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_85 = mau_1_io_pipe_phv_out_data_85; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_86 = mau_1_io_pipe_phv_out_data_86; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_87 = mau_1_io_pipe_phv_out_data_87; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_88 = mau_1_io_pipe_phv_out_data_88; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_89 = mau_1_io_pipe_phv_out_data_89; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_90 = mau_1_io_pipe_phv_out_data_90; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_91 = mau_1_io_pipe_phv_out_data_91; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_92 = mau_1_io_pipe_phv_out_data_92; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_93 = mau_1_io_pipe_phv_out_data_93; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_94 = mau_1_io_pipe_phv_out_data_94; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_95 = mau_1_io_pipe_phv_out_data_95; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_96 = mau_1_io_pipe_phv_out_data_96; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_97 = mau_1_io_pipe_phv_out_data_97; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_98 = mau_1_io_pipe_phv_out_data_98; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_99 = mau_1_io_pipe_phv_out_data_99; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_100 = mau_1_io_pipe_phv_out_data_100; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_101 = mau_1_io_pipe_phv_out_data_101; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_102 = mau_1_io_pipe_phv_out_data_102; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_103 = mau_1_io_pipe_phv_out_data_103; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_104 = mau_1_io_pipe_phv_out_data_104; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_105 = mau_1_io_pipe_phv_out_data_105; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_106 = mau_1_io_pipe_phv_out_data_106; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_107 = mau_1_io_pipe_phv_out_data_107; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_108 = mau_1_io_pipe_phv_out_data_108; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_109 = mau_1_io_pipe_phv_out_data_109; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_110 = mau_1_io_pipe_phv_out_data_110; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_111 = mau_1_io_pipe_phv_out_data_111; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_112 = mau_1_io_pipe_phv_out_data_112; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_113 = mau_1_io_pipe_phv_out_data_113; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_114 = mau_1_io_pipe_phv_out_data_114; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_115 = mau_1_io_pipe_phv_out_data_115; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_116 = mau_1_io_pipe_phv_out_data_116; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_117 = mau_1_io_pipe_phv_out_data_117; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_118 = mau_1_io_pipe_phv_out_data_118; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_119 = mau_1_io_pipe_phv_out_data_119; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_120 = mau_1_io_pipe_phv_out_data_120; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_121 = mau_1_io_pipe_phv_out_data_121; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_122 = mau_1_io_pipe_phv_out_data_122; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_123 = mau_1_io_pipe_phv_out_data_123; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_124 = mau_1_io_pipe_phv_out_data_124; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_125 = mau_1_io_pipe_phv_out_data_125; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_126 = mau_1_io_pipe_phv_out_data_126; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_127 = mau_1_io_pipe_phv_out_data_127; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_128 = mau_1_io_pipe_phv_out_data_128; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_129 = mau_1_io_pipe_phv_out_data_129; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_130 = mau_1_io_pipe_phv_out_data_130; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_131 = mau_1_io_pipe_phv_out_data_131; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_132 = mau_1_io_pipe_phv_out_data_132; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_133 = mau_1_io_pipe_phv_out_data_133; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_134 = mau_1_io_pipe_phv_out_data_134; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_135 = mau_1_io_pipe_phv_out_data_135; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_136 = mau_1_io_pipe_phv_out_data_136; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_137 = mau_1_io_pipe_phv_out_data_137; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_138 = mau_1_io_pipe_phv_out_data_138; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_139 = mau_1_io_pipe_phv_out_data_139; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_140 = mau_1_io_pipe_phv_out_data_140; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_141 = mau_1_io_pipe_phv_out_data_141; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_142 = mau_1_io_pipe_phv_out_data_142; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_143 = mau_1_io_pipe_phv_out_data_143; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_144 = mau_1_io_pipe_phv_out_data_144; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_145 = mau_1_io_pipe_phv_out_data_145; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_146 = mau_1_io_pipe_phv_out_data_146; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_147 = mau_1_io_pipe_phv_out_data_147; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_148 = mau_1_io_pipe_phv_out_data_148; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_149 = mau_1_io_pipe_phv_out_data_149; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_150 = mau_1_io_pipe_phv_out_data_150; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_151 = mau_1_io_pipe_phv_out_data_151; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_152 = mau_1_io_pipe_phv_out_data_152; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_153 = mau_1_io_pipe_phv_out_data_153; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_154 = mau_1_io_pipe_phv_out_data_154; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_155 = mau_1_io_pipe_phv_out_data_155; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_156 = mau_1_io_pipe_phv_out_data_156; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_157 = mau_1_io_pipe_phv_out_data_157; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_158 = mau_1_io_pipe_phv_out_data_158; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_data_159 = mau_1_io_pipe_phv_out_data_159; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_0 = mau_1_io_pipe_phv_out_header_0; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_1 = mau_1_io_pipe_phv_out_header_1; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_2 = mau_1_io_pipe_phv_out_header_2; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_3 = mau_1_io_pipe_phv_out_header_3; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_4 = mau_1_io_pipe_phv_out_header_4; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_5 = mau_1_io_pipe_phv_out_header_5; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_6 = mau_1_io_pipe_phv_out_header_6; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_7 = mau_1_io_pipe_phv_out_header_7; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_8 = mau_1_io_pipe_phv_out_header_8; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_9 = mau_1_io_pipe_phv_out_header_9; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_10 = mau_1_io_pipe_phv_out_header_10; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_11 = mau_1_io_pipe_phv_out_header_11; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_12 = mau_1_io_pipe_phv_out_header_12; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_13 = mau_1_io_pipe_phv_out_header_13; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_14 = mau_1_io_pipe_phv_out_header_14; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_header_15 = mau_1_io_pipe_phv_out_header_15; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_parse_current_state = mau_1_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_parse_current_offset = mau_1_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_parse_transition_field = mau_1_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_next_processor_id = mau_1_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_next_config_id = mau_1_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_is_valid_processor = mau_1_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 42:35]
  assign mau_2_io_pipe_phv_in_valid = mau_1_io_pipe_phv_out_valid; // @[parser_pisa.scala 42:35]
  assign mau_2_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_2 :
    io_mod_module_mod_state_id_mod; // @[parser_pisa.scala 51:22 parser_pisa.scala 58:40 parser_pisa.scala 47:23]
  assign mau_2_io_mod_state_id = io_mod_module_mod_state_id; // @[parser_pisa.scala 47:23]
  assign mau_2_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser_pisa.scala 47:23]
  assign mau_2_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_2 : io_mod_module_mod_sram_w_en; // @[parser_pisa.scala 51:22 parser_pisa.scala 57:40 parser_pisa.scala 47:23]
  assign mau_2_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser_pisa.scala 47:23]
  assign mau_2_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser_pisa.scala 47:23]
  assign mau_3_clock = clock;
  assign mau_3_io_pipe_phv_in_data_0 = mau_2_io_pipe_phv_out_data_0; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_1 = mau_2_io_pipe_phv_out_data_1; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_2 = mau_2_io_pipe_phv_out_data_2; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_3 = mau_2_io_pipe_phv_out_data_3; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_4 = mau_2_io_pipe_phv_out_data_4; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_5 = mau_2_io_pipe_phv_out_data_5; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_6 = mau_2_io_pipe_phv_out_data_6; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_7 = mau_2_io_pipe_phv_out_data_7; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_8 = mau_2_io_pipe_phv_out_data_8; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_9 = mau_2_io_pipe_phv_out_data_9; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_10 = mau_2_io_pipe_phv_out_data_10; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_11 = mau_2_io_pipe_phv_out_data_11; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_12 = mau_2_io_pipe_phv_out_data_12; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_13 = mau_2_io_pipe_phv_out_data_13; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_14 = mau_2_io_pipe_phv_out_data_14; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_15 = mau_2_io_pipe_phv_out_data_15; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_16 = mau_2_io_pipe_phv_out_data_16; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_17 = mau_2_io_pipe_phv_out_data_17; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_18 = mau_2_io_pipe_phv_out_data_18; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_19 = mau_2_io_pipe_phv_out_data_19; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_20 = mau_2_io_pipe_phv_out_data_20; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_21 = mau_2_io_pipe_phv_out_data_21; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_22 = mau_2_io_pipe_phv_out_data_22; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_23 = mau_2_io_pipe_phv_out_data_23; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_24 = mau_2_io_pipe_phv_out_data_24; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_25 = mau_2_io_pipe_phv_out_data_25; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_26 = mau_2_io_pipe_phv_out_data_26; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_27 = mau_2_io_pipe_phv_out_data_27; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_28 = mau_2_io_pipe_phv_out_data_28; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_29 = mau_2_io_pipe_phv_out_data_29; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_30 = mau_2_io_pipe_phv_out_data_30; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_31 = mau_2_io_pipe_phv_out_data_31; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_32 = mau_2_io_pipe_phv_out_data_32; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_33 = mau_2_io_pipe_phv_out_data_33; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_34 = mau_2_io_pipe_phv_out_data_34; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_35 = mau_2_io_pipe_phv_out_data_35; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_36 = mau_2_io_pipe_phv_out_data_36; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_37 = mau_2_io_pipe_phv_out_data_37; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_38 = mau_2_io_pipe_phv_out_data_38; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_39 = mau_2_io_pipe_phv_out_data_39; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_40 = mau_2_io_pipe_phv_out_data_40; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_41 = mau_2_io_pipe_phv_out_data_41; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_42 = mau_2_io_pipe_phv_out_data_42; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_43 = mau_2_io_pipe_phv_out_data_43; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_44 = mau_2_io_pipe_phv_out_data_44; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_45 = mau_2_io_pipe_phv_out_data_45; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_46 = mau_2_io_pipe_phv_out_data_46; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_47 = mau_2_io_pipe_phv_out_data_47; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_48 = mau_2_io_pipe_phv_out_data_48; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_49 = mau_2_io_pipe_phv_out_data_49; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_50 = mau_2_io_pipe_phv_out_data_50; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_51 = mau_2_io_pipe_phv_out_data_51; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_52 = mau_2_io_pipe_phv_out_data_52; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_53 = mau_2_io_pipe_phv_out_data_53; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_54 = mau_2_io_pipe_phv_out_data_54; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_55 = mau_2_io_pipe_phv_out_data_55; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_56 = mau_2_io_pipe_phv_out_data_56; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_57 = mau_2_io_pipe_phv_out_data_57; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_58 = mau_2_io_pipe_phv_out_data_58; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_59 = mau_2_io_pipe_phv_out_data_59; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_60 = mau_2_io_pipe_phv_out_data_60; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_61 = mau_2_io_pipe_phv_out_data_61; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_62 = mau_2_io_pipe_phv_out_data_62; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_63 = mau_2_io_pipe_phv_out_data_63; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_64 = mau_2_io_pipe_phv_out_data_64; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_65 = mau_2_io_pipe_phv_out_data_65; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_66 = mau_2_io_pipe_phv_out_data_66; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_67 = mau_2_io_pipe_phv_out_data_67; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_68 = mau_2_io_pipe_phv_out_data_68; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_69 = mau_2_io_pipe_phv_out_data_69; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_70 = mau_2_io_pipe_phv_out_data_70; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_71 = mau_2_io_pipe_phv_out_data_71; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_72 = mau_2_io_pipe_phv_out_data_72; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_73 = mau_2_io_pipe_phv_out_data_73; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_74 = mau_2_io_pipe_phv_out_data_74; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_75 = mau_2_io_pipe_phv_out_data_75; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_76 = mau_2_io_pipe_phv_out_data_76; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_77 = mau_2_io_pipe_phv_out_data_77; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_78 = mau_2_io_pipe_phv_out_data_78; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_79 = mau_2_io_pipe_phv_out_data_79; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_80 = mau_2_io_pipe_phv_out_data_80; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_81 = mau_2_io_pipe_phv_out_data_81; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_82 = mau_2_io_pipe_phv_out_data_82; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_83 = mau_2_io_pipe_phv_out_data_83; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_84 = mau_2_io_pipe_phv_out_data_84; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_85 = mau_2_io_pipe_phv_out_data_85; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_86 = mau_2_io_pipe_phv_out_data_86; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_87 = mau_2_io_pipe_phv_out_data_87; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_88 = mau_2_io_pipe_phv_out_data_88; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_89 = mau_2_io_pipe_phv_out_data_89; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_90 = mau_2_io_pipe_phv_out_data_90; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_91 = mau_2_io_pipe_phv_out_data_91; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_92 = mau_2_io_pipe_phv_out_data_92; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_93 = mau_2_io_pipe_phv_out_data_93; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_94 = mau_2_io_pipe_phv_out_data_94; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_95 = mau_2_io_pipe_phv_out_data_95; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_96 = mau_2_io_pipe_phv_out_data_96; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_97 = mau_2_io_pipe_phv_out_data_97; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_98 = mau_2_io_pipe_phv_out_data_98; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_99 = mau_2_io_pipe_phv_out_data_99; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_100 = mau_2_io_pipe_phv_out_data_100; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_101 = mau_2_io_pipe_phv_out_data_101; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_102 = mau_2_io_pipe_phv_out_data_102; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_103 = mau_2_io_pipe_phv_out_data_103; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_104 = mau_2_io_pipe_phv_out_data_104; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_105 = mau_2_io_pipe_phv_out_data_105; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_106 = mau_2_io_pipe_phv_out_data_106; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_107 = mau_2_io_pipe_phv_out_data_107; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_108 = mau_2_io_pipe_phv_out_data_108; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_109 = mau_2_io_pipe_phv_out_data_109; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_110 = mau_2_io_pipe_phv_out_data_110; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_111 = mau_2_io_pipe_phv_out_data_111; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_112 = mau_2_io_pipe_phv_out_data_112; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_113 = mau_2_io_pipe_phv_out_data_113; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_114 = mau_2_io_pipe_phv_out_data_114; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_115 = mau_2_io_pipe_phv_out_data_115; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_116 = mau_2_io_pipe_phv_out_data_116; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_117 = mau_2_io_pipe_phv_out_data_117; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_118 = mau_2_io_pipe_phv_out_data_118; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_119 = mau_2_io_pipe_phv_out_data_119; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_120 = mau_2_io_pipe_phv_out_data_120; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_121 = mau_2_io_pipe_phv_out_data_121; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_122 = mau_2_io_pipe_phv_out_data_122; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_123 = mau_2_io_pipe_phv_out_data_123; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_124 = mau_2_io_pipe_phv_out_data_124; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_125 = mau_2_io_pipe_phv_out_data_125; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_126 = mau_2_io_pipe_phv_out_data_126; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_127 = mau_2_io_pipe_phv_out_data_127; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_128 = mau_2_io_pipe_phv_out_data_128; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_129 = mau_2_io_pipe_phv_out_data_129; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_130 = mau_2_io_pipe_phv_out_data_130; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_131 = mau_2_io_pipe_phv_out_data_131; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_132 = mau_2_io_pipe_phv_out_data_132; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_133 = mau_2_io_pipe_phv_out_data_133; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_134 = mau_2_io_pipe_phv_out_data_134; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_135 = mau_2_io_pipe_phv_out_data_135; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_136 = mau_2_io_pipe_phv_out_data_136; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_137 = mau_2_io_pipe_phv_out_data_137; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_138 = mau_2_io_pipe_phv_out_data_138; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_139 = mau_2_io_pipe_phv_out_data_139; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_140 = mau_2_io_pipe_phv_out_data_140; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_141 = mau_2_io_pipe_phv_out_data_141; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_142 = mau_2_io_pipe_phv_out_data_142; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_143 = mau_2_io_pipe_phv_out_data_143; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_144 = mau_2_io_pipe_phv_out_data_144; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_145 = mau_2_io_pipe_phv_out_data_145; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_146 = mau_2_io_pipe_phv_out_data_146; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_147 = mau_2_io_pipe_phv_out_data_147; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_148 = mau_2_io_pipe_phv_out_data_148; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_149 = mau_2_io_pipe_phv_out_data_149; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_150 = mau_2_io_pipe_phv_out_data_150; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_151 = mau_2_io_pipe_phv_out_data_151; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_152 = mau_2_io_pipe_phv_out_data_152; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_153 = mau_2_io_pipe_phv_out_data_153; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_154 = mau_2_io_pipe_phv_out_data_154; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_155 = mau_2_io_pipe_phv_out_data_155; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_156 = mau_2_io_pipe_phv_out_data_156; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_157 = mau_2_io_pipe_phv_out_data_157; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_158 = mau_2_io_pipe_phv_out_data_158; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_data_159 = mau_2_io_pipe_phv_out_data_159; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_0 = mau_2_io_pipe_phv_out_header_0; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_1 = mau_2_io_pipe_phv_out_header_1; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_2 = mau_2_io_pipe_phv_out_header_2; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_3 = mau_2_io_pipe_phv_out_header_3; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_4 = mau_2_io_pipe_phv_out_header_4; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_5 = mau_2_io_pipe_phv_out_header_5; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_6 = mau_2_io_pipe_phv_out_header_6; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_7 = mau_2_io_pipe_phv_out_header_7; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_8 = mau_2_io_pipe_phv_out_header_8; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_9 = mau_2_io_pipe_phv_out_header_9; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_10 = mau_2_io_pipe_phv_out_header_10; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_11 = mau_2_io_pipe_phv_out_header_11; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_12 = mau_2_io_pipe_phv_out_header_12; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_13 = mau_2_io_pipe_phv_out_header_13; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_14 = mau_2_io_pipe_phv_out_header_14; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_header_15 = mau_2_io_pipe_phv_out_header_15; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_parse_current_state = mau_2_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_parse_current_offset = mau_2_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_parse_transition_field = mau_2_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_next_processor_id = mau_2_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_next_config_id = mau_2_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_is_valid_processor = mau_2_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 42:35]
  assign mau_3_io_pipe_phv_in_valid = mau_2_io_pipe_phv_out_valid; // @[parser_pisa.scala 42:35]
  assign mau_3_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_3 :
    io_mod_module_mod_state_id_mod; // @[parser_pisa.scala 51:22 parser_pisa.scala 58:40 parser_pisa.scala 47:23]
  assign mau_3_io_mod_state_id = io_mod_module_mod_state_id; // @[parser_pisa.scala 47:23]
  assign mau_3_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser_pisa.scala 47:23]
  assign mau_3_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_3 : io_mod_module_mod_sram_w_en; // @[parser_pisa.scala 51:22 parser_pisa.scala 57:40 parser_pisa.scala 47:23]
  assign mau_3_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser_pisa.scala 47:23]
  assign mau_3_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser_pisa.scala 47:23]
  assign mau_4_clock = clock;
  assign mau_4_io_pipe_phv_in_data_0 = mau_3_io_pipe_phv_out_data_0; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_1 = mau_3_io_pipe_phv_out_data_1; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_2 = mau_3_io_pipe_phv_out_data_2; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_3 = mau_3_io_pipe_phv_out_data_3; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_4 = mau_3_io_pipe_phv_out_data_4; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_5 = mau_3_io_pipe_phv_out_data_5; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_6 = mau_3_io_pipe_phv_out_data_6; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_7 = mau_3_io_pipe_phv_out_data_7; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_8 = mau_3_io_pipe_phv_out_data_8; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_9 = mau_3_io_pipe_phv_out_data_9; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_10 = mau_3_io_pipe_phv_out_data_10; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_11 = mau_3_io_pipe_phv_out_data_11; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_12 = mau_3_io_pipe_phv_out_data_12; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_13 = mau_3_io_pipe_phv_out_data_13; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_14 = mau_3_io_pipe_phv_out_data_14; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_15 = mau_3_io_pipe_phv_out_data_15; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_16 = mau_3_io_pipe_phv_out_data_16; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_17 = mau_3_io_pipe_phv_out_data_17; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_18 = mau_3_io_pipe_phv_out_data_18; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_19 = mau_3_io_pipe_phv_out_data_19; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_20 = mau_3_io_pipe_phv_out_data_20; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_21 = mau_3_io_pipe_phv_out_data_21; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_22 = mau_3_io_pipe_phv_out_data_22; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_23 = mau_3_io_pipe_phv_out_data_23; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_24 = mau_3_io_pipe_phv_out_data_24; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_25 = mau_3_io_pipe_phv_out_data_25; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_26 = mau_3_io_pipe_phv_out_data_26; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_27 = mau_3_io_pipe_phv_out_data_27; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_28 = mau_3_io_pipe_phv_out_data_28; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_29 = mau_3_io_pipe_phv_out_data_29; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_30 = mau_3_io_pipe_phv_out_data_30; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_31 = mau_3_io_pipe_phv_out_data_31; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_32 = mau_3_io_pipe_phv_out_data_32; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_33 = mau_3_io_pipe_phv_out_data_33; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_34 = mau_3_io_pipe_phv_out_data_34; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_35 = mau_3_io_pipe_phv_out_data_35; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_36 = mau_3_io_pipe_phv_out_data_36; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_37 = mau_3_io_pipe_phv_out_data_37; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_38 = mau_3_io_pipe_phv_out_data_38; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_39 = mau_3_io_pipe_phv_out_data_39; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_40 = mau_3_io_pipe_phv_out_data_40; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_41 = mau_3_io_pipe_phv_out_data_41; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_42 = mau_3_io_pipe_phv_out_data_42; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_43 = mau_3_io_pipe_phv_out_data_43; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_44 = mau_3_io_pipe_phv_out_data_44; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_45 = mau_3_io_pipe_phv_out_data_45; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_46 = mau_3_io_pipe_phv_out_data_46; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_47 = mau_3_io_pipe_phv_out_data_47; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_48 = mau_3_io_pipe_phv_out_data_48; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_49 = mau_3_io_pipe_phv_out_data_49; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_50 = mau_3_io_pipe_phv_out_data_50; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_51 = mau_3_io_pipe_phv_out_data_51; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_52 = mau_3_io_pipe_phv_out_data_52; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_53 = mau_3_io_pipe_phv_out_data_53; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_54 = mau_3_io_pipe_phv_out_data_54; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_55 = mau_3_io_pipe_phv_out_data_55; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_56 = mau_3_io_pipe_phv_out_data_56; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_57 = mau_3_io_pipe_phv_out_data_57; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_58 = mau_3_io_pipe_phv_out_data_58; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_59 = mau_3_io_pipe_phv_out_data_59; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_60 = mau_3_io_pipe_phv_out_data_60; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_61 = mau_3_io_pipe_phv_out_data_61; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_62 = mau_3_io_pipe_phv_out_data_62; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_63 = mau_3_io_pipe_phv_out_data_63; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_64 = mau_3_io_pipe_phv_out_data_64; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_65 = mau_3_io_pipe_phv_out_data_65; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_66 = mau_3_io_pipe_phv_out_data_66; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_67 = mau_3_io_pipe_phv_out_data_67; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_68 = mau_3_io_pipe_phv_out_data_68; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_69 = mau_3_io_pipe_phv_out_data_69; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_70 = mau_3_io_pipe_phv_out_data_70; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_71 = mau_3_io_pipe_phv_out_data_71; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_72 = mau_3_io_pipe_phv_out_data_72; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_73 = mau_3_io_pipe_phv_out_data_73; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_74 = mau_3_io_pipe_phv_out_data_74; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_75 = mau_3_io_pipe_phv_out_data_75; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_76 = mau_3_io_pipe_phv_out_data_76; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_77 = mau_3_io_pipe_phv_out_data_77; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_78 = mau_3_io_pipe_phv_out_data_78; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_79 = mau_3_io_pipe_phv_out_data_79; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_80 = mau_3_io_pipe_phv_out_data_80; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_81 = mau_3_io_pipe_phv_out_data_81; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_82 = mau_3_io_pipe_phv_out_data_82; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_83 = mau_3_io_pipe_phv_out_data_83; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_84 = mau_3_io_pipe_phv_out_data_84; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_85 = mau_3_io_pipe_phv_out_data_85; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_86 = mau_3_io_pipe_phv_out_data_86; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_87 = mau_3_io_pipe_phv_out_data_87; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_88 = mau_3_io_pipe_phv_out_data_88; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_89 = mau_3_io_pipe_phv_out_data_89; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_90 = mau_3_io_pipe_phv_out_data_90; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_91 = mau_3_io_pipe_phv_out_data_91; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_92 = mau_3_io_pipe_phv_out_data_92; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_93 = mau_3_io_pipe_phv_out_data_93; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_94 = mau_3_io_pipe_phv_out_data_94; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_95 = mau_3_io_pipe_phv_out_data_95; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_96 = mau_3_io_pipe_phv_out_data_96; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_97 = mau_3_io_pipe_phv_out_data_97; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_98 = mau_3_io_pipe_phv_out_data_98; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_99 = mau_3_io_pipe_phv_out_data_99; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_100 = mau_3_io_pipe_phv_out_data_100; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_101 = mau_3_io_pipe_phv_out_data_101; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_102 = mau_3_io_pipe_phv_out_data_102; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_103 = mau_3_io_pipe_phv_out_data_103; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_104 = mau_3_io_pipe_phv_out_data_104; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_105 = mau_3_io_pipe_phv_out_data_105; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_106 = mau_3_io_pipe_phv_out_data_106; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_107 = mau_3_io_pipe_phv_out_data_107; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_108 = mau_3_io_pipe_phv_out_data_108; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_109 = mau_3_io_pipe_phv_out_data_109; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_110 = mau_3_io_pipe_phv_out_data_110; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_111 = mau_3_io_pipe_phv_out_data_111; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_112 = mau_3_io_pipe_phv_out_data_112; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_113 = mau_3_io_pipe_phv_out_data_113; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_114 = mau_3_io_pipe_phv_out_data_114; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_115 = mau_3_io_pipe_phv_out_data_115; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_116 = mau_3_io_pipe_phv_out_data_116; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_117 = mau_3_io_pipe_phv_out_data_117; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_118 = mau_3_io_pipe_phv_out_data_118; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_119 = mau_3_io_pipe_phv_out_data_119; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_120 = mau_3_io_pipe_phv_out_data_120; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_121 = mau_3_io_pipe_phv_out_data_121; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_122 = mau_3_io_pipe_phv_out_data_122; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_123 = mau_3_io_pipe_phv_out_data_123; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_124 = mau_3_io_pipe_phv_out_data_124; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_125 = mau_3_io_pipe_phv_out_data_125; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_126 = mau_3_io_pipe_phv_out_data_126; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_127 = mau_3_io_pipe_phv_out_data_127; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_128 = mau_3_io_pipe_phv_out_data_128; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_129 = mau_3_io_pipe_phv_out_data_129; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_130 = mau_3_io_pipe_phv_out_data_130; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_131 = mau_3_io_pipe_phv_out_data_131; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_132 = mau_3_io_pipe_phv_out_data_132; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_133 = mau_3_io_pipe_phv_out_data_133; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_134 = mau_3_io_pipe_phv_out_data_134; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_135 = mau_3_io_pipe_phv_out_data_135; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_136 = mau_3_io_pipe_phv_out_data_136; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_137 = mau_3_io_pipe_phv_out_data_137; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_138 = mau_3_io_pipe_phv_out_data_138; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_139 = mau_3_io_pipe_phv_out_data_139; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_140 = mau_3_io_pipe_phv_out_data_140; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_141 = mau_3_io_pipe_phv_out_data_141; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_142 = mau_3_io_pipe_phv_out_data_142; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_143 = mau_3_io_pipe_phv_out_data_143; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_144 = mau_3_io_pipe_phv_out_data_144; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_145 = mau_3_io_pipe_phv_out_data_145; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_146 = mau_3_io_pipe_phv_out_data_146; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_147 = mau_3_io_pipe_phv_out_data_147; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_148 = mau_3_io_pipe_phv_out_data_148; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_149 = mau_3_io_pipe_phv_out_data_149; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_150 = mau_3_io_pipe_phv_out_data_150; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_151 = mau_3_io_pipe_phv_out_data_151; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_152 = mau_3_io_pipe_phv_out_data_152; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_153 = mau_3_io_pipe_phv_out_data_153; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_154 = mau_3_io_pipe_phv_out_data_154; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_155 = mau_3_io_pipe_phv_out_data_155; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_156 = mau_3_io_pipe_phv_out_data_156; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_157 = mau_3_io_pipe_phv_out_data_157; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_158 = mau_3_io_pipe_phv_out_data_158; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_data_159 = mau_3_io_pipe_phv_out_data_159; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_0 = mau_3_io_pipe_phv_out_header_0; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_1 = mau_3_io_pipe_phv_out_header_1; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_2 = mau_3_io_pipe_phv_out_header_2; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_3 = mau_3_io_pipe_phv_out_header_3; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_4 = mau_3_io_pipe_phv_out_header_4; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_5 = mau_3_io_pipe_phv_out_header_5; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_6 = mau_3_io_pipe_phv_out_header_6; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_7 = mau_3_io_pipe_phv_out_header_7; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_8 = mau_3_io_pipe_phv_out_header_8; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_9 = mau_3_io_pipe_phv_out_header_9; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_10 = mau_3_io_pipe_phv_out_header_10; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_11 = mau_3_io_pipe_phv_out_header_11; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_12 = mau_3_io_pipe_phv_out_header_12; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_13 = mau_3_io_pipe_phv_out_header_13; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_14 = mau_3_io_pipe_phv_out_header_14; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_header_15 = mau_3_io_pipe_phv_out_header_15; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_parse_current_state = mau_3_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_parse_current_offset = mau_3_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_parse_transition_field = mau_3_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_next_processor_id = mau_3_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_next_config_id = mau_3_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_is_valid_processor = mau_3_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 42:35]
  assign mau_4_io_pipe_phv_in_valid = mau_3_io_pipe_phv_out_valid; // @[parser_pisa.scala 42:35]
  assign mau_4_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_4 :
    io_mod_module_mod_state_id_mod; // @[parser_pisa.scala 51:22 parser_pisa.scala 58:40 parser_pisa.scala 47:23]
  assign mau_4_io_mod_state_id = io_mod_module_mod_state_id; // @[parser_pisa.scala 47:23]
  assign mau_4_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser_pisa.scala 47:23]
  assign mau_4_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_4 : io_mod_module_mod_sram_w_en; // @[parser_pisa.scala 51:22 parser_pisa.scala 57:40 parser_pisa.scala 47:23]
  assign mau_4_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser_pisa.scala 47:23]
  assign mau_4_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser_pisa.scala 47:23]
  assign mau_5_clock = clock;
  assign mau_5_io_pipe_phv_in_data_0 = mau_4_io_pipe_phv_out_data_0; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_1 = mau_4_io_pipe_phv_out_data_1; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_2 = mau_4_io_pipe_phv_out_data_2; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_3 = mau_4_io_pipe_phv_out_data_3; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_4 = mau_4_io_pipe_phv_out_data_4; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_5 = mau_4_io_pipe_phv_out_data_5; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_6 = mau_4_io_pipe_phv_out_data_6; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_7 = mau_4_io_pipe_phv_out_data_7; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_8 = mau_4_io_pipe_phv_out_data_8; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_9 = mau_4_io_pipe_phv_out_data_9; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_10 = mau_4_io_pipe_phv_out_data_10; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_11 = mau_4_io_pipe_phv_out_data_11; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_12 = mau_4_io_pipe_phv_out_data_12; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_13 = mau_4_io_pipe_phv_out_data_13; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_14 = mau_4_io_pipe_phv_out_data_14; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_15 = mau_4_io_pipe_phv_out_data_15; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_16 = mau_4_io_pipe_phv_out_data_16; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_17 = mau_4_io_pipe_phv_out_data_17; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_18 = mau_4_io_pipe_phv_out_data_18; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_19 = mau_4_io_pipe_phv_out_data_19; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_20 = mau_4_io_pipe_phv_out_data_20; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_21 = mau_4_io_pipe_phv_out_data_21; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_22 = mau_4_io_pipe_phv_out_data_22; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_23 = mau_4_io_pipe_phv_out_data_23; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_24 = mau_4_io_pipe_phv_out_data_24; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_25 = mau_4_io_pipe_phv_out_data_25; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_26 = mau_4_io_pipe_phv_out_data_26; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_27 = mau_4_io_pipe_phv_out_data_27; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_28 = mau_4_io_pipe_phv_out_data_28; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_29 = mau_4_io_pipe_phv_out_data_29; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_30 = mau_4_io_pipe_phv_out_data_30; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_31 = mau_4_io_pipe_phv_out_data_31; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_32 = mau_4_io_pipe_phv_out_data_32; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_33 = mau_4_io_pipe_phv_out_data_33; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_34 = mau_4_io_pipe_phv_out_data_34; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_35 = mau_4_io_pipe_phv_out_data_35; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_36 = mau_4_io_pipe_phv_out_data_36; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_37 = mau_4_io_pipe_phv_out_data_37; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_38 = mau_4_io_pipe_phv_out_data_38; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_39 = mau_4_io_pipe_phv_out_data_39; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_40 = mau_4_io_pipe_phv_out_data_40; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_41 = mau_4_io_pipe_phv_out_data_41; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_42 = mau_4_io_pipe_phv_out_data_42; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_43 = mau_4_io_pipe_phv_out_data_43; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_44 = mau_4_io_pipe_phv_out_data_44; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_45 = mau_4_io_pipe_phv_out_data_45; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_46 = mau_4_io_pipe_phv_out_data_46; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_47 = mau_4_io_pipe_phv_out_data_47; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_48 = mau_4_io_pipe_phv_out_data_48; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_49 = mau_4_io_pipe_phv_out_data_49; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_50 = mau_4_io_pipe_phv_out_data_50; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_51 = mau_4_io_pipe_phv_out_data_51; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_52 = mau_4_io_pipe_phv_out_data_52; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_53 = mau_4_io_pipe_phv_out_data_53; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_54 = mau_4_io_pipe_phv_out_data_54; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_55 = mau_4_io_pipe_phv_out_data_55; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_56 = mau_4_io_pipe_phv_out_data_56; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_57 = mau_4_io_pipe_phv_out_data_57; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_58 = mau_4_io_pipe_phv_out_data_58; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_59 = mau_4_io_pipe_phv_out_data_59; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_60 = mau_4_io_pipe_phv_out_data_60; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_61 = mau_4_io_pipe_phv_out_data_61; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_62 = mau_4_io_pipe_phv_out_data_62; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_63 = mau_4_io_pipe_phv_out_data_63; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_64 = mau_4_io_pipe_phv_out_data_64; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_65 = mau_4_io_pipe_phv_out_data_65; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_66 = mau_4_io_pipe_phv_out_data_66; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_67 = mau_4_io_pipe_phv_out_data_67; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_68 = mau_4_io_pipe_phv_out_data_68; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_69 = mau_4_io_pipe_phv_out_data_69; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_70 = mau_4_io_pipe_phv_out_data_70; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_71 = mau_4_io_pipe_phv_out_data_71; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_72 = mau_4_io_pipe_phv_out_data_72; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_73 = mau_4_io_pipe_phv_out_data_73; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_74 = mau_4_io_pipe_phv_out_data_74; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_75 = mau_4_io_pipe_phv_out_data_75; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_76 = mau_4_io_pipe_phv_out_data_76; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_77 = mau_4_io_pipe_phv_out_data_77; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_78 = mau_4_io_pipe_phv_out_data_78; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_79 = mau_4_io_pipe_phv_out_data_79; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_80 = mau_4_io_pipe_phv_out_data_80; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_81 = mau_4_io_pipe_phv_out_data_81; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_82 = mau_4_io_pipe_phv_out_data_82; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_83 = mau_4_io_pipe_phv_out_data_83; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_84 = mau_4_io_pipe_phv_out_data_84; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_85 = mau_4_io_pipe_phv_out_data_85; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_86 = mau_4_io_pipe_phv_out_data_86; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_87 = mau_4_io_pipe_phv_out_data_87; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_88 = mau_4_io_pipe_phv_out_data_88; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_89 = mau_4_io_pipe_phv_out_data_89; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_90 = mau_4_io_pipe_phv_out_data_90; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_91 = mau_4_io_pipe_phv_out_data_91; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_92 = mau_4_io_pipe_phv_out_data_92; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_93 = mau_4_io_pipe_phv_out_data_93; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_94 = mau_4_io_pipe_phv_out_data_94; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_95 = mau_4_io_pipe_phv_out_data_95; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_96 = mau_4_io_pipe_phv_out_data_96; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_97 = mau_4_io_pipe_phv_out_data_97; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_98 = mau_4_io_pipe_phv_out_data_98; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_99 = mau_4_io_pipe_phv_out_data_99; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_100 = mau_4_io_pipe_phv_out_data_100; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_101 = mau_4_io_pipe_phv_out_data_101; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_102 = mau_4_io_pipe_phv_out_data_102; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_103 = mau_4_io_pipe_phv_out_data_103; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_104 = mau_4_io_pipe_phv_out_data_104; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_105 = mau_4_io_pipe_phv_out_data_105; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_106 = mau_4_io_pipe_phv_out_data_106; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_107 = mau_4_io_pipe_phv_out_data_107; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_108 = mau_4_io_pipe_phv_out_data_108; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_109 = mau_4_io_pipe_phv_out_data_109; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_110 = mau_4_io_pipe_phv_out_data_110; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_111 = mau_4_io_pipe_phv_out_data_111; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_112 = mau_4_io_pipe_phv_out_data_112; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_113 = mau_4_io_pipe_phv_out_data_113; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_114 = mau_4_io_pipe_phv_out_data_114; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_115 = mau_4_io_pipe_phv_out_data_115; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_116 = mau_4_io_pipe_phv_out_data_116; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_117 = mau_4_io_pipe_phv_out_data_117; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_118 = mau_4_io_pipe_phv_out_data_118; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_119 = mau_4_io_pipe_phv_out_data_119; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_120 = mau_4_io_pipe_phv_out_data_120; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_121 = mau_4_io_pipe_phv_out_data_121; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_122 = mau_4_io_pipe_phv_out_data_122; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_123 = mau_4_io_pipe_phv_out_data_123; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_124 = mau_4_io_pipe_phv_out_data_124; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_125 = mau_4_io_pipe_phv_out_data_125; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_126 = mau_4_io_pipe_phv_out_data_126; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_127 = mau_4_io_pipe_phv_out_data_127; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_128 = mau_4_io_pipe_phv_out_data_128; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_129 = mau_4_io_pipe_phv_out_data_129; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_130 = mau_4_io_pipe_phv_out_data_130; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_131 = mau_4_io_pipe_phv_out_data_131; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_132 = mau_4_io_pipe_phv_out_data_132; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_133 = mau_4_io_pipe_phv_out_data_133; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_134 = mau_4_io_pipe_phv_out_data_134; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_135 = mau_4_io_pipe_phv_out_data_135; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_136 = mau_4_io_pipe_phv_out_data_136; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_137 = mau_4_io_pipe_phv_out_data_137; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_138 = mau_4_io_pipe_phv_out_data_138; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_139 = mau_4_io_pipe_phv_out_data_139; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_140 = mau_4_io_pipe_phv_out_data_140; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_141 = mau_4_io_pipe_phv_out_data_141; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_142 = mau_4_io_pipe_phv_out_data_142; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_143 = mau_4_io_pipe_phv_out_data_143; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_144 = mau_4_io_pipe_phv_out_data_144; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_145 = mau_4_io_pipe_phv_out_data_145; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_146 = mau_4_io_pipe_phv_out_data_146; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_147 = mau_4_io_pipe_phv_out_data_147; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_148 = mau_4_io_pipe_phv_out_data_148; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_149 = mau_4_io_pipe_phv_out_data_149; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_150 = mau_4_io_pipe_phv_out_data_150; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_151 = mau_4_io_pipe_phv_out_data_151; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_152 = mau_4_io_pipe_phv_out_data_152; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_153 = mau_4_io_pipe_phv_out_data_153; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_154 = mau_4_io_pipe_phv_out_data_154; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_155 = mau_4_io_pipe_phv_out_data_155; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_156 = mau_4_io_pipe_phv_out_data_156; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_157 = mau_4_io_pipe_phv_out_data_157; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_158 = mau_4_io_pipe_phv_out_data_158; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_data_159 = mau_4_io_pipe_phv_out_data_159; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_0 = mau_4_io_pipe_phv_out_header_0; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_1 = mau_4_io_pipe_phv_out_header_1; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_2 = mau_4_io_pipe_phv_out_header_2; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_3 = mau_4_io_pipe_phv_out_header_3; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_4 = mau_4_io_pipe_phv_out_header_4; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_5 = mau_4_io_pipe_phv_out_header_5; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_6 = mau_4_io_pipe_phv_out_header_6; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_7 = mau_4_io_pipe_phv_out_header_7; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_8 = mau_4_io_pipe_phv_out_header_8; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_9 = mau_4_io_pipe_phv_out_header_9; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_10 = mau_4_io_pipe_phv_out_header_10; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_11 = mau_4_io_pipe_phv_out_header_11; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_12 = mau_4_io_pipe_phv_out_header_12; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_13 = mau_4_io_pipe_phv_out_header_13; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_14 = mau_4_io_pipe_phv_out_header_14; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_header_15 = mau_4_io_pipe_phv_out_header_15; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_parse_current_state = mau_4_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_parse_current_offset = mau_4_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_parse_transition_field = mau_4_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_next_processor_id = mau_4_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_next_config_id = mau_4_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_is_valid_processor = mau_4_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 42:35]
  assign mau_5_io_pipe_phv_in_valid = mau_4_io_pipe_phv_out_valid; // @[parser_pisa.scala 42:35]
  assign mau_5_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_5 :
    io_mod_module_mod_state_id_mod; // @[parser_pisa.scala 51:22 parser_pisa.scala 58:40 parser_pisa.scala 47:23]
  assign mau_5_io_mod_state_id = io_mod_module_mod_state_id; // @[parser_pisa.scala 47:23]
  assign mau_5_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser_pisa.scala 47:23]
  assign mau_5_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_5 : io_mod_module_mod_sram_w_en; // @[parser_pisa.scala 51:22 parser_pisa.scala 57:40 parser_pisa.scala 47:23]
  assign mau_5_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser_pisa.scala 47:23]
  assign mau_5_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser_pisa.scala 47:23]
  assign mau_6_clock = clock;
  assign mau_6_io_pipe_phv_in_data_0 = mau_5_io_pipe_phv_out_data_0; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_1 = mau_5_io_pipe_phv_out_data_1; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_2 = mau_5_io_pipe_phv_out_data_2; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_3 = mau_5_io_pipe_phv_out_data_3; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_4 = mau_5_io_pipe_phv_out_data_4; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_5 = mau_5_io_pipe_phv_out_data_5; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_6 = mau_5_io_pipe_phv_out_data_6; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_7 = mau_5_io_pipe_phv_out_data_7; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_8 = mau_5_io_pipe_phv_out_data_8; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_9 = mau_5_io_pipe_phv_out_data_9; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_10 = mau_5_io_pipe_phv_out_data_10; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_11 = mau_5_io_pipe_phv_out_data_11; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_12 = mau_5_io_pipe_phv_out_data_12; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_13 = mau_5_io_pipe_phv_out_data_13; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_14 = mau_5_io_pipe_phv_out_data_14; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_15 = mau_5_io_pipe_phv_out_data_15; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_16 = mau_5_io_pipe_phv_out_data_16; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_17 = mau_5_io_pipe_phv_out_data_17; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_18 = mau_5_io_pipe_phv_out_data_18; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_19 = mau_5_io_pipe_phv_out_data_19; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_20 = mau_5_io_pipe_phv_out_data_20; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_21 = mau_5_io_pipe_phv_out_data_21; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_22 = mau_5_io_pipe_phv_out_data_22; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_23 = mau_5_io_pipe_phv_out_data_23; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_24 = mau_5_io_pipe_phv_out_data_24; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_25 = mau_5_io_pipe_phv_out_data_25; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_26 = mau_5_io_pipe_phv_out_data_26; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_27 = mau_5_io_pipe_phv_out_data_27; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_28 = mau_5_io_pipe_phv_out_data_28; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_29 = mau_5_io_pipe_phv_out_data_29; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_30 = mau_5_io_pipe_phv_out_data_30; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_31 = mau_5_io_pipe_phv_out_data_31; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_32 = mau_5_io_pipe_phv_out_data_32; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_33 = mau_5_io_pipe_phv_out_data_33; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_34 = mau_5_io_pipe_phv_out_data_34; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_35 = mau_5_io_pipe_phv_out_data_35; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_36 = mau_5_io_pipe_phv_out_data_36; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_37 = mau_5_io_pipe_phv_out_data_37; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_38 = mau_5_io_pipe_phv_out_data_38; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_39 = mau_5_io_pipe_phv_out_data_39; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_40 = mau_5_io_pipe_phv_out_data_40; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_41 = mau_5_io_pipe_phv_out_data_41; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_42 = mau_5_io_pipe_phv_out_data_42; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_43 = mau_5_io_pipe_phv_out_data_43; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_44 = mau_5_io_pipe_phv_out_data_44; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_45 = mau_5_io_pipe_phv_out_data_45; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_46 = mau_5_io_pipe_phv_out_data_46; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_47 = mau_5_io_pipe_phv_out_data_47; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_48 = mau_5_io_pipe_phv_out_data_48; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_49 = mau_5_io_pipe_phv_out_data_49; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_50 = mau_5_io_pipe_phv_out_data_50; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_51 = mau_5_io_pipe_phv_out_data_51; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_52 = mau_5_io_pipe_phv_out_data_52; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_53 = mau_5_io_pipe_phv_out_data_53; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_54 = mau_5_io_pipe_phv_out_data_54; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_55 = mau_5_io_pipe_phv_out_data_55; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_56 = mau_5_io_pipe_phv_out_data_56; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_57 = mau_5_io_pipe_phv_out_data_57; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_58 = mau_5_io_pipe_phv_out_data_58; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_59 = mau_5_io_pipe_phv_out_data_59; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_60 = mau_5_io_pipe_phv_out_data_60; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_61 = mau_5_io_pipe_phv_out_data_61; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_62 = mau_5_io_pipe_phv_out_data_62; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_63 = mau_5_io_pipe_phv_out_data_63; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_64 = mau_5_io_pipe_phv_out_data_64; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_65 = mau_5_io_pipe_phv_out_data_65; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_66 = mau_5_io_pipe_phv_out_data_66; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_67 = mau_5_io_pipe_phv_out_data_67; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_68 = mau_5_io_pipe_phv_out_data_68; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_69 = mau_5_io_pipe_phv_out_data_69; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_70 = mau_5_io_pipe_phv_out_data_70; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_71 = mau_5_io_pipe_phv_out_data_71; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_72 = mau_5_io_pipe_phv_out_data_72; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_73 = mau_5_io_pipe_phv_out_data_73; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_74 = mau_5_io_pipe_phv_out_data_74; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_75 = mau_5_io_pipe_phv_out_data_75; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_76 = mau_5_io_pipe_phv_out_data_76; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_77 = mau_5_io_pipe_phv_out_data_77; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_78 = mau_5_io_pipe_phv_out_data_78; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_79 = mau_5_io_pipe_phv_out_data_79; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_80 = mau_5_io_pipe_phv_out_data_80; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_81 = mau_5_io_pipe_phv_out_data_81; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_82 = mau_5_io_pipe_phv_out_data_82; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_83 = mau_5_io_pipe_phv_out_data_83; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_84 = mau_5_io_pipe_phv_out_data_84; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_85 = mau_5_io_pipe_phv_out_data_85; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_86 = mau_5_io_pipe_phv_out_data_86; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_87 = mau_5_io_pipe_phv_out_data_87; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_88 = mau_5_io_pipe_phv_out_data_88; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_89 = mau_5_io_pipe_phv_out_data_89; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_90 = mau_5_io_pipe_phv_out_data_90; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_91 = mau_5_io_pipe_phv_out_data_91; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_92 = mau_5_io_pipe_phv_out_data_92; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_93 = mau_5_io_pipe_phv_out_data_93; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_94 = mau_5_io_pipe_phv_out_data_94; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_95 = mau_5_io_pipe_phv_out_data_95; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_96 = mau_5_io_pipe_phv_out_data_96; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_97 = mau_5_io_pipe_phv_out_data_97; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_98 = mau_5_io_pipe_phv_out_data_98; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_99 = mau_5_io_pipe_phv_out_data_99; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_100 = mau_5_io_pipe_phv_out_data_100; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_101 = mau_5_io_pipe_phv_out_data_101; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_102 = mau_5_io_pipe_phv_out_data_102; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_103 = mau_5_io_pipe_phv_out_data_103; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_104 = mau_5_io_pipe_phv_out_data_104; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_105 = mau_5_io_pipe_phv_out_data_105; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_106 = mau_5_io_pipe_phv_out_data_106; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_107 = mau_5_io_pipe_phv_out_data_107; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_108 = mau_5_io_pipe_phv_out_data_108; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_109 = mau_5_io_pipe_phv_out_data_109; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_110 = mau_5_io_pipe_phv_out_data_110; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_111 = mau_5_io_pipe_phv_out_data_111; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_112 = mau_5_io_pipe_phv_out_data_112; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_113 = mau_5_io_pipe_phv_out_data_113; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_114 = mau_5_io_pipe_phv_out_data_114; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_115 = mau_5_io_pipe_phv_out_data_115; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_116 = mau_5_io_pipe_phv_out_data_116; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_117 = mau_5_io_pipe_phv_out_data_117; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_118 = mau_5_io_pipe_phv_out_data_118; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_119 = mau_5_io_pipe_phv_out_data_119; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_120 = mau_5_io_pipe_phv_out_data_120; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_121 = mau_5_io_pipe_phv_out_data_121; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_122 = mau_5_io_pipe_phv_out_data_122; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_123 = mau_5_io_pipe_phv_out_data_123; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_124 = mau_5_io_pipe_phv_out_data_124; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_125 = mau_5_io_pipe_phv_out_data_125; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_126 = mau_5_io_pipe_phv_out_data_126; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_127 = mau_5_io_pipe_phv_out_data_127; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_128 = mau_5_io_pipe_phv_out_data_128; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_129 = mau_5_io_pipe_phv_out_data_129; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_130 = mau_5_io_pipe_phv_out_data_130; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_131 = mau_5_io_pipe_phv_out_data_131; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_132 = mau_5_io_pipe_phv_out_data_132; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_133 = mau_5_io_pipe_phv_out_data_133; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_134 = mau_5_io_pipe_phv_out_data_134; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_135 = mau_5_io_pipe_phv_out_data_135; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_136 = mau_5_io_pipe_phv_out_data_136; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_137 = mau_5_io_pipe_phv_out_data_137; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_138 = mau_5_io_pipe_phv_out_data_138; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_139 = mau_5_io_pipe_phv_out_data_139; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_140 = mau_5_io_pipe_phv_out_data_140; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_141 = mau_5_io_pipe_phv_out_data_141; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_142 = mau_5_io_pipe_phv_out_data_142; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_143 = mau_5_io_pipe_phv_out_data_143; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_144 = mau_5_io_pipe_phv_out_data_144; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_145 = mau_5_io_pipe_phv_out_data_145; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_146 = mau_5_io_pipe_phv_out_data_146; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_147 = mau_5_io_pipe_phv_out_data_147; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_148 = mau_5_io_pipe_phv_out_data_148; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_149 = mau_5_io_pipe_phv_out_data_149; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_150 = mau_5_io_pipe_phv_out_data_150; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_151 = mau_5_io_pipe_phv_out_data_151; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_152 = mau_5_io_pipe_phv_out_data_152; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_153 = mau_5_io_pipe_phv_out_data_153; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_154 = mau_5_io_pipe_phv_out_data_154; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_155 = mau_5_io_pipe_phv_out_data_155; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_156 = mau_5_io_pipe_phv_out_data_156; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_157 = mau_5_io_pipe_phv_out_data_157; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_158 = mau_5_io_pipe_phv_out_data_158; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_data_159 = mau_5_io_pipe_phv_out_data_159; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_0 = mau_5_io_pipe_phv_out_header_0; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_1 = mau_5_io_pipe_phv_out_header_1; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_2 = mau_5_io_pipe_phv_out_header_2; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_3 = mau_5_io_pipe_phv_out_header_3; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_4 = mau_5_io_pipe_phv_out_header_4; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_5 = mau_5_io_pipe_phv_out_header_5; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_6 = mau_5_io_pipe_phv_out_header_6; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_7 = mau_5_io_pipe_phv_out_header_7; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_8 = mau_5_io_pipe_phv_out_header_8; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_9 = mau_5_io_pipe_phv_out_header_9; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_10 = mau_5_io_pipe_phv_out_header_10; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_11 = mau_5_io_pipe_phv_out_header_11; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_12 = mau_5_io_pipe_phv_out_header_12; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_13 = mau_5_io_pipe_phv_out_header_13; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_14 = mau_5_io_pipe_phv_out_header_14; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_header_15 = mau_5_io_pipe_phv_out_header_15; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_parse_current_state = mau_5_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_parse_current_offset = mau_5_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_parse_transition_field = mau_5_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_next_processor_id = mau_5_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_next_config_id = mau_5_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_is_valid_processor = mau_5_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 42:35]
  assign mau_6_io_pipe_phv_in_valid = mau_5_io_pipe_phv_out_valid; // @[parser_pisa.scala 42:35]
  assign mau_6_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_6 :
    io_mod_module_mod_state_id_mod; // @[parser_pisa.scala 51:22 parser_pisa.scala 58:40 parser_pisa.scala 47:23]
  assign mau_6_io_mod_state_id = io_mod_module_mod_state_id; // @[parser_pisa.scala 47:23]
  assign mau_6_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser_pisa.scala 47:23]
  assign mau_6_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_6 : io_mod_module_mod_sram_w_en; // @[parser_pisa.scala 51:22 parser_pisa.scala 57:40 parser_pisa.scala 47:23]
  assign mau_6_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser_pisa.scala 47:23]
  assign mau_6_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser_pisa.scala 47:23]
  assign mau_7_clock = clock;
  assign mau_7_io_pipe_phv_in_data_0 = mau_6_io_pipe_phv_out_data_0; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_1 = mau_6_io_pipe_phv_out_data_1; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_2 = mau_6_io_pipe_phv_out_data_2; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_3 = mau_6_io_pipe_phv_out_data_3; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_4 = mau_6_io_pipe_phv_out_data_4; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_5 = mau_6_io_pipe_phv_out_data_5; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_6 = mau_6_io_pipe_phv_out_data_6; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_7 = mau_6_io_pipe_phv_out_data_7; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_8 = mau_6_io_pipe_phv_out_data_8; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_9 = mau_6_io_pipe_phv_out_data_9; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_10 = mau_6_io_pipe_phv_out_data_10; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_11 = mau_6_io_pipe_phv_out_data_11; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_12 = mau_6_io_pipe_phv_out_data_12; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_13 = mau_6_io_pipe_phv_out_data_13; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_14 = mau_6_io_pipe_phv_out_data_14; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_15 = mau_6_io_pipe_phv_out_data_15; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_16 = mau_6_io_pipe_phv_out_data_16; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_17 = mau_6_io_pipe_phv_out_data_17; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_18 = mau_6_io_pipe_phv_out_data_18; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_19 = mau_6_io_pipe_phv_out_data_19; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_20 = mau_6_io_pipe_phv_out_data_20; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_21 = mau_6_io_pipe_phv_out_data_21; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_22 = mau_6_io_pipe_phv_out_data_22; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_23 = mau_6_io_pipe_phv_out_data_23; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_24 = mau_6_io_pipe_phv_out_data_24; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_25 = mau_6_io_pipe_phv_out_data_25; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_26 = mau_6_io_pipe_phv_out_data_26; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_27 = mau_6_io_pipe_phv_out_data_27; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_28 = mau_6_io_pipe_phv_out_data_28; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_29 = mau_6_io_pipe_phv_out_data_29; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_30 = mau_6_io_pipe_phv_out_data_30; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_31 = mau_6_io_pipe_phv_out_data_31; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_32 = mau_6_io_pipe_phv_out_data_32; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_33 = mau_6_io_pipe_phv_out_data_33; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_34 = mau_6_io_pipe_phv_out_data_34; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_35 = mau_6_io_pipe_phv_out_data_35; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_36 = mau_6_io_pipe_phv_out_data_36; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_37 = mau_6_io_pipe_phv_out_data_37; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_38 = mau_6_io_pipe_phv_out_data_38; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_39 = mau_6_io_pipe_phv_out_data_39; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_40 = mau_6_io_pipe_phv_out_data_40; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_41 = mau_6_io_pipe_phv_out_data_41; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_42 = mau_6_io_pipe_phv_out_data_42; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_43 = mau_6_io_pipe_phv_out_data_43; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_44 = mau_6_io_pipe_phv_out_data_44; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_45 = mau_6_io_pipe_phv_out_data_45; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_46 = mau_6_io_pipe_phv_out_data_46; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_47 = mau_6_io_pipe_phv_out_data_47; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_48 = mau_6_io_pipe_phv_out_data_48; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_49 = mau_6_io_pipe_phv_out_data_49; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_50 = mau_6_io_pipe_phv_out_data_50; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_51 = mau_6_io_pipe_phv_out_data_51; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_52 = mau_6_io_pipe_phv_out_data_52; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_53 = mau_6_io_pipe_phv_out_data_53; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_54 = mau_6_io_pipe_phv_out_data_54; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_55 = mau_6_io_pipe_phv_out_data_55; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_56 = mau_6_io_pipe_phv_out_data_56; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_57 = mau_6_io_pipe_phv_out_data_57; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_58 = mau_6_io_pipe_phv_out_data_58; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_59 = mau_6_io_pipe_phv_out_data_59; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_60 = mau_6_io_pipe_phv_out_data_60; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_61 = mau_6_io_pipe_phv_out_data_61; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_62 = mau_6_io_pipe_phv_out_data_62; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_63 = mau_6_io_pipe_phv_out_data_63; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_64 = mau_6_io_pipe_phv_out_data_64; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_65 = mau_6_io_pipe_phv_out_data_65; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_66 = mau_6_io_pipe_phv_out_data_66; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_67 = mau_6_io_pipe_phv_out_data_67; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_68 = mau_6_io_pipe_phv_out_data_68; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_69 = mau_6_io_pipe_phv_out_data_69; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_70 = mau_6_io_pipe_phv_out_data_70; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_71 = mau_6_io_pipe_phv_out_data_71; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_72 = mau_6_io_pipe_phv_out_data_72; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_73 = mau_6_io_pipe_phv_out_data_73; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_74 = mau_6_io_pipe_phv_out_data_74; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_75 = mau_6_io_pipe_phv_out_data_75; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_76 = mau_6_io_pipe_phv_out_data_76; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_77 = mau_6_io_pipe_phv_out_data_77; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_78 = mau_6_io_pipe_phv_out_data_78; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_79 = mau_6_io_pipe_phv_out_data_79; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_80 = mau_6_io_pipe_phv_out_data_80; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_81 = mau_6_io_pipe_phv_out_data_81; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_82 = mau_6_io_pipe_phv_out_data_82; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_83 = mau_6_io_pipe_phv_out_data_83; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_84 = mau_6_io_pipe_phv_out_data_84; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_85 = mau_6_io_pipe_phv_out_data_85; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_86 = mau_6_io_pipe_phv_out_data_86; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_87 = mau_6_io_pipe_phv_out_data_87; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_88 = mau_6_io_pipe_phv_out_data_88; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_89 = mau_6_io_pipe_phv_out_data_89; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_90 = mau_6_io_pipe_phv_out_data_90; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_91 = mau_6_io_pipe_phv_out_data_91; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_92 = mau_6_io_pipe_phv_out_data_92; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_93 = mau_6_io_pipe_phv_out_data_93; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_94 = mau_6_io_pipe_phv_out_data_94; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_95 = mau_6_io_pipe_phv_out_data_95; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_96 = mau_6_io_pipe_phv_out_data_96; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_97 = mau_6_io_pipe_phv_out_data_97; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_98 = mau_6_io_pipe_phv_out_data_98; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_99 = mau_6_io_pipe_phv_out_data_99; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_100 = mau_6_io_pipe_phv_out_data_100; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_101 = mau_6_io_pipe_phv_out_data_101; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_102 = mau_6_io_pipe_phv_out_data_102; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_103 = mau_6_io_pipe_phv_out_data_103; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_104 = mau_6_io_pipe_phv_out_data_104; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_105 = mau_6_io_pipe_phv_out_data_105; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_106 = mau_6_io_pipe_phv_out_data_106; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_107 = mau_6_io_pipe_phv_out_data_107; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_108 = mau_6_io_pipe_phv_out_data_108; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_109 = mau_6_io_pipe_phv_out_data_109; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_110 = mau_6_io_pipe_phv_out_data_110; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_111 = mau_6_io_pipe_phv_out_data_111; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_112 = mau_6_io_pipe_phv_out_data_112; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_113 = mau_6_io_pipe_phv_out_data_113; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_114 = mau_6_io_pipe_phv_out_data_114; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_115 = mau_6_io_pipe_phv_out_data_115; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_116 = mau_6_io_pipe_phv_out_data_116; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_117 = mau_6_io_pipe_phv_out_data_117; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_118 = mau_6_io_pipe_phv_out_data_118; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_119 = mau_6_io_pipe_phv_out_data_119; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_120 = mau_6_io_pipe_phv_out_data_120; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_121 = mau_6_io_pipe_phv_out_data_121; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_122 = mau_6_io_pipe_phv_out_data_122; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_123 = mau_6_io_pipe_phv_out_data_123; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_124 = mau_6_io_pipe_phv_out_data_124; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_125 = mau_6_io_pipe_phv_out_data_125; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_126 = mau_6_io_pipe_phv_out_data_126; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_127 = mau_6_io_pipe_phv_out_data_127; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_128 = mau_6_io_pipe_phv_out_data_128; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_129 = mau_6_io_pipe_phv_out_data_129; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_130 = mau_6_io_pipe_phv_out_data_130; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_131 = mau_6_io_pipe_phv_out_data_131; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_132 = mau_6_io_pipe_phv_out_data_132; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_133 = mau_6_io_pipe_phv_out_data_133; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_134 = mau_6_io_pipe_phv_out_data_134; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_135 = mau_6_io_pipe_phv_out_data_135; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_136 = mau_6_io_pipe_phv_out_data_136; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_137 = mau_6_io_pipe_phv_out_data_137; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_138 = mau_6_io_pipe_phv_out_data_138; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_139 = mau_6_io_pipe_phv_out_data_139; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_140 = mau_6_io_pipe_phv_out_data_140; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_141 = mau_6_io_pipe_phv_out_data_141; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_142 = mau_6_io_pipe_phv_out_data_142; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_143 = mau_6_io_pipe_phv_out_data_143; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_144 = mau_6_io_pipe_phv_out_data_144; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_145 = mau_6_io_pipe_phv_out_data_145; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_146 = mau_6_io_pipe_phv_out_data_146; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_147 = mau_6_io_pipe_phv_out_data_147; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_148 = mau_6_io_pipe_phv_out_data_148; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_149 = mau_6_io_pipe_phv_out_data_149; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_150 = mau_6_io_pipe_phv_out_data_150; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_151 = mau_6_io_pipe_phv_out_data_151; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_152 = mau_6_io_pipe_phv_out_data_152; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_153 = mau_6_io_pipe_phv_out_data_153; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_154 = mau_6_io_pipe_phv_out_data_154; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_155 = mau_6_io_pipe_phv_out_data_155; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_156 = mau_6_io_pipe_phv_out_data_156; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_157 = mau_6_io_pipe_phv_out_data_157; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_158 = mau_6_io_pipe_phv_out_data_158; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_data_159 = mau_6_io_pipe_phv_out_data_159; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_0 = mau_6_io_pipe_phv_out_header_0; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_1 = mau_6_io_pipe_phv_out_header_1; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_2 = mau_6_io_pipe_phv_out_header_2; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_3 = mau_6_io_pipe_phv_out_header_3; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_4 = mau_6_io_pipe_phv_out_header_4; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_5 = mau_6_io_pipe_phv_out_header_5; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_6 = mau_6_io_pipe_phv_out_header_6; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_7 = mau_6_io_pipe_phv_out_header_7; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_8 = mau_6_io_pipe_phv_out_header_8; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_9 = mau_6_io_pipe_phv_out_header_9; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_10 = mau_6_io_pipe_phv_out_header_10; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_11 = mau_6_io_pipe_phv_out_header_11; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_12 = mau_6_io_pipe_phv_out_header_12; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_13 = mau_6_io_pipe_phv_out_header_13; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_14 = mau_6_io_pipe_phv_out_header_14; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_header_15 = mau_6_io_pipe_phv_out_header_15; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_parse_current_state = mau_6_io_pipe_phv_out_parse_current_state; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_parse_current_offset = mau_6_io_pipe_phv_out_parse_current_offset; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_parse_transition_field = mau_6_io_pipe_phv_out_parse_transition_field; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_next_processor_id = mau_6_io_pipe_phv_out_next_processor_id; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_next_config_id = mau_6_io_pipe_phv_out_next_config_id; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_is_valid_processor = mau_6_io_pipe_phv_out_is_valid_processor; // @[parser_pisa.scala 42:35]
  assign mau_7_io_pipe_phv_in_valid = mau_6_io_pipe_phv_out_valid; // @[parser_pisa.scala 42:35]
  assign mau_7_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_7 :
    io_mod_module_mod_state_id_mod; // @[parser_pisa.scala 51:22 parser_pisa.scala 58:40 parser_pisa.scala 47:23]
  assign mau_7_io_mod_state_id = io_mod_module_mod_state_id; // @[parser_pisa.scala 47:23]
  assign mau_7_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser_pisa.scala 47:23]
  assign mau_7_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_7 : io_mod_module_mod_sram_w_en; // @[parser_pisa.scala 51:22 parser_pisa.scala 57:40 parser_pisa.scala 47:23]
  assign mau_7_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser_pisa.scala 47:23]
  assign mau_7_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser_pisa.scala 47:23]
  always @(posedge clock) begin
    if (io_mod_en) begin // @[parser_pisa.scala 51:22]
      if (io_mod_last_mau_id_mod) begin // @[parser_pisa.scala 52:39]
        last_mau_id <= io_mod_last_mau_id; // @[parser_pisa.scala 53:25]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  last_mau_id = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
