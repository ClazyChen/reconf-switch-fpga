module AXISIdle(
  input          clock,
  input          reset,
  input          io_s_axis_tvalid,
  output         io_s_axis_tready,
  input  [511:0] io_s_axis_tdata,
  input  [63:0]  io_s_axis_tkeep,
  input          io_s_axis_tlast,
  output         io_m_axis_tvalid,
  input          io_m_axis_tready,
  output [511:0] io_m_axis_tdata,
  output [63:0]  io_m_axis_tkeep,
  output         io_m_axis_tlast
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
`endif // RANDOMIZE_REG_INIT
  wire  in_axi_clock; // @[tester.scala 16:24]
  wire  in_axi_reset; // @[tester.scala 16:24]
  wire  in_axi_io_s_axis_tvalid; // @[tester.scala 16:24]
  wire [511:0] in_axi_io_s_axis_tdata; // @[tester.scala 16:24]
  wire  in_axi_io_s_axis_tlast; // @[tester.scala 16:24]
  wire  in_axi_io_ipsa_en_in; // @[tester.scala 16:24]
  wire  in_axi_io_ipsa_last_in; // @[tester.scala 16:24]
  wire [1023:0] in_axi_io_ipsa_data_in; // @[tester.scala 16:24]
  wire  out_axi_clock; // @[tester.scala 17:25]
  wire  out_axi_reset; // @[tester.scala 17:25]
  wire  out_axi_io_m_axis_tready; // @[tester.scala 17:25]
  wire [511:0] out_axi_io_m_axis_tdata; // @[tester.scala 17:25]
  wire  out_axi_io_m_axis_tlast; // @[tester.scala 17:25]
  wire  out_axi_io_ipsa_last_out; // @[tester.scala 17:25]
  wire  out_axi_io_ipsa_en_out; // @[tester.scala 17:25]
  wire [1023:0] out_axi_io_ipsa_data_out; // @[tester.scala 17:25]
  wire  in_port_io_en; // @[tester.scala 18:25]
  wire  in_port_io_last; // @[tester.scala 18:25]
  wire [1023:0] in_port_io_data; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_0; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_1; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_2; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_3; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_4; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_5; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_6; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_7; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_8; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_9; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_10; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_11; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_12; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_13; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_14; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_15; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_16; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_17; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_18; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_19; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_20; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_21; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_22; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_23; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_24; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_25; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_26; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_27; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_28; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_29; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_30; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_31; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_32; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_33; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_34; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_35; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_36; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_37; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_38; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_39; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_40; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_41; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_42; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_43; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_44; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_45; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_46; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_47; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_48; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_49; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_50; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_51; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_52; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_53; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_54; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_55; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_56; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_57; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_58; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_59; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_60; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_61; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_62; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_63; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_64; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_65; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_66; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_67; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_68; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_69; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_70; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_71; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_72; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_73; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_74; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_75; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_76; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_77; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_78; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_79; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_80; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_81; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_82; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_83; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_84; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_85; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_86; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_87; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_88; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_89; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_90; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_91; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_92; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_93; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_94; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_95; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_96; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_97; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_98; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_99; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_100; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_101; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_102; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_103; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_104; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_105; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_106; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_107; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_108; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_109; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_110; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_111; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_112; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_113; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_114; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_115; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_116; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_117; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_118; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_119; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_120; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_121; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_122; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_123; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_124; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_125; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_126; // @[tester.scala 18:25]
  wire [7:0] in_port_io_phv_out_data_127; // @[tester.scala 18:25]
  wire  in_port_io_phv_out_valid; // @[tester.scala 18:25]
  wire  in_port_io_phv_out_last; // @[tester.scala 18:25]
  wire [7:0] out_port_io_phv_in_data_0; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_1; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_2; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_3; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_4; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_5; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_6; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_7; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_8; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_9; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_10; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_11; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_12; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_13; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_14; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_15; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_16; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_17; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_18; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_19; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_20; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_21; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_22; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_23; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_24; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_25; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_26; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_27; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_28; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_29; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_30; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_31; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_32; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_33; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_34; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_35; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_36; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_37; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_38; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_39; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_40; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_41; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_42; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_43; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_44; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_45; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_46; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_47; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_48; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_49; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_50; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_51; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_52; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_53; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_54; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_55; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_56; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_57; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_58; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_59; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_60; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_61; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_62; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_63; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_64; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_65; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_66; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_67; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_68; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_69; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_70; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_71; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_72; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_73; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_74; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_75; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_76; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_77; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_78; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_79; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_80; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_81; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_82; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_83; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_84; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_85; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_86; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_87; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_88; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_89; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_90; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_91; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_92; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_93; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_94; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_95; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_96; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_97; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_98; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_99; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_100; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_101; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_102; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_103; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_104; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_105; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_106; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_107; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_108; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_109; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_110; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_111; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_112; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_113; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_114; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_115; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_116; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_117; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_118; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_119; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_120; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_121; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_122; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_123; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_124; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_125; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_126; // @[tester.scala 19:26]
  wire [7:0] out_port_io_phv_in_data_127; // @[tester.scala 19:26]
  wire  out_port_io_phv_in_valid; // @[tester.scala 19:26]
  wire  out_port_io_phv_in_last; // @[tester.scala 19:26]
  wire [1023:0] out_port_io_data; // @[tester.scala 19:26]
  wire  out_port_io_last; // @[tester.scala 19:26]
  wire  out_port_io_en; // @[tester.scala 19:26]
  reg [7:0] phv1_data_0; // @[tester.scala 21:19]
  reg [7:0] phv1_data_1; // @[tester.scala 21:19]
  reg [7:0] phv1_data_2; // @[tester.scala 21:19]
  reg [7:0] phv1_data_3; // @[tester.scala 21:19]
  reg [7:0] phv1_data_4; // @[tester.scala 21:19]
  reg [7:0] phv1_data_5; // @[tester.scala 21:19]
  reg [7:0] phv1_data_6; // @[tester.scala 21:19]
  reg [7:0] phv1_data_7; // @[tester.scala 21:19]
  reg [7:0] phv1_data_8; // @[tester.scala 21:19]
  reg [7:0] phv1_data_9; // @[tester.scala 21:19]
  reg [7:0] phv1_data_10; // @[tester.scala 21:19]
  reg [7:0] phv1_data_11; // @[tester.scala 21:19]
  reg [7:0] phv1_data_12; // @[tester.scala 21:19]
  reg [7:0] phv1_data_13; // @[tester.scala 21:19]
  reg [7:0] phv1_data_14; // @[tester.scala 21:19]
  reg [7:0] phv1_data_15; // @[tester.scala 21:19]
  reg [7:0] phv1_data_16; // @[tester.scala 21:19]
  reg [7:0] phv1_data_17; // @[tester.scala 21:19]
  reg [7:0] phv1_data_18; // @[tester.scala 21:19]
  reg [7:0] phv1_data_19; // @[tester.scala 21:19]
  reg [7:0] phv1_data_20; // @[tester.scala 21:19]
  reg [7:0] phv1_data_21; // @[tester.scala 21:19]
  reg [7:0] phv1_data_22; // @[tester.scala 21:19]
  reg [7:0] phv1_data_23; // @[tester.scala 21:19]
  reg [7:0] phv1_data_24; // @[tester.scala 21:19]
  reg [7:0] phv1_data_25; // @[tester.scala 21:19]
  reg [7:0] phv1_data_26; // @[tester.scala 21:19]
  reg [7:0] phv1_data_27; // @[tester.scala 21:19]
  reg [7:0] phv1_data_28; // @[tester.scala 21:19]
  reg [7:0] phv1_data_29; // @[tester.scala 21:19]
  reg [7:0] phv1_data_30; // @[tester.scala 21:19]
  reg [7:0] phv1_data_31; // @[tester.scala 21:19]
  reg [7:0] phv1_data_32; // @[tester.scala 21:19]
  reg [7:0] phv1_data_33; // @[tester.scala 21:19]
  reg [7:0] phv1_data_34; // @[tester.scala 21:19]
  reg [7:0] phv1_data_35; // @[tester.scala 21:19]
  reg [7:0] phv1_data_36; // @[tester.scala 21:19]
  reg [7:0] phv1_data_37; // @[tester.scala 21:19]
  reg [7:0] phv1_data_38; // @[tester.scala 21:19]
  reg [7:0] phv1_data_39; // @[tester.scala 21:19]
  reg [7:0] phv1_data_40; // @[tester.scala 21:19]
  reg [7:0] phv1_data_41; // @[tester.scala 21:19]
  reg [7:0] phv1_data_42; // @[tester.scala 21:19]
  reg [7:0] phv1_data_43; // @[tester.scala 21:19]
  reg [7:0] phv1_data_44; // @[tester.scala 21:19]
  reg [7:0] phv1_data_45; // @[tester.scala 21:19]
  reg [7:0] phv1_data_46; // @[tester.scala 21:19]
  reg [7:0] phv1_data_47; // @[tester.scala 21:19]
  reg [7:0] phv1_data_48; // @[tester.scala 21:19]
  reg [7:0] phv1_data_49; // @[tester.scala 21:19]
  reg [7:0] phv1_data_50; // @[tester.scala 21:19]
  reg [7:0] phv1_data_51; // @[tester.scala 21:19]
  reg [7:0] phv1_data_52; // @[tester.scala 21:19]
  reg [7:0] phv1_data_53; // @[tester.scala 21:19]
  reg [7:0] phv1_data_54; // @[tester.scala 21:19]
  reg [7:0] phv1_data_55; // @[tester.scala 21:19]
  reg [7:0] phv1_data_56; // @[tester.scala 21:19]
  reg [7:0] phv1_data_57; // @[tester.scala 21:19]
  reg [7:0] phv1_data_58; // @[tester.scala 21:19]
  reg [7:0] phv1_data_59; // @[tester.scala 21:19]
  reg [7:0] phv1_data_60; // @[tester.scala 21:19]
  reg [7:0] phv1_data_61; // @[tester.scala 21:19]
  reg [7:0] phv1_data_62; // @[tester.scala 21:19]
  reg [7:0] phv1_data_63; // @[tester.scala 21:19]
  reg [7:0] phv1_data_64; // @[tester.scala 21:19]
  reg [7:0] phv1_data_65; // @[tester.scala 21:19]
  reg [7:0] phv1_data_66; // @[tester.scala 21:19]
  reg [7:0] phv1_data_67; // @[tester.scala 21:19]
  reg [7:0] phv1_data_68; // @[tester.scala 21:19]
  reg [7:0] phv1_data_69; // @[tester.scala 21:19]
  reg [7:0] phv1_data_70; // @[tester.scala 21:19]
  reg [7:0] phv1_data_71; // @[tester.scala 21:19]
  reg [7:0] phv1_data_72; // @[tester.scala 21:19]
  reg [7:0] phv1_data_73; // @[tester.scala 21:19]
  reg [7:0] phv1_data_74; // @[tester.scala 21:19]
  reg [7:0] phv1_data_75; // @[tester.scala 21:19]
  reg [7:0] phv1_data_76; // @[tester.scala 21:19]
  reg [7:0] phv1_data_77; // @[tester.scala 21:19]
  reg [7:0] phv1_data_78; // @[tester.scala 21:19]
  reg [7:0] phv1_data_79; // @[tester.scala 21:19]
  reg [7:0] phv1_data_80; // @[tester.scala 21:19]
  reg [7:0] phv1_data_81; // @[tester.scala 21:19]
  reg [7:0] phv1_data_82; // @[tester.scala 21:19]
  reg [7:0] phv1_data_83; // @[tester.scala 21:19]
  reg [7:0] phv1_data_84; // @[tester.scala 21:19]
  reg [7:0] phv1_data_85; // @[tester.scala 21:19]
  reg [7:0] phv1_data_86; // @[tester.scala 21:19]
  reg [7:0] phv1_data_87; // @[tester.scala 21:19]
  reg [7:0] phv1_data_88; // @[tester.scala 21:19]
  reg [7:0] phv1_data_89; // @[tester.scala 21:19]
  reg [7:0] phv1_data_90; // @[tester.scala 21:19]
  reg [7:0] phv1_data_91; // @[tester.scala 21:19]
  reg [7:0] phv1_data_92; // @[tester.scala 21:19]
  reg [7:0] phv1_data_93; // @[tester.scala 21:19]
  reg [7:0] phv1_data_94; // @[tester.scala 21:19]
  reg [7:0] phv1_data_95; // @[tester.scala 21:19]
  reg [7:0] phv1_data_96; // @[tester.scala 21:19]
  reg [7:0] phv1_data_97; // @[tester.scala 21:19]
  reg [7:0] phv1_data_98; // @[tester.scala 21:19]
  reg [7:0] phv1_data_99; // @[tester.scala 21:19]
  reg [7:0] phv1_data_100; // @[tester.scala 21:19]
  reg [7:0] phv1_data_101; // @[tester.scala 21:19]
  reg [7:0] phv1_data_102; // @[tester.scala 21:19]
  reg [7:0] phv1_data_103; // @[tester.scala 21:19]
  reg [7:0] phv1_data_104; // @[tester.scala 21:19]
  reg [7:0] phv1_data_105; // @[tester.scala 21:19]
  reg [7:0] phv1_data_106; // @[tester.scala 21:19]
  reg [7:0] phv1_data_107; // @[tester.scala 21:19]
  reg [7:0] phv1_data_108; // @[tester.scala 21:19]
  reg [7:0] phv1_data_109; // @[tester.scala 21:19]
  reg [7:0] phv1_data_110; // @[tester.scala 21:19]
  reg [7:0] phv1_data_111; // @[tester.scala 21:19]
  reg [7:0] phv1_data_112; // @[tester.scala 21:19]
  reg [7:0] phv1_data_113; // @[tester.scala 21:19]
  reg [7:0] phv1_data_114; // @[tester.scala 21:19]
  reg [7:0] phv1_data_115; // @[tester.scala 21:19]
  reg [7:0] phv1_data_116; // @[tester.scala 21:19]
  reg [7:0] phv1_data_117; // @[tester.scala 21:19]
  reg [7:0] phv1_data_118; // @[tester.scala 21:19]
  reg [7:0] phv1_data_119; // @[tester.scala 21:19]
  reg [7:0] phv1_data_120; // @[tester.scala 21:19]
  reg [7:0] phv1_data_121; // @[tester.scala 21:19]
  reg [7:0] phv1_data_122; // @[tester.scala 21:19]
  reg [7:0] phv1_data_123; // @[tester.scala 21:19]
  reg [7:0] phv1_data_124; // @[tester.scala 21:19]
  reg [7:0] phv1_data_125; // @[tester.scala 21:19]
  reg [7:0] phv1_data_126; // @[tester.scala 21:19]
  reg [7:0] phv1_data_127; // @[tester.scala 21:19]
  reg  phv1_valid; // @[tester.scala 21:19]
  reg  phv1_last; // @[tester.scala 21:19]
  reg [7:0] phv2_data_0; // @[tester.scala 22:19]
  reg [7:0] phv2_data_1; // @[tester.scala 22:19]
  reg [7:0] phv2_data_2; // @[tester.scala 22:19]
  reg [7:0] phv2_data_3; // @[tester.scala 22:19]
  reg [7:0] phv2_data_4; // @[tester.scala 22:19]
  reg [7:0] phv2_data_5; // @[tester.scala 22:19]
  reg [7:0] phv2_data_6; // @[tester.scala 22:19]
  reg [7:0] phv2_data_7; // @[tester.scala 22:19]
  reg [7:0] phv2_data_8; // @[tester.scala 22:19]
  reg [7:0] phv2_data_9; // @[tester.scala 22:19]
  reg [7:0] phv2_data_10; // @[tester.scala 22:19]
  reg [7:0] phv2_data_11; // @[tester.scala 22:19]
  reg [7:0] phv2_data_12; // @[tester.scala 22:19]
  reg [7:0] phv2_data_13; // @[tester.scala 22:19]
  reg [7:0] phv2_data_14; // @[tester.scala 22:19]
  reg [7:0] phv2_data_15; // @[tester.scala 22:19]
  reg [7:0] phv2_data_16; // @[tester.scala 22:19]
  reg [7:0] phv2_data_17; // @[tester.scala 22:19]
  reg [7:0] phv2_data_18; // @[tester.scala 22:19]
  reg [7:0] phv2_data_19; // @[tester.scala 22:19]
  reg [7:0] phv2_data_20; // @[tester.scala 22:19]
  reg [7:0] phv2_data_21; // @[tester.scala 22:19]
  reg [7:0] phv2_data_22; // @[tester.scala 22:19]
  reg [7:0] phv2_data_23; // @[tester.scala 22:19]
  reg [7:0] phv2_data_24; // @[tester.scala 22:19]
  reg [7:0] phv2_data_25; // @[tester.scala 22:19]
  reg [7:0] phv2_data_26; // @[tester.scala 22:19]
  reg [7:0] phv2_data_27; // @[tester.scala 22:19]
  reg [7:0] phv2_data_28; // @[tester.scala 22:19]
  reg [7:0] phv2_data_29; // @[tester.scala 22:19]
  reg [7:0] phv2_data_30; // @[tester.scala 22:19]
  reg [7:0] phv2_data_31; // @[tester.scala 22:19]
  reg [7:0] phv2_data_32; // @[tester.scala 22:19]
  reg [7:0] phv2_data_33; // @[tester.scala 22:19]
  reg [7:0] phv2_data_34; // @[tester.scala 22:19]
  reg [7:0] phv2_data_35; // @[tester.scala 22:19]
  reg [7:0] phv2_data_36; // @[tester.scala 22:19]
  reg [7:0] phv2_data_37; // @[tester.scala 22:19]
  reg [7:0] phv2_data_38; // @[tester.scala 22:19]
  reg [7:0] phv2_data_39; // @[tester.scala 22:19]
  reg [7:0] phv2_data_40; // @[tester.scala 22:19]
  reg [7:0] phv2_data_41; // @[tester.scala 22:19]
  reg [7:0] phv2_data_42; // @[tester.scala 22:19]
  reg [7:0] phv2_data_43; // @[tester.scala 22:19]
  reg [7:0] phv2_data_44; // @[tester.scala 22:19]
  reg [7:0] phv2_data_45; // @[tester.scala 22:19]
  reg [7:0] phv2_data_46; // @[tester.scala 22:19]
  reg [7:0] phv2_data_47; // @[tester.scala 22:19]
  reg [7:0] phv2_data_48; // @[tester.scala 22:19]
  reg [7:0] phv2_data_49; // @[tester.scala 22:19]
  reg [7:0] phv2_data_50; // @[tester.scala 22:19]
  reg [7:0] phv2_data_51; // @[tester.scala 22:19]
  reg [7:0] phv2_data_52; // @[tester.scala 22:19]
  reg [7:0] phv2_data_53; // @[tester.scala 22:19]
  reg [7:0] phv2_data_54; // @[tester.scala 22:19]
  reg [7:0] phv2_data_55; // @[tester.scala 22:19]
  reg [7:0] phv2_data_56; // @[tester.scala 22:19]
  reg [7:0] phv2_data_57; // @[tester.scala 22:19]
  reg [7:0] phv2_data_58; // @[tester.scala 22:19]
  reg [7:0] phv2_data_59; // @[tester.scala 22:19]
  reg [7:0] phv2_data_60; // @[tester.scala 22:19]
  reg [7:0] phv2_data_61; // @[tester.scala 22:19]
  reg [7:0] phv2_data_62; // @[tester.scala 22:19]
  reg [7:0] phv2_data_63; // @[tester.scala 22:19]
  reg [7:0] phv2_data_64; // @[tester.scala 22:19]
  reg [7:0] phv2_data_65; // @[tester.scala 22:19]
  reg [7:0] phv2_data_66; // @[tester.scala 22:19]
  reg [7:0] phv2_data_67; // @[tester.scala 22:19]
  reg [7:0] phv2_data_68; // @[tester.scala 22:19]
  reg [7:0] phv2_data_69; // @[tester.scala 22:19]
  reg [7:0] phv2_data_70; // @[tester.scala 22:19]
  reg [7:0] phv2_data_71; // @[tester.scala 22:19]
  reg [7:0] phv2_data_72; // @[tester.scala 22:19]
  reg [7:0] phv2_data_73; // @[tester.scala 22:19]
  reg [7:0] phv2_data_74; // @[tester.scala 22:19]
  reg [7:0] phv2_data_75; // @[tester.scala 22:19]
  reg [7:0] phv2_data_76; // @[tester.scala 22:19]
  reg [7:0] phv2_data_77; // @[tester.scala 22:19]
  reg [7:0] phv2_data_78; // @[tester.scala 22:19]
  reg [7:0] phv2_data_79; // @[tester.scala 22:19]
  reg [7:0] phv2_data_80; // @[tester.scala 22:19]
  reg [7:0] phv2_data_81; // @[tester.scala 22:19]
  reg [7:0] phv2_data_82; // @[tester.scala 22:19]
  reg [7:0] phv2_data_83; // @[tester.scala 22:19]
  reg [7:0] phv2_data_84; // @[tester.scala 22:19]
  reg [7:0] phv2_data_85; // @[tester.scala 22:19]
  reg [7:0] phv2_data_86; // @[tester.scala 22:19]
  reg [7:0] phv2_data_87; // @[tester.scala 22:19]
  reg [7:0] phv2_data_88; // @[tester.scala 22:19]
  reg [7:0] phv2_data_89; // @[tester.scala 22:19]
  reg [7:0] phv2_data_90; // @[tester.scala 22:19]
  reg [7:0] phv2_data_91; // @[tester.scala 22:19]
  reg [7:0] phv2_data_92; // @[tester.scala 22:19]
  reg [7:0] phv2_data_93; // @[tester.scala 22:19]
  reg [7:0] phv2_data_94; // @[tester.scala 22:19]
  reg [7:0] phv2_data_95; // @[tester.scala 22:19]
  reg [7:0] phv2_data_96; // @[tester.scala 22:19]
  reg [7:0] phv2_data_97; // @[tester.scala 22:19]
  reg [7:0] phv2_data_98; // @[tester.scala 22:19]
  reg [7:0] phv2_data_99; // @[tester.scala 22:19]
  reg [7:0] phv2_data_100; // @[tester.scala 22:19]
  reg [7:0] phv2_data_101; // @[tester.scala 22:19]
  reg [7:0] phv2_data_102; // @[tester.scala 22:19]
  reg [7:0] phv2_data_103; // @[tester.scala 22:19]
  reg [7:0] phv2_data_104; // @[tester.scala 22:19]
  reg [7:0] phv2_data_105; // @[tester.scala 22:19]
  reg [7:0] phv2_data_106; // @[tester.scala 22:19]
  reg [7:0] phv2_data_107; // @[tester.scala 22:19]
  reg [7:0] phv2_data_108; // @[tester.scala 22:19]
  reg [7:0] phv2_data_109; // @[tester.scala 22:19]
  reg [7:0] phv2_data_110; // @[tester.scala 22:19]
  reg [7:0] phv2_data_111; // @[tester.scala 22:19]
  reg [7:0] phv2_data_112; // @[tester.scala 22:19]
  reg [7:0] phv2_data_113; // @[tester.scala 22:19]
  reg [7:0] phv2_data_114; // @[tester.scala 22:19]
  reg [7:0] phv2_data_115; // @[tester.scala 22:19]
  reg [7:0] phv2_data_116; // @[tester.scala 22:19]
  reg [7:0] phv2_data_117; // @[tester.scala 22:19]
  reg [7:0] phv2_data_118; // @[tester.scala 22:19]
  reg [7:0] phv2_data_119; // @[tester.scala 22:19]
  reg [7:0] phv2_data_120; // @[tester.scala 22:19]
  reg [7:0] phv2_data_121; // @[tester.scala 22:19]
  reg [7:0] phv2_data_122; // @[tester.scala 22:19]
  reg [7:0] phv2_data_123; // @[tester.scala 22:19]
  reg [7:0] phv2_data_124; // @[tester.scala 22:19]
  reg [7:0] phv2_data_125; // @[tester.scala 22:19]
  reg [7:0] phv2_data_126; // @[tester.scala 22:19]
  reg [7:0] phv2_data_127; // @[tester.scala 22:19]
  reg  phv2_valid; // @[tester.scala 22:19]
  reg  phv2_last; // @[tester.scala 22:19]
  InAXI in_axi ( // @[tester.scala 16:24]
    .clock(in_axi_clock),
    .reset(in_axi_reset),
    .io_s_axis_tvalid(in_axi_io_s_axis_tvalid),
    .io_s_axis_tdata(in_axi_io_s_axis_tdata),
    .io_s_axis_tlast(in_axi_io_s_axis_tlast),
    .io_ipsa_en_in(in_axi_io_ipsa_en_in),
    .io_ipsa_last_in(in_axi_io_ipsa_last_in),
    .io_ipsa_data_in(in_axi_io_ipsa_data_in)
  );
  OutAXI out_axi ( // @[tester.scala 17:25]
    .clock(out_axi_clock),
    .reset(out_axi_reset),
    .io_m_axis_tready(out_axi_io_m_axis_tready),
    .io_m_axis_tdata(out_axi_io_m_axis_tdata),
    .io_m_axis_tlast(out_axi_io_m_axis_tlast),
    .io_ipsa_last_out(out_axi_io_ipsa_last_out),
    .io_ipsa_en_out(out_axi_io_ipsa_en_out),
    .io_ipsa_data_out(out_axi_io_ipsa_data_out)
  );
  InPort in_port ( // @[tester.scala 18:25]
    .io_en(in_port_io_en),
    .io_last(in_port_io_last),
    .io_data(in_port_io_data),
    .io_phv_out_data_0(in_port_io_phv_out_data_0),
    .io_phv_out_data_1(in_port_io_phv_out_data_1),
    .io_phv_out_data_2(in_port_io_phv_out_data_2),
    .io_phv_out_data_3(in_port_io_phv_out_data_3),
    .io_phv_out_data_4(in_port_io_phv_out_data_4),
    .io_phv_out_data_5(in_port_io_phv_out_data_5),
    .io_phv_out_data_6(in_port_io_phv_out_data_6),
    .io_phv_out_data_7(in_port_io_phv_out_data_7),
    .io_phv_out_data_8(in_port_io_phv_out_data_8),
    .io_phv_out_data_9(in_port_io_phv_out_data_9),
    .io_phv_out_data_10(in_port_io_phv_out_data_10),
    .io_phv_out_data_11(in_port_io_phv_out_data_11),
    .io_phv_out_data_12(in_port_io_phv_out_data_12),
    .io_phv_out_data_13(in_port_io_phv_out_data_13),
    .io_phv_out_data_14(in_port_io_phv_out_data_14),
    .io_phv_out_data_15(in_port_io_phv_out_data_15),
    .io_phv_out_data_16(in_port_io_phv_out_data_16),
    .io_phv_out_data_17(in_port_io_phv_out_data_17),
    .io_phv_out_data_18(in_port_io_phv_out_data_18),
    .io_phv_out_data_19(in_port_io_phv_out_data_19),
    .io_phv_out_data_20(in_port_io_phv_out_data_20),
    .io_phv_out_data_21(in_port_io_phv_out_data_21),
    .io_phv_out_data_22(in_port_io_phv_out_data_22),
    .io_phv_out_data_23(in_port_io_phv_out_data_23),
    .io_phv_out_data_24(in_port_io_phv_out_data_24),
    .io_phv_out_data_25(in_port_io_phv_out_data_25),
    .io_phv_out_data_26(in_port_io_phv_out_data_26),
    .io_phv_out_data_27(in_port_io_phv_out_data_27),
    .io_phv_out_data_28(in_port_io_phv_out_data_28),
    .io_phv_out_data_29(in_port_io_phv_out_data_29),
    .io_phv_out_data_30(in_port_io_phv_out_data_30),
    .io_phv_out_data_31(in_port_io_phv_out_data_31),
    .io_phv_out_data_32(in_port_io_phv_out_data_32),
    .io_phv_out_data_33(in_port_io_phv_out_data_33),
    .io_phv_out_data_34(in_port_io_phv_out_data_34),
    .io_phv_out_data_35(in_port_io_phv_out_data_35),
    .io_phv_out_data_36(in_port_io_phv_out_data_36),
    .io_phv_out_data_37(in_port_io_phv_out_data_37),
    .io_phv_out_data_38(in_port_io_phv_out_data_38),
    .io_phv_out_data_39(in_port_io_phv_out_data_39),
    .io_phv_out_data_40(in_port_io_phv_out_data_40),
    .io_phv_out_data_41(in_port_io_phv_out_data_41),
    .io_phv_out_data_42(in_port_io_phv_out_data_42),
    .io_phv_out_data_43(in_port_io_phv_out_data_43),
    .io_phv_out_data_44(in_port_io_phv_out_data_44),
    .io_phv_out_data_45(in_port_io_phv_out_data_45),
    .io_phv_out_data_46(in_port_io_phv_out_data_46),
    .io_phv_out_data_47(in_port_io_phv_out_data_47),
    .io_phv_out_data_48(in_port_io_phv_out_data_48),
    .io_phv_out_data_49(in_port_io_phv_out_data_49),
    .io_phv_out_data_50(in_port_io_phv_out_data_50),
    .io_phv_out_data_51(in_port_io_phv_out_data_51),
    .io_phv_out_data_52(in_port_io_phv_out_data_52),
    .io_phv_out_data_53(in_port_io_phv_out_data_53),
    .io_phv_out_data_54(in_port_io_phv_out_data_54),
    .io_phv_out_data_55(in_port_io_phv_out_data_55),
    .io_phv_out_data_56(in_port_io_phv_out_data_56),
    .io_phv_out_data_57(in_port_io_phv_out_data_57),
    .io_phv_out_data_58(in_port_io_phv_out_data_58),
    .io_phv_out_data_59(in_port_io_phv_out_data_59),
    .io_phv_out_data_60(in_port_io_phv_out_data_60),
    .io_phv_out_data_61(in_port_io_phv_out_data_61),
    .io_phv_out_data_62(in_port_io_phv_out_data_62),
    .io_phv_out_data_63(in_port_io_phv_out_data_63),
    .io_phv_out_data_64(in_port_io_phv_out_data_64),
    .io_phv_out_data_65(in_port_io_phv_out_data_65),
    .io_phv_out_data_66(in_port_io_phv_out_data_66),
    .io_phv_out_data_67(in_port_io_phv_out_data_67),
    .io_phv_out_data_68(in_port_io_phv_out_data_68),
    .io_phv_out_data_69(in_port_io_phv_out_data_69),
    .io_phv_out_data_70(in_port_io_phv_out_data_70),
    .io_phv_out_data_71(in_port_io_phv_out_data_71),
    .io_phv_out_data_72(in_port_io_phv_out_data_72),
    .io_phv_out_data_73(in_port_io_phv_out_data_73),
    .io_phv_out_data_74(in_port_io_phv_out_data_74),
    .io_phv_out_data_75(in_port_io_phv_out_data_75),
    .io_phv_out_data_76(in_port_io_phv_out_data_76),
    .io_phv_out_data_77(in_port_io_phv_out_data_77),
    .io_phv_out_data_78(in_port_io_phv_out_data_78),
    .io_phv_out_data_79(in_port_io_phv_out_data_79),
    .io_phv_out_data_80(in_port_io_phv_out_data_80),
    .io_phv_out_data_81(in_port_io_phv_out_data_81),
    .io_phv_out_data_82(in_port_io_phv_out_data_82),
    .io_phv_out_data_83(in_port_io_phv_out_data_83),
    .io_phv_out_data_84(in_port_io_phv_out_data_84),
    .io_phv_out_data_85(in_port_io_phv_out_data_85),
    .io_phv_out_data_86(in_port_io_phv_out_data_86),
    .io_phv_out_data_87(in_port_io_phv_out_data_87),
    .io_phv_out_data_88(in_port_io_phv_out_data_88),
    .io_phv_out_data_89(in_port_io_phv_out_data_89),
    .io_phv_out_data_90(in_port_io_phv_out_data_90),
    .io_phv_out_data_91(in_port_io_phv_out_data_91),
    .io_phv_out_data_92(in_port_io_phv_out_data_92),
    .io_phv_out_data_93(in_port_io_phv_out_data_93),
    .io_phv_out_data_94(in_port_io_phv_out_data_94),
    .io_phv_out_data_95(in_port_io_phv_out_data_95),
    .io_phv_out_data_96(in_port_io_phv_out_data_96),
    .io_phv_out_data_97(in_port_io_phv_out_data_97),
    .io_phv_out_data_98(in_port_io_phv_out_data_98),
    .io_phv_out_data_99(in_port_io_phv_out_data_99),
    .io_phv_out_data_100(in_port_io_phv_out_data_100),
    .io_phv_out_data_101(in_port_io_phv_out_data_101),
    .io_phv_out_data_102(in_port_io_phv_out_data_102),
    .io_phv_out_data_103(in_port_io_phv_out_data_103),
    .io_phv_out_data_104(in_port_io_phv_out_data_104),
    .io_phv_out_data_105(in_port_io_phv_out_data_105),
    .io_phv_out_data_106(in_port_io_phv_out_data_106),
    .io_phv_out_data_107(in_port_io_phv_out_data_107),
    .io_phv_out_data_108(in_port_io_phv_out_data_108),
    .io_phv_out_data_109(in_port_io_phv_out_data_109),
    .io_phv_out_data_110(in_port_io_phv_out_data_110),
    .io_phv_out_data_111(in_port_io_phv_out_data_111),
    .io_phv_out_data_112(in_port_io_phv_out_data_112),
    .io_phv_out_data_113(in_port_io_phv_out_data_113),
    .io_phv_out_data_114(in_port_io_phv_out_data_114),
    .io_phv_out_data_115(in_port_io_phv_out_data_115),
    .io_phv_out_data_116(in_port_io_phv_out_data_116),
    .io_phv_out_data_117(in_port_io_phv_out_data_117),
    .io_phv_out_data_118(in_port_io_phv_out_data_118),
    .io_phv_out_data_119(in_port_io_phv_out_data_119),
    .io_phv_out_data_120(in_port_io_phv_out_data_120),
    .io_phv_out_data_121(in_port_io_phv_out_data_121),
    .io_phv_out_data_122(in_port_io_phv_out_data_122),
    .io_phv_out_data_123(in_port_io_phv_out_data_123),
    .io_phv_out_data_124(in_port_io_phv_out_data_124),
    .io_phv_out_data_125(in_port_io_phv_out_data_125),
    .io_phv_out_data_126(in_port_io_phv_out_data_126),
    .io_phv_out_data_127(in_port_io_phv_out_data_127),
    .io_phv_out_valid(in_port_io_phv_out_valid),
    .io_phv_out_last(in_port_io_phv_out_last)
  );
  OutPort out_port ( // @[tester.scala 19:26]
    .io_phv_in_data_0(out_port_io_phv_in_data_0),
    .io_phv_in_data_1(out_port_io_phv_in_data_1),
    .io_phv_in_data_2(out_port_io_phv_in_data_2),
    .io_phv_in_data_3(out_port_io_phv_in_data_3),
    .io_phv_in_data_4(out_port_io_phv_in_data_4),
    .io_phv_in_data_5(out_port_io_phv_in_data_5),
    .io_phv_in_data_6(out_port_io_phv_in_data_6),
    .io_phv_in_data_7(out_port_io_phv_in_data_7),
    .io_phv_in_data_8(out_port_io_phv_in_data_8),
    .io_phv_in_data_9(out_port_io_phv_in_data_9),
    .io_phv_in_data_10(out_port_io_phv_in_data_10),
    .io_phv_in_data_11(out_port_io_phv_in_data_11),
    .io_phv_in_data_12(out_port_io_phv_in_data_12),
    .io_phv_in_data_13(out_port_io_phv_in_data_13),
    .io_phv_in_data_14(out_port_io_phv_in_data_14),
    .io_phv_in_data_15(out_port_io_phv_in_data_15),
    .io_phv_in_data_16(out_port_io_phv_in_data_16),
    .io_phv_in_data_17(out_port_io_phv_in_data_17),
    .io_phv_in_data_18(out_port_io_phv_in_data_18),
    .io_phv_in_data_19(out_port_io_phv_in_data_19),
    .io_phv_in_data_20(out_port_io_phv_in_data_20),
    .io_phv_in_data_21(out_port_io_phv_in_data_21),
    .io_phv_in_data_22(out_port_io_phv_in_data_22),
    .io_phv_in_data_23(out_port_io_phv_in_data_23),
    .io_phv_in_data_24(out_port_io_phv_in_data_24),
    .io_phv_in_data_25(out_port_io_phv_in_data_25),
    .io_phv_in_data_26(out_port_io_phv_in_data_26),
    .io_phv_in_data_27(out_port_io_phv_in_data_27),
    .io_phv_in_data_28(out_port_io_phv_in_data_28),
    .io_phv_in_data_29(out_port_io_phv_in_data_29),
    .io_phv_in_data_30(out_port_io_phv_in_data_30),
    .io_phv_in_data_31(out_port_io_phv_in_data_31),
    .io_phv_in_data_32(out_port_io_phv_in_data_32),
    .io_phv_in_data_33(out_port_io_phv_in_data_33),
    .io_phv_in_data_34(out_port_io_phv_in_data_34),
    .io_phv_in_data_35(out_port_io_phv_in_data_35),
    .io_phv_in_data_36(out_port_io_phv_in_data_36),
    .io_phv_in_data_37(out_port_io_phv_in_data_37),
    .io_phv_in_data_38(out_port_io_phv_in_data_38),
    .io_phv_in_data_39(out_port_io_phv_in_data_39),
    .io_phv_in_data_40(out_port_io_phv_in_data_40),
    .io_phv_in_data_41(out_port_io_phv_in_data_41),
    .io_phv_in_data_42(out_port_io_phv_in_data_42),
    .io_phv_in_data_43(out_port_io_phv_in_data_43),
    .io_phv_in_data_44(out_port_io_phv_in_data_44),
    .io_phv_in_data_45(out_port_io_phv_in_data_45),
    .io_phv_in_data_46(out_port_io_phv_in_data_46),
    .io_phv_in_data_47(out_port_io_phv_in_data_47),
    .io_phv_in_data_48(out_port_io_phv_in_data_48),
    .io_phv_in_data_49(out_port_io_phv_in_data_49),
    .io_phv_in_data_50(out_port_io_phv_in_data_50),
    .io_phv_in_data_51(out_port_io_phv_in_data_51),
    .io_phv_in_data_52(out_port_io_phv_in_data_52),
    .io_phv_in_data_53(out_port_io_phv_in_data_53),
    .io_phv_in_data_54(out_port_io_phv_in_data_54),
    .io_phv_in_data_55(out_port_io_phv_in_data_55),
    .io_phv_in_data_56(out_port_io_phv_in_data_56),
    .io_phv_in_data_57(out_port_io_phv_in_data_57),
    .io_phv_in_data_58(out_port_io_phv_in_data_58),
    .io_phv_in_data_59(out_port_io_phv_in_data_59),
    .io_phv_in_data_60(out_port_io_phv_in_data_60),
    .io_phv_in_data_61(out_port_io_phv_in_data_61),
    .io_phv_in_data_62(out_port_io_phv_in_data_62),
    .io_phv_in_data_63(out_port_io_phv_in_data_63),
    .io_phv_in_data_64(out_port_io_phv_in_data_64),
    .io_phv_in_data_65(out_port_io_phv_in_data_65),
    .io_phv_in_data_66(out_port_io_phv_in_data_66),
    .io_phv_in_data_67(out_port_io_phv_in_data_67),
    .io_phv_in_data_68(out_port_io_phv_in_data_68),
    .io_phv_in_data_69(out_port_io_phv_in_data_69),
    .io_phv_in_data_70(out_port_io_phv_in_data_70),
    .io_phv_in_data_71(out_port_io_phv_in_data_71),
    .io_phv_in_data_72(out_port_io_phv_in_data_72),
    .io_phv_in_data_73(out_port_io_phv_in_data_73),
    .io_phv_in_data_74(out_port_io_phv_in_data_74),
    .io_phv_in_data_75(out_port_io_phv_in_data_75),
    .io_phv_in_data_76(out_port_io_phv_in_data_76),
    .io_phv_in_data_77(out_port_io_phv_in_data_77),
    .io_phv_in_data_78(out_port_io_phv_in_data_78),
    .io_phv_in_data_79(out_port_io_phv_in_data_79),
    .io_phv_in_data_80(out_port_io_phv_in_data_80),
    .io_phv_in_data_81(out_port_io_phv_in_data_81),
    .io_phv_in_data_82(out_port_io_phv_in_data_82),
    .io_phv_in_data_83(out_port_io_phv_in_data_83),
    .io_phv_in_data_84(out_port_io_phv_in_data_84),
    .io_phv_in_data_85(out_port_io_phv_in_data_85),
    .io_phv_in_data_86(out_port_io_phv_in_data_86),
    .io_phv_in_data_87(out_port_io_phv_in_data_87),
    .io_phv_in_data_88(out_port_io_phv_in_data_88),
    .io_phv_in_data_89(out_port_io_phv_in_data_89),
    .io_phv_in_data_90(out_port_io_phv_in_data_90),
    .io_phv_in_data_91(out_port_io_phv_in_data_91),
    .io_phv_in_data_92(out_port_io_phv_in_data_92),
    .io_phv_in_data_93(out_port_io_phv_in_data_93),
    .io_phv_in_data_94(out_port_io_phv_in_data_94),
    .io_phv_in_data_95(out_port_io_phv_in_data_95),
    .io_phv_in_data_96(out_port_io_phv_in_data_96),
    .io_phv_in_data_97(out_port_io_phv_in_data_97),
    .io_phv_in_data_98(out_port_io_phv_in_data_98),
    .io_phv_in_data_99(out_port_io_phv_in_data_99),
    .io_phv_in_data_100(out_port_io_phv_in_data_100),
    .io_phv_in_data_101(out_port_io_phv_in_data_101),
    .io_phv_in_data_102(out_port_io_phv_in_data_102),
    .io_phv_in_data_103(out_port_io_phv_in_data_103),
    .io_phv_in_data_104(out_port_io_phv_in_data_104),
    .io_phv_in_data_105(out_port_io_phv_in_data_105),
    .io_phv_in_data_106(out_port_io_phv_in_data_106),
    .io_phv_in_data_107(out_port_io_phv_in_data_107),
    .io_phv_in_data_108(out_port_io_phv_in_data_108),
    .io_phv_in_data_109(out_port_io_phv_in_data_109),
    .io_phv_in_data_110(out_port_io_phv_in_data_110),
    .io_phv_in_data_111(out_port_io_phv_in_data_111),
    .io_phv_in_data_112(out_port_io_phv_in_data_112),
    .io_phv_in_data_113(out_port_io_phv_in_data_113),
    .io_phv_in_data_114(out_port_io_phv_in_data_114),
    .io_phv_in_data_115(out_port_io_phv_in_data_115),
    .io_phv_in_data_116(out_port_io_phv_in_data_116),
    .io_phv_in_data_117(out_port_io_phv_in_data_117),
    .io_phv_in_data_118(out_port_io_phv_in_data_118),
    .io_phv_in_data_119(out_port_io_phv_in_data_119),
    .io_phv_in_data_120(out_port_io_phv_in_data_120),
    .io_phv_in_data_121(out_port_io_phv_in_data_121),
    .io_phv_in_data_122(out_port_io_phv_in_data_122),
    .io_phv_in_data_123(out_port_io_phv_in_data_123),
    .io_phv_in_data_124(out_port_io_phv_in_data_124),
    .io_phv_in_data_125(out_port_io_phv_in_data_125),
    .io_phv_in_data_126(out_port_io_phv_in_data_126),
    .io_phv_in_data_127(out_port_io_phv_in_data_127),
    .io_phv_in_valid(out_port_io_phv_in_valid),
    .io_phv_in_last(out_port_io_phv_in_last),
    .io_data(out_port_io_data),
    .io_last(out_port_io_last),
    .io_en(out_port_io_en)
  );
  assign io_s_axis_tready = 1'h1; // @[tester.scala 23:22]
  assign io_m_axis_tvalid = 1'h1; // @[tester.scala 39:23]
  assign io_m_axis_tdata = out_axi_io_m_axis_tdata; // @[tester.scala 39:23]
  assign io_m_axis_tkeep = 64'hffffffffffffffff; // @[tester.scala 39:23]
  assign io_m_axis_tlast = out_axi_io_m_axis_tlast; // @[tester.scala 39:23]
  assign in_axi_clock = clock;
  assign in_axi_reset = reset;
  assign in_axi_io_s_axis_tvalid = io_s_axis_tvalid; // @[tester.scala 23:22]
  assign in_axi_io_s_axis_tdata = io_s_axis_tdata; // @[tester.scala 23:22]
  assign in_axi_io_s_axis_tlast = io_s_axis_tlast; // @[tester.scala 23:22]
  assign out_axi_clock = clock;
  assign out_axi_reset = reset;
  assign out_axi_io_m_axis_tready = io_m_axis_tready; // @[tester.scala 39:23]
  assign out_axi_io_ipsa_last_out = out_port_io_last; // @[tester.scala 41:30]
  assign out_axi_io_ipsa_en_out = out_port_io_en; // @[tester.scala 40:28]
  assign out_axi_io_ipsa_data_out = out_port_io_data; // @[tester.scala 42:30]
  assign in_port_io_en = in_axi_io_ipsa_en_in; // @[tester.scala 24:26]
  assign in_port_io_last = in_axi_io_ipsa_last_in; // @[tester.scala 25:28]
  assign in_port_io_data = in_axi_io_ipsa_data_in; // @[tester.scala 26:28]
  assign out_port_io_phv_in_data_0 = phv2_data_0; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_1 = phv2_data_1; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_2 = phv2_data_2; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_3 = phv2_data_3; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_4 = phv2_data_4; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_5 = phv2_data_5; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_6 = phv2_data_6; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_7 = phv2_data_7; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_8 = phv2_data_8; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_9 = phv2_data_9; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_10 = phv2_data_10; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_11 = phv2_data_11; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_12 = phv2_data_12; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_13 = phv2_data_13; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_14 = phv2_data_14; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_15 = phv2_data_15; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_16 = phv2_data_16; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_17 = phv2_data_17; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_18 = phv2_data_18; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_19 = phv2_data_19; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_20 = phv2_data_20; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_21 = phv2_data_21; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_22 = phv2_data_22; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_23 = phv2_data_23; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_24 = phv2_data_24; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_25 = phv2_data_25; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_26 = phv2_data_26; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_27 = phv2_data_27; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_28 = phv2_data_28; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_29 = phv2_data_29; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_30 = phv2_data_30; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_31 = phv2_data_31; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_32 = phv2_data_32; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_33 = phv2_data_33; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_34 = phv2_data_34; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_35 = phv2_data_35; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_36 = phv2_data_36; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_37 = phv2_data_37; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_38 = phv2_data_38; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_39 = phv2_data_39; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_40 = phv2_data_40; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_41 = phv2_data_41; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_42 = phv2_data_42; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_43 = phv2_data_43; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_44 = phv2_data_44; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_45 = phv2_data_45; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_46 = phv2_data_46; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_47 = phv2_data_47; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_48 = phv2_data_48; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_49 = phv2_data_49; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_50 = phv2_data_50; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_51 = phv2_data_51; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_52 = phv2_data_52; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_53 = phv2_data_53; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_54 = phv2_data_54; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_55 = phv2_data_55; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_56 = phv2_data_56; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_57 = phv2_data_57; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_58 = phv2_data_58; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_59 = phv2_data_59; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_60 = phv2_data_60; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_61 = phv2_data_61; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_62 = phv2_data_62; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_63 = phv2_data_63; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_64 = phv2_data_64; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_65 = phv2_data_65; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_66 = phv2_data_66; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_67 = phv2_data_67; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_68 = phv2_data_68; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_69 = phv2_data_69; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_70 = phv2_data_70; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_71 = phv2_data_71; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_72 = phv2_data_72; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_73 = phv2_data_73; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_74 = phv2_data_74; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_75 = phv2_data_75; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_76 = phv2_data_76; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_77 = phv2_data_77; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_78 = phv2_data_78; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_79 = phv2_data_79; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_80 = phv2_data_80; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_81 = phv2_data_81; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_82 = phv2_data_82; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_83 = phv2_data_83; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_84 = phv2_data_84; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_85 = phv2_data_85; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_86 = phv2_data_86; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_87 = phv2_data_87; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_88 = phv2_data_88; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_89 = phv2_data_89; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_90 = phv2_data_90; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_91 = phv2_data_91; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_92 = phv2_data_92; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_93 = phv2_data_93; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_94 = phv2_data_94; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_95 = phv2_data_95; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_96 = phv2_data_96; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_97 = phv2_data_97; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_98 = phv2_data_98; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_99 = phv2_data_99; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_100 = phv2_data_100; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_101 = phv2_data_101; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_102 = phv2_data_102; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_103 = phv2_data_103; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_104 = phv2_data_104; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_105 = phv2_data_105; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_106 = phv2_data_106; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_107 = phv2_data_107; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_108 = phv2_data_108; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_109 = phv2_data_109; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_110 = phv2_data_110; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_111 = phv2_data_111; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_112 = phv2_data_112; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_113 = phv2_data_113; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_114 = phv2_data_114; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_115 = phv2_data_115; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_116 = phv2_data_116; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_117 = phv2_data_117; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_118 = phv2_data_118; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_119 = phv2_data_119; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_120 = phv2_data_120; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_121 = phv2_data_121; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_122 = phv2_data_122; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_123 = phv2_data_123; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_124 = phv2_data_124; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_125 = phv2_data_125; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_126 = phv2_data_126; // @[tester.scala 33:24]
  assign out_port_io_phv_in_data_127 = phv2_data_127; // @[tester.scala 33:24]
  assign out_port_io_phv_in_valid = phv2_valid; // @[tester.scala 33:24]
  assign out_port_io_phv_in_last = phv2_last; // @[tester.scala 33:24]
  always @(posedge clock) begin
    phv1_data_0 <= in_port_io_phv_out_data_0; // @[tester.scala 31:10]
    phv1_data_1 <= in_port_io_phv_out_data_1; // @[tester.scala 31:10]
    phv1_data_2 <= in_port_io_phv_out_data_2; // @[tester.scala 31:10]
    phv1_data_3 <= in_port_io_phv_out_data_3; // @[tester.scala 31:10]
    phv1_data_4 <= in_port_io_phv_out_data_4; // @[tester.scala 31:10]
    phv1_data_5 <= in_port_io_phv_out_data_5; // @[tester.scala 31:10]
    phv1_data_6 <= in_port_io_phv_out_data_6; // @[tester.scala 31:10]
    phv1_data_7 <= in_port_io_phv_out_data_7; // @[tester.scala 31:10]
    phv1_data_8 <= in_port_io_phv_out_data_8; // @[tester.scala 31:10]
    phv1_data_9 <= in_port_io_phv_out_data_9; // @[tester.scala 31:10]
    phv1_data_10 <= in_port_io_phv_out_data_10; // @[tester.scala 31:10]
    phv1_data_11 <= in_port_io_phv_out_data_11; // @[tester.scala 31:10]
    phv1_data_12 <= in_port_io_phv_out_data_12; // @[tester.scala 31:10]
    phv1_data_13 <= in_port_io_phv_out_data_13; // @[tester.scala 31:10]
    phv1_data_14 <= in_port_io_phv_out_data_14; // @[tester.scala 31:10]
    phv1_data_15 <= in_port_io_phv_out_data_15; // @[tester.scala 31:10]
    phv1_data_16 <= in_port_io_phv_out_data_16; // @[tester.scala 31:10]
    phv1_data_17 <= in_port_io_phv_out_data_17; // @[tester.scala 31:10]
    phv1_data_18 <= in_port_io_phv_out_data_18; // @[tester.scala 31:10]
    phv1_data_19 <= in_port_io_phv_out_data_19; // @[tester.scala 31:10]
    phv1_data_20 <= in_port_io_phv_out_data_20; // @[tester.scala 31:10]
    phv1_data_21 <= in_port_io_phv_out_data_21; // @[tester.scala 31:10]
    phv1_data_22 <= in_port_io_phv_out_data_22; // @[tester.scala 31:10]
    phv1_data_23 <= in_port_io_phv_out_data_23; // @[tester.scala 31:10]
    phv1_data_24 <= in_port_io_phv_out_data_24; // @[tester.scala 31:10]
    phv1_data_25 <= in_port_io_phv_out_data_25; // @[tester.scala 31:10]
    phv1_data_26 <= in_port_io_phv_out_data_26; // @[tester.scala 31:10]
    phv1_data_27 <= in_port_io_phv_out_data_27; // @[tester.scala 31:10]
    phv1_data_28 <= in_port_io_phv_out_data_28; // @[tester.scala 31:10]
    phv1_data_29 <= in_port_io_phv_out_data_29; // @[tester.scala 31:10]
    phv1_data_30 <= in_port_io_phv_out_data_30; // @[tester.scala 31:10]
    phv1_data_31 <= in_port_io_phv_out_data_31; // @[tester.scala 31:10]
    phv1_data_32 <= in_port_io_phv_out_data_32; // @[tester.scala 31:10]
    phv1_data_33 <= in_port_io_phv_out_data_33; // @[tester.scala 31:10]
    phv1_data_34 <= in_port_io_phv_out_data_34; // @[tester.scala 31:10]
    phv1_data_35 <= in_port_io_phv_out_data_35; // @[tester.scala 31:10]
    phv1_data_36 <= in_port_io_phv_out_data_36; // @[tester.scala 31:10]
    phv1_data_37 <= in_port_io_phv_out_data_37; // @[tester.scala 31:10]
    phv1_data_38 <= in_port_io_phv_out_data_38; // @[tester.scala 31:10]
    phv1_data_39 <= in_port_io_phv_out_data_39; // @[tester.scala 31:10]
    phv1_data_40 <= in_port_io_phv_out_data_40; // @[tester.scala 31:10]
    phv1_data_41 <= in_port_io_phv_out_data_41; // @[tester.scala 31:10]
    phv1_data_42 <= in_port_io_phv_out_data_42; // @[tester.scala 31:10]
    phv1_data_43 <= in_port_io_phv_out_data_43; // @[tester.scala 31:10]
    phv1_data_44 <= in_port_io_phv_out_data_44; // @[tester.scala 31:10]
    phv1_data_45 <= in_port_io_phv_out_data_45; // @[tester.scala 31:10]
    phv1_data_46 <= in_port_io_phv_out_data_46; // @[tester.scala 31:10]
    phv1_data_47 <= in_port_io_phv_out_data_47; // @[tester.scala 31:10]
    phv1_data_48 <= in_port_io_phv_out_data_48; // @[tester.scala 31:10]
    phv1_data_49 <= in_port_io_phv_out_data_49; // @[tester.scala 31:10]
    phv1_data_50 <= in_port_io_phv_out_data_50; // @[tester.scala 31:10]
    phv1_data_51 <= in_port_io_phv_out_data_51; // @[tester.scala 31:10]
    phv1_data_52 <= in_port_io_phv_out_data_52; // @[tester.scala 31:10]
    phv1_data_53 <= in_port_io_phv_out_data_53; // @[tester.scala 31:10]
    phv1_data_54 <= in_port_io_phv_out_data_54; // @[tester.scala 31:10]
    phv1_data_55 <= in_port_io_phv_out_data_55; // @[tester.scala 31:10]
    phv1_data_56 <= in_port_io_phv_out_data_56; // @[tester.scala 31:10]
    phv1_data_57 <= in_port_io_phv_out_data_57; // @[tester.scala 31:10]
    phv1_data_58 <= in_port_io_phv_out_data_58; // @[tester.scala 31:10]
    phv1_data_59 <= in_port_io_phv_out_data_59; // @[tester.scala 31:10]
    phv1_data_60 <= in_port_io_phv_out_data_60; // @[tester.scala 31:10]
    phv1_data_61 <= in_port_io_phv_out_data_61; // @[tester.scala 31:10]
    phv1_data_62 <= in_port_io_phv_out_data_62; // @[tester.scala 31:10]
    phv1_data_63 <= in_port_io_phv_out_data_63; // @[tester.scala 31:10]
    phv1_data_64 <= in_port_io_phv_out_data_64; // @[tester.scala 31:10]
    phv1_data_65 <= in_port_io_phv_out_data_65; // @[tester.scala 31:10]
    phv1_data_66 <= in_port_io_phv_out_data_66; // @[tester.scala 31:10]
    phv1_data_67 <= in_port_io_phv_out_data_67; // @[tester.scala 31:10]
    phv1_data_68 <= in_port_io_phv_out_data_68; // @[tester.scala 31:10]
    phv1_data_69 <= in_port_io_phv_out_data_69; // @[tester.scala 31:10]
    phv1_data_70 <= in_port_io_phv_out_data_70; // @[tester.scala 31:10]
    phv1_data_71 <= in_port_io_phv_out_data_71; // @[tester.scala 31:10]
    phv1_data_72 <= in_port_io_phv_out_data_72; // @[tester.scala 31:10]
    phv1_data_73 <= in_port_io_phv_out_data_73; // @[tester.scala 31:10]
    phv1_data_74 <= in_port_io_phv_out_data_74; // @[tester.scala 31:10]
    phv1_data_75 <= in_port_io_phv_out_data_75; // @[tester.scala 31:10]
    phv1_data_76 <= in_port_io_phv_out_data_76; // @[tester.scala 31:10]
    phv1_data_77 <= in_port_io_phv_out_data_77; // @[tester.scala 31:10]
    phv1_data_78 <= in_port_io_phv_out_data_78; // @[tester.scala 31:10]
    phv1_data_79 <= in_port_io_phv_out_data_79; // @[tester.scala 31:10]
    phv1_data_80 <= in_port_io_phv_out_data_80; // @[tester.scala 31:10]
    phv1_data_81 <= in_port_io_phv_out_data_81; // @[tester.scala 31:10]
    phv1_data_82 <= in_port_io_phv_out_data_82; // @[tester.scala 31:10]
    phv1_data_83 <= in_port_io_phv_out_data_83; // @[tester.scala 31:10]
    phv1_data_84 <= in_port_io_phv_out_data_84; // @[tester.scala 31:10]
    phv1_data_85 <= in_port_io_phv_out_data_85; // @[tester.scala 31:10]
    phv1_data_86 <= in_port_io_phv_out_data_86; // @[tester.scala 31:10]
    phv1_data_87 <= in_port_io_phv_out_data_87; // @[tester.scala 31:10]
    phv1_data_88 <= in_port_io_phv_out_data_88; // @[tester.scala 31:10]
    phv1_data_89 <= in_port_io_phv_out_data_89; // @[tester.scala 31:10]
    phv1_data_90 <= in_port_io_phv_out_data_90; // @[tester.scala 31:10]
    phv1_data_91 <= in_port_io_phv_out_data_91; // @[tester.scala 31:10]
    phv1_data_92 <= in_port_io_phv_out_data_92; // @[tester.scala 31:10]
    phv1_data_93 <= in_port_io_phv_out_data_93; // @[tester.scala 31:10]
    phv1_data_94 <= in_port_io_phv_out_data_94; // @[tester.scala 31:10]
    phv1_data_95 <= in_port_io_phv_out_data_95; // @[tester.scala 31:10]
    phv1_data_96 <= in_port_io_phv_out_data_96; // @[tester.scala 31:10]
    phv1_data_97 <= in_port_io_phv_out_data_97; // @[tester.scala 31:10]
    phv1_data_98 <= in_port_io_phv_out_data_98; // @[tester.scala 31:10]
    phv1_data_99 <= in_port_io_phv_out_data_99; // @[tester.scala 31:10]
    phv1_data_100 <= in_port_io_phv_out_data_100; // @[tester.scala 31:10]
    phv1_data_101 <= in_port_io_phv_out_data_101; // @[tester.scala 31:10]
    phv1_data_102 <= in_port_io_phv_out_data_102; // @[tester.scala 31:10]
    phv1_data_103 <= in_port_io_phv_out_data_103; // @[tester.scala 31:10]
    phv1_data_104 <= in_port_io_phv_out_data_104; // @[tester.scala 31:10]
    phv1_data_105 <= in_port_io_phv_out_data_105; // @[tester.scala 31:10]
    phv1_data_106 <= in_port_io_phv_out_data_106; // @[tester.scala 31:10]
    phv1_data_107 <= in_port_io_phv_out_data_107; // @[tester.scala 31:10]
    phv1_data_108 <= in_port_io_phv_out_data_108; // @[tester.scala 31:10]
    phv1_data_109 <= in_port_io_phv_out_data_109; // @[tester.scala 31:10]
    phv1_data_110 <= in_port_io_phv_out_data_110; // @[tester.scala 31:10]
    phv1_data_111 <= in_port_io_phv_out_data_111; // @[tester.scala 31:10]
    phv1_data_112 <= in_port_io_phv_out_data_112; // @[tester.scala 31:10]
    phv1_data_113 <= in_port_io_phv_out_data_113; // @[tester.scala 31:10]
    phv1_data_114 <= in_port_io_phv_out_data_114; // @[tester.scala 31:10]
    phv1_data_115 <= in_port_io_phv_out_data_115; // @[tester.scala 31:10]
    phv1_data_116 <= in_port_io_phv_out_data_116; // @[tester.scala 31:10]
    phv1_data_117 <= in_port_io_phv_out_data_117; // @[tester.scala 31:10]
    phv1_data_118 <= in_port_io_phv_out_data_118; // @[tester.scala 31:10]
    phv1_data_119 <= in_port_io_phv_out_data_119; // @[tester.scala 31:10]
    phv1_data_120 <= in_port_io_phv_out_data_120; // @[tester.scala 31:10]
    phv1_data_121 <= in_port_io_phv_out_data_121; // @[tester.scala 31:10]
    phv1_data_122 <= in_port_io_phv_out_data_122; // @[tester.scala 31:10]
    phv1_data_123 <= in_port_io_phv_out_data_123; // @[tester.scala 31:10]
    phv1_data_124 <= in_port_io_phv_out_data_124; // @[tester.scala 31:10]
    phv1_data_125 <= in_port_io_phv_out_data_125; // @[tester.scala 31:10]
    phv1_data_126 <= in_port_io_phv_out_data_126; // @[tester.scala 31:10]
    phv1_data_127 <= in_port_io_phv_out_data_127; // @[tester.scala 31:10]
    phv1_valid <= in_port_io_phv_out_valid; // @[tester.scala 31:10]
    phv1_last <= in_port_io_phv_out_last; // @[tester.scala 31:10]
    phv2_data_0 <= phv1_data_0; // @[tester.scala 32:10]
    phv2_data_1 <= phv1_data_1; // @[tester.scala 32:10]
    phv2_data_2 <= phv1_data_2; // @[tester.scala 32:10]
    phv2_data_3 <= phv1_data_3; // @[tester.scala 32:10]
    phv2_data_4 <= phv1_data_4; // @[tester.scala 32:10]
    phv2_data_5 <= phv1_data_5; // @[tester.scala 32:10]
    phv2_data_6 <= phv1_data_6; // @[tester.scala 32:10]
    phv2_data_7 <= phv1_data_7; // @[tester.scala 32:10]
    phv2_data_8 <= phv1_data_8; // @[tester.scala 32:10]
    phv2_data_9 <= phv1_data_9; // @[tester.scala 32:10]
    phv2_data_10 <= phv1_data_10; // @[tester.scala 32:10]
    phv2_data_11 <= phv1_data_11; // @[tester.scala 32:10]
    phv2_data_12 <= phv1_data_12; // @[tester.scala 32:10]
    phv2_data_13 <= phv1_data_13; // @[tester.scala 32:10]
    phv2_data_14 <= phv1_data_14; // @[tester.scala 32:10]
    phv2_data_15 <= phv1_data_15; // @[tester.scala 32:10]
    phv2_data_16 <= phv1_data_16; // @[tester.scala 32:10]
    phv2_data_17 <= phv1_data_17; // @[tester.scala 32:10]
    phv2_data_18 <= phv1_data_18; // @[tester.scala 32:10]
    phv2_data_19 <= phv1_data_19; // @[tester.scala 32:10]
    phv2_data_20 <= phv1_data_20; // @[tester.scala 32:10]
    phv2_data_21 <= phv1_data_21; // @[tester.scala 32:10]
    phv2_data_22 <= phv1_data_22; // @[tester.scala 32:10]
    phv2_data_23 <= phv1_data_23; // @[tester.scala 32:10]
    phv2_data_24 <= phv1_data_24; // @[tester.scala 32:10]
    phv2_data_25 <= phv1_data_25; // @[tester.scala 32:10]
    phv2_data_26 <= phv1_data_26; // @[tester.scala 32:10]
    phv2_data_27 <= phv1_data_27; // @[tester.scala 32:10]
    phv2_data_28 <= phv1_data_28; // @[tester.scala 32:10]
    phv2_data_29 <= phv1_data_29; // @[tester.scala 32:10]
    phv2_data_30 <= phv1_data_30; // @[tester.scala 32:10]
    phv2_data_31 <= phv1_data_31; // @[tester.scala 32:10]
    phv2_data_32 <= phv1_data_32; // @[tester.scala 32:10]
    phv2_data_33 <= phv1_data_33; // @[tester.scala 32:10]
    phv2_data_34 <= phv1_data_34; // @[tester.scala 32:10]
    phv2_data_35 <= phv1_data_35; // @[tester.scala 32:10]
    phv2_data_36 <= phv1_data_36; // @[tester.scala 32:10]
    phv2_data_37 <= phv1_data_37; // @[tester.scala 32:10]
    phv2_data_38 <= phv1_data_38; // @[tester.scala 32:10]
    phv2_data_39 <= phv1_data_39; // @[tester.scala 32:10]
    phv2_data_40 <= phv1_data_40; // @[tester.scala 32:10]
    phv2_data_41 <= phv1_data_41; // @[tester.scala 32:10]
    phv2_data_42 <= phv1_data_42; // @[tester.scala 32:10]
    phv2_data_43 <= phv1_data_43; // @[tester.scala 32:10]
    phv2_data_44 <= phv1_data_44; // @[tester.scala 32:10]
    phv2_data_45 <= phv1_data_45; // @[tester.scala 32:10]
    phv2_data_46 <= phv1_data_46; // @[tester.scala 32:10]
    phv2_data_47 <= phv1_data_47; // @[tester.scala 32:10]
    phv2_data_48 <= phv1_data_48; // @[tester.scala 32:10]
    phv2_data_49 <= phv1_data_49; // @[tester.scala 32:10]
    phv2_data_50 <= phv1_data_50; // @[tester.scala 32:10]
    phv2_data_51 <= phv1_data_51; // @[tester.scala 32:10]
    phv2_data_52 <= phv1_data_52; // @[tester.scala 32:10]
    phv2_data_53 <= phv1_data_53; // @[tester.scala 32:10]
    phv2_data_54 <= phv1_data_54; // @[tester.scala 32:10]
    phv2_data_55 <= phv1_data_55; // @[tester.scala 32:10]
    phv2_data_56 <= phv1_data_56; // @[tester.scala 32:10]
    phv2_data_57 <= phv1_data_57; // @[tester.scala 32:10]
    phv2_data_58 <= phv1_data_58; // @[tester.scala 32:10]
    phv2_data_59 <= phv1_data_59; // @[tester.scala 32:10]
    phv2_data_60 <= phv1_data_60; // @[tester.scala 32:10]
    phv2_data_61 <= phv1_data_61; // @[tester.scala 32:10]
    phv2_data_62 <= phv1_data_62; // @[tester.scala 32:10]
    phv2_data_63 <= phv1_data_63; // @[tester.scala 32:10]
    phv2_data_64 <= phv1_data_64; // @[tester.scala 32:10]
    phv2_data_65 <= phv1_data_65; // @[tester.scala 32:10]
    phv2_data_66 <= phv1_data_66; // @[tester.scala 32:10]
    phv2_data_67 <= phv1_data_67; // @[tester.scala 32:10]
    phv2_data_68 <= phv1_data_68; // @[tester.scala 32:10]
    phv2_data_69 <= phv1_data_69; // @[tester.scala 32:10]
    phv2_data_70 <= phv1_data_70; // @[tester.scala 32:10]
    phv2_data_71 <= phv1_data_71; // @[tester.scala 32:10]
    phv2_data_72 <= phv1_data_72; // @[tester.scala 32:10]
    phv2_data_73 <= phv1_data_73; // @[tester.scala 32:10]
    phv2_data_74 <= phv1_data_74; // @[tester.scala 32:10]
    phv2_data_75 <= phv1_data_75; // @[tester.scala 32:10]
    phv2_data_76 <= phv1_data_76; // @[tester.scala 32:10]
    phv2_data_77 <= phv1_data_77; // @[tester.scala 32:10]
    phv2_data_78 <= phv1_data_78; // @[tester.scala 32:10]
    phv2_data_79 <= phv1_data_79; // @[tester.scala 32:10]
    phv2_data_80 <= phv1_data_80; // @[tester.scala 32:10]
    phv2_data_81 <= phv1_data_81; // @[tester.scala 32:10]
    phv2_data_82 <= phv1_data_82; // @[tester.scala 32:10]
    phv2_data_83 <= phv1_data_83; // @[tester.scala 32:10]
    phv2_data_84 <= phv1_data_84; // @[tester.scala 32:10]
    phv2_data_85 <= phv1_data_85; // @[tester.scala 32:10]
    phv2_data_86 <= phv1_data_86; // @[tester.scala 32:10]
    phv2_data_87 <= phv1_data_87; // @[tester.scala 32:10]
    phv2_data_88 <= phv1_data_88; // @[tester.scala 32:10]
    phv2_data_89 <= phv1_data_89; // @[tester.scala 32:10]
    phv2_data_90 <= phv1_data_90; // @[tester.scala 32:10]
    phv2_data_91 <= phv1_data_91; // @[tester.scala 32:10]
    phv2_data_92 <= phv1_data_92; // @[tester.scala 32:10]
    phv2_data_93 <= phv1_data_93; // @[tester.scala 32:10]
    phv2_data_94 <= phv1_data_94; // @[tester.scala 32:10]
    phv2_data_95 <= phv1_data_95; // @[tester.scala 32:10]
    phv2_data_96 <= phv1_data_96; // @[tester.scala 32:10]
    phv2_data_97 <= phv1_data_97; // @[tester.scala 32:10]
    phv2_data_98 <= phv1_data_98; // @[tester.scala 32:10]
    phv2_data_99 <= phv1_data_99; // @[tester.scala 32:10]
    phv2_data_100 <= phv1_data_100; // @[tester.scala 32:10]
    phv2_data_101 <= phv1_data_101; // @[tester.scala 32:10]
    phv2_data_102 <= phv1_data_102; // @[tester.scala 32:10]
    phv2_data_103 <= phv1_data_103; // @[tester.scala 32:10]
    phv2_data_104 <= phv1_data_104; // @[tester.scala 32:10]
    phv2_data_105 <= phv1_data_105; // @[tester.scala 32:10]
    phv2_data_106 <= phv1_data_106; // @[tester.scala 32:10]
    phv2_data_107 <= phv1_data_107; // @[tester.scala 32:10]
    phv2_data_108 <= phv1_data_108; // @[tester.scala 32:10]
    phv2_data_109 <= phv1_data_109; // @[tester.scala 32:10]
    phv2_data_110 <= phv1_data_110; // @[tester.scala 32:10]
    phv2_data_111 <= phv1_data_111; // @[tester.scala 32:10]
    phv2_data_112 <= phv1_data_112; // @[tester.scala 32:10]
    phv2_data_113 <= phv1_data_113; // @[tester.scala 32:10]
    phv2_data_114 <= phv1_data_114; // @[tester.scala 32:10]
    phv2_data_115 <= phv1_data_115; // @[tester.scala 32:10]
    phv2_data_116 <= phv1_data_116; // @[tester.scala 32:10]
    phv2_data_117 <= phv1_data_117; // @[tester.scala 32:10]
    phv2_data_118 <= phv1_data_118; // @[tester.scala 32:10]
    phv2_data_119 <= phv1_data_119; // @[tester.scala 32:10]
    phv2_data_120 <= phv1_data_120; // @[tester.scala 32:10]
    phv2_data_121 <= phv1_data_121; // @[tester.scala 32:10]
    phv2_data_122 <= phv1_data_122; // @[tester.scala 32:10]
    phv2_data_123 <= phv1_data_123; // @[tester.scala 32:10]
    phv2_data_124 <= phv1_data_124; // @[tester.scala 32:10]
    phv2_data_125 <= phv1_data_125; // @[tester.scala 32:10]
    phv2_data_126 <= phv1_data_126; // @[tester.scala 32:10]
    phv2_data_127 <= phv1_data_127; // @[tester.scala 32:10]
    phv2_valid <= phv1_valid; // @[tester.scala 32:10]
    phv2_last <= phv1_last; // @[tester.scala 32:10]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv1_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv1_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv1_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv1_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv1_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv1_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv1_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv1_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv1_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv1_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv1_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv1_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv1_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv1_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv1_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv1_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv1_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv1_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv1_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv1_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv1_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv1_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv1_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv1_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv1_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv1_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv1_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv1_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv1_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv1_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv1_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv1_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv1_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv1_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv1_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv1_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv1_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv1_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv1_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv1_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv1_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv1_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv1_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv1_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv1_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv1_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv1_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv1_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv1_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv1_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv1_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv1_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv1_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv1_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv1_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv1_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv1_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv1_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv1_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv1_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv1_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv1_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv1_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv1_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv1_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv1_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv1_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv1_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv1_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv1_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv1_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv1_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv1_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv1_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv1_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv1_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv1_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv1_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv1_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv1_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv1_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv1_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv1_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv1_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv1_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv1_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv1_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv1_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv1_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv1_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv1_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv1_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv1_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv1_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv1_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv1_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv1_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv1_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv1_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv1_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv1_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv1_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv1_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv1_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv1_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv1_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv1_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv1_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv1_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv1_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv1_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv1_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv1_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv1_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv1_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv1_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv1_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv1_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv1_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv1_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv1_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv1_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv1_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv1_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv1_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv1_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv1_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv1_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv1_valid = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  phv1_last = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  phv2_data_0 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv2_data_1 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv2_data_2 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv2_data_3 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv2_data_4 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv2_data_5 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv2_data_6 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv2_data_7 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv2_data_8 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv2_data_9 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv2_data_10 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv2_data_11 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv2_data_12 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv2_data_13 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv2_data_14 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv2_data_15 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv2_data_16 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv2_data_17 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv2_data_18 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv2_data_19 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv2_data_20 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv2_data_21 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv2_data_22 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv2_data_23 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv2_data_24 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv2_data_25 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv2_data_26 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv2_data_27 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv2_data_28 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv2_data_29 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv2_data_30 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  phv2_data_31 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  phv2_data_32 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  phv2_data_33 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  phv2_data_34 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  phv2_data_35 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  phv2_data_36 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  phv2_data_37 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  phv2_data_38 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  phv2_data_39 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  phv2_data_40 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  phv2_data_41 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  phv2_data_42 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  phv2_data_43 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  phv2_data_44 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  phv2_data_45 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  phv2_data_46 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv2_data_47 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv2_data_48 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  phv2_data_49 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  phv2_data_50 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  phv2_data_51 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  phv2_data_52 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  phv2_data_53 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  phv2_data_54 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  phv2_data_55 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  phv2_data_56 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  phv2_data_57 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  phv2_data_58 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  phv2_data_59 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  phv2_data_60 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  phv2_data_61 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  phv2_data_62 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  phv2_data_63 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  phv2_data_64 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  phv2_data_65 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  phv2_data_66 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  phv2_data_67 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  phv2_data_68 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  phv2_data_69 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  phv2_data_70 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  phv2_data_71 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  phv2_data_72 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  phv2_data_73 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  phv2_data_74 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  phv2_data_75 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  phv2_data_76 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  phv2_data_77 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  phv2_data_78 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  phv2_data_79 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  phv2_data_80 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  phv2_data_81 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  phv2_data_82 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  phv2_data_83 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  phv2_data_84 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  phv2_data_85 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  phv2_data_86 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  phv2_data_87 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  phv2_data_88 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  phv2_data_89 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  phv2_data_90 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  phv2_data_91 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  phv2_data_92 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  phv2_data_93 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  phv2_data_94 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  phv2_data_95 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  phv2_data_96 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  phv2_data_97 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  phv2_data_98 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  phv2_data_99 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  phv2_data_100 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  phv2_data_101 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  phv2_data_102 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  phv2_data_103 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  phv2_data_104 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  phv2_data_105 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  phv2_data_106 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  phv2_data_107 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  phv2_data_108 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  phv2_data_109 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  phv2_data_110 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  phv2_data_111 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  phv2_data_112 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  phv2_data_113 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  phv2_data_114 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  phv2_data_115 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  phv2_data_116 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  phv2_data_117 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  phv2_data_118 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  phv2_data_119 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  phv2_data_120 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  phv2_data_121 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  phv2_data_122 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  phv2_data_123 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  phv2_data_124 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  phv2_data_125 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  phv2_data_126 = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  phv2_data_127 = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  phv2_valid = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  phv2_last = _RAND_259[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
