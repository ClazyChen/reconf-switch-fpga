module Matcher(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [7:0]  io_pipe_phv_in_data_256,
  input  [7:0]  io_pipe_phv_in_data_257,
  input  [7:0]  io_pipe_phv_in_data_258,
  input  [7:0]  io_pipe_phv_in_data_259,
  input  [7:0]  io_pipe_phv_in_data_260,
  input  [7:0]  io_pipe_phv_in_data_261,
  input  [7:0]  io_pipe_phv_in_data_262,
  input  [7:0]  io_pipe_phv_in_data_263,
  input  [7:0]  io_pipe_phv_in_data_264,
  input  [7:0]  io_pipe_phv_in_data_265,
  input  [7:0]  io_pipe_phv_in_data_266,
  input  [7:0]  io_pipe_phv_in_data_267,
  input  [7:0]  io_pipe_phv_in_data_268,
  input  [7:0]  io_pipe_phv_in_data_269,
  input  [7:0]  io_pipe_phv_in_data_270,
  input  [7:0]  io_pipe_phv_in_data_271,
  input  [7:0]  io_pipe_phv_in_data_272,
  input  [7:0]  io_pipe_phv_in_data_273,
  input  [7:0]  io_pipe_phv_in_data_274,
  input  [7:0]  io_pipe_phv_in_data_275,
  input  [7:0]  io_pipe_phv_in_data_276,
  input  [7:0]  io_pipe_phv_in_data_277,
  input  [7:0]  io_pipe_phv_in_data_278,
  input  [7:0]  io_pipe_phv_in_data_279,
  input  [7:0]  io_pipe_phv_in_data_280,
  input  [7:0]  io_pipe_phv_in_data_281,
  input  [7:0]  io_pipe_phv_in_data_282,
  input  [7:0]  io_pipe_phv_in_data_283,
  input  [7:0]  io_pipe_phv_in_data_284,
  input  [7:0]  io_pipe_phv_in_data_285,
  input  [7:0]  io_pipe_phv_in_data_286,
  input  [7:0]  io_pipe_phv_in_data_287,
  input  [7:0]  io_pipe_phv_in_data_288,
  input  [7:0]  io_pipe_phv_in_data_289,
  input  [7:0]  io_pipe_phv_in_data_290,
  input  [7:0]  io_pipe_phv_in_data_291,
  input  [7:0]  io_pipe_phv_in_data_292,
  input  [7:0]  io_pipe_phv_in_data_293,
  input  [7:0]  io_pipe_phv_in_data_294,
  input  [7:0]  io_pipe_phv_in_data_295,
  input  [7:0]  io_pipe_phv_in_data_296,
  input  [7:0]  io_pipe_phv_in_data_297,
  input  [7:0]  io_pipe_phv_in_data_298,
  input  [7:0]  io_pipe_phv_in_data_299,
  input  [7:0]  io_pipe_phv_in_data_300,
  input  [7:0]  io_pipe_phv_in_data_301,
  input  [7:0]  io_pipe_phv_in_data_302,
  input  [7:0]  io_pipe_phv_in_data_303,
  input  [7:0]  io_pipe_phv_in_data_304,
  input  [7:0]  io_pipe_phv_in_data_305,
  input  [7:0]  io_pipe_phv_in_data_306,
  input  [7:0]  io_pipe_phv_in_data_307,
  input  [7:0]  io_pipe_phv_in_data_308,
  input  [7:0]  io_pipe_phv_in_data_309,
  input  [7:0]  io_pipe_phv_in_data_310,
  input  [7:0]  io_pipe_phv_in_data_311,
  input  [7:0]  io_pipe_phv_in_data_312,
  input  [7:0]  io_pipe_phv_in_data_313,
  input  [7:0]  io_pipe_phv_in_data_314,
  input  [7:0]  io_pipe_phv_in_data_315,
  input  [7:0]  io_pipe_phv_in_data_316,
  input  [7:0]  io_pipe_phv_in_data_317,
  input  [7:0]  io_pipe_phv_in_data_318,
  input  [7:0]  io_pipe_phv_in_data_319,
  input  [7:0]  io_pipe_phv_in_data_320,
  input  [7:0]  io_pipe_phv_in_data_321,
  input  [7:0]  io_pipe_phv_in_data_322,
  input  [7:0]  io_pipe_phv_in_data_323,
  input  [7:0]  io_pipe_phv_in_data_324,
  input  [7:0]  io_pipe_phv_in_data_325,
  input  [7:0]  io_pipe_phv_in_data_326,
  input  [7:0]  io_pipe_phv_in_data_327,
  input  [7:0]  io_pipe_phv_in_data_328,
  input  [7:0]  io_pipe_phv_in_data_329,
  input  [7:0]  io_pipe_phv_in_data_330,
  input  [7:0]  io_pipe_phv_in_data_331,
  input  [7:0]  io_pipe_phv_in_data_332,
  input  [7:0]  io_pipe_phv_in_data_333,
  input  [7:0]  io_pipe_phv_in_data_334,
  input  [7:0]  io_pipe_phv_in_data_335,
  input  [7:0]  io_pipe_phv_in_data_336,
  input  [7:0]  io_pipe_phv_in_data_337,
  input  [7:0]  io_pipe_phv_in_data_338,
  input  [7:0]  io_pipe_phv_in_data_339,
  input  [7:0]  io_pipe_phv_in_data_340,
  input  [7:0]  io_pipe_phv_in_data_341,
  input  [7:0]  io_pipe_phv_in_data_342,
  input  [7:0]  io_pipe_phv_in_data_343,
  input  [7:0]  io_pipe_phv_in_data_344,
  input  [7:0]  io_pipe_phv_in_data_345,
  input  [7:0]  io_pipe_phv_in_data_346,
  input  [7:0]  io_pipe_phv_in_data_347,
  input  [7:0]  io_pipe_phv_in_data_348,
  input  [7:0]  io_pipe_phv_in_data_349,
  input  [7:0]  io_pipe_phv_in_data_350,
  input  [7:0]  io_pipe_phv_in_data_351,
  input  [7:0]  io_pipe_phv_in_data_352,
  input  [7:0]  io_pipe_phv_in_data_353,
  input  [7:0]  io_pipe_phv_in_data_354,
  input  [7:0]  io_pipe_phv_in_data_355,
  input  [7:0]  io_pipe_phv_in_data_356,
  input  [7:0]  io_pipe_phv_in_data_357,
  input  [7:0]  io_pipe_phv_in_data_358,
  input  [7:0]  io_pipe_phv_in_data_359,
  input  [7:0]  io_pipe_phv_in_data_360,
  input  [7:0]  io_pipe_phv_in_data_361,
  input  [7:0]  io_pipe_phv_in_data_362,
  input  [7:0]  io_pipe_phv_in_data_363,
  input  [7:0]  io_pipe_phv_in_data_364,
  input  [7:0]  io_pipe_phv_in_data_365,
  input  [7:0]  io_pipe_phv_in_data_366,
  input  [7:0]  io_pipe_phv_in_data_367,
  input  [7:0]  io_pipe_phv_in_data_368,
  input  [7:0]  io_pipe_phv_in_data_369,
  input  [7:0]  io_pipe_phv_in_data_370,
  input  [7:0]  io_pipe_phv_in_data_371,
  input  [7:0]  io_pipe_phv_in_data_372,
  input  [7:0]  io_pipe_phv_in_data_373,
  input  [7:0]  io_pipe_phv_in_data_374,
  input  [7:0]  io_pipe_phv_in_data_375,
  input  [7:0]  io_pipe_phv_in_data_376,
  input  [7:0]  io_pipe_phv_in_data_377,
  input  [7:0]  io_pipe_phv_in_data_378,
  input  [7:0]  io_pipe_phv_in_data_379,
  input  [7:0]  io_pipe_phv_in_data_380,
  input  [7:0]  io_pipe_phv_in_data_381,
  input  [7:0]  io_pipe_phv_in_data_382,
  input  [7:0]  io_pipe_phv_in_data_383,
  input  [7:0]  io_pipe_phv_in_data_384,
  input  [7:0]  io_pipe_phv_in_data_385,
  input  [7:0]  io_pipe_phv_in_data_386,
  input  [7:0]  io_pipe_phv_in_data_387,
  input  [7:0]  io_pipe_phv_in_data_388,
  input  [7:0]  io_pipe_phv_in_data_389,
  input  [7:0]  io_pipe_phv_in_data_390,
  input  [7:0]  io_pipe_phv_in_data_391,
  input  [7:0]  io_pipe_phv_in_data_392,
  input  [7:0]  io_pipe_phv_in_data_393,
  input  [7:0]  io_pipe_phv_in_data_394,
  input  [7:0]  io_pipe_phv_in_data_395,
  input  [7:0]  io_pipe_phv_in_data_396,
  input  [7:0]  io_pipe_phv_in_data_397,
  input  [7:0]  io_pipe_phv_in_data_398,
  input  [7:0]  io_pipe_phv_in_data_399,
  input  [7:0]  io_pipe_phv_in_data_400,
  input  [7:0]  io_pipe_phv_in_data_401,
  input  [7:0]  io_pipe_phv_in_data_402,
  input  [7:0]  io_pipe_phv_in_data_403,
  input  [7:0]  io_pipe_phv_in_data_404,
  input  [7:0]  io_pipe_phv_in_data_405,
  input  [7:0]  io_pipe_phv_in_data_406,
  input  [7:0]  io_pipe_phv_in_data_407,
  input  [7:0]  io_pipe_phv_in_data_408,
  input  [7:0]  io_pipe_phv_in_data_409,
  input  [7:0]  io_pipe_phv_in_data_410,
  input  [7:0]  io_pipe_phv_in_data_411,
  input  [7:0]  io_pipe_phv_in_data_412,
  input  [7:0]  io_pipe_phv_in_data_413,
  input  [7:0]  io_pipe_phv_in_data_414,
  input  [7:0]  io_pipe_phv_in_data_415,
  input  [7:0]  io_pipe_phv_in_data_416,
  input  [7:0]  io_pipe_phv_in_data_417,
  input  [7:0]  io_pipe_phv_in_data_418,
  input  [7:0]  io_pipe_phv_in_data_419,
  input  [7:0]  io_pipe_phv_in_data_420,
  input  [7:0]  io_pipe_phv_in_data_421,
  input  [7:0]  io_pipe_phv_in_data_422,
  input  [7:0]  io_pipe_phv_in_data_423,
  input  [7:0]  io_pipe_phv_in_data_424,
  input  [7:0]  io_pipe_phv_in_data_425,
  input  [7:0]  io_pipe_phv_in_data_426,
  input  [7:0]  io_pipe_phv_in_data_427,
  input  [7:0]  io_pipe_phv_in_data_428,
  input  [7:0]  io_pipe_phv_in_data_429,
  input  [7:0]  io_pipe_phv_in_data_430,
  input  [7:0]  io_pipe_phv_in_data_431,
  input  [7:0]  io_pipe_phv_in_data_432,
  input  [7:0]  io_pipe_phv_in_data_433,
  input  [7:0]  io_pipe_phv_in_data_434,
  input  [7:0]  io_pipe_phv_in_data_435,
  input  [7:0]  io_pipe_phv_in_data_436,
  input  [7:0]  io_pipe_phv_in_data_437,
  input  [7:0]  io_pipe_phv_in_data_438,
  input  [7:0]  io_pipe_phv_in_data_439,
  input  [7:0]  io_pipe_phv_in_data_440,
  input  [7:0]  io_pipe_phv_in_data_441,
  input  [7:0]  io_pipe_phv_in_data_442,
  input  [7:0]  io_pipe_phv_in_data_443,
  input  [7:0]  io_pipe_phv_in_data_444,
  input  [7:0]  io_pipe_phv_in_data_445,
  input  [7:0]  io_pipe_phv_in_data_446,
  input  [7:0]  io_pipe_phv_in_data_447,
  input  [7:0]  io_pipe_phv_in_data_448,
  input  [7:0]  io_pipe_phv_in_data_449,
  input  [7:0]  io_pipe_phv_in_data_450,
  input  [7:0]  io_pipe_phv_in_data_451,
  input  [7:0]  io_pipe_phv_in_data_452,
  input  [7:0]  io_pipe_phv_in_data_453,
  input  [7:0]  io_pipe_phv_in_data_454,
  input  [7:0]  io_pipe_phv_in_data_455,
  input  [7:0]  io_pipe_phv_in_data_456,
  input  [7:0]  io_pipe_phv_in_data_457,
  input  [7:0]  io_pipe_phv_in_data_458,
  input  [7:0]  io_pipe_phv_in_data_459,
  input  [7:0]  io_pipe_phv_in_data_460,
  input  [7:0]  io_pipe_phv_in_data_461,
  input  [7:0]  io_pipe_phv_in_data_462,
  input  [7:0]  io_pipe_phv_in_data_463,
  input  [7:0]  io_pipe_phv_in_data_464,
  input  [7:0]  io_pipe_phv_in_data_465,
  input  [7:0]  io_pipe_phv_in_data_466,
  input  [7:0]  io_pipe_phv_in_data_467,
  input  [7:0]  io_pipe_phv_in_data_468,
  input  [7:0]  io_pipe_phv_in_data_469,
  input  [7:0]  io_pipe_phv_in_data_470,
  input  [7:0]  io_pipe_phv_in_data_471,
  input  [7:0]  io_pipe_phv_in_data_472,
  input  [7:0]  io_pipe_phv_in_data_473,
  input  [7:0]  io_pipe_phv_in_data_474,
  input  [7:0]  io_pipe_phv_in_data_475,
  input  [7:0]  io_pipe_phv_in_data_476,
  input  [7:0]  io_pipe_phv_in_data_477,
  input  [7:0]  io_pipe_phv_in_data_478,
  input  [7:0]  io_pipe_phv_in_data_479,
  input  [7:0]  io_pipe_phv_in_data_480,
  input  [7:0]  io_pipe_phv_in_data_481,
  input  [7:0]  io_pipe_phv_in_data_482,
  input  [7:0]  io_pipe_phv_in_data_483,
  input  [7:0]  io_pipe_phv_in_data_484,
  input  [7:0]  io_pipe_phv_in_data_485,
  input  [7:0]  io_pipe_phv_in_data_486,
  input  [7:0]  io_pipe_phv_in_data_487,
  input  [7:0]  io_pipe_phv_in_data_488,
  input  [7:0]  io_pipe_phv_in_data_489,
  input  [7:0]  io_pipe_phv_in_data_490,
  input  [7:0]  io_pipe_phv_in_data_491,
  input  [7:0]  io_pipe_phv_in_data_492,
  input  [7:0]  io_pipe_phv_in_data_493,
  input  [7:0]  io_pipe_phv_in_data_494,
  input  [7:0]  io_pipe_phv_in_data_495,
  input  [7:0]  io_pipe_phv_in_data_496,
  input  [7:0]  io_pipe_phv_in_data_497,
  input  [7:0]  io_pipe_phv_in_data_498,
  input  [7:0]  io_pipe_phv_in_data_499,
  input  [7:0]  io_pipe_phv_in_data_500,
  input  [7:0]  io_pipe_phv_in_data_501,
  input  [7:0]  io_pipe_phv_in_data_502,
  input  [7:0]  io_pipe_phv_in_data_503,
  input  [7:0]  io_pipe_phv_in_data_504,
  input  [7:0]  io_pipe_phv_in_data_505,
  input  [7:0]  io_pipe_phv_in_data_506,
  input  [7:0]  io_pipe_phv_in_data_507,
  input  [7:0]  io_pipe_phv_in_data_508,
  input  [7:0]  io_pipe_phv_in_data_509,
  input  [7:0]  io_pipe_phv_in_data_510,
  input  [7:0]  io_pipe_phv_in_data_511,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [7:0]  io_pipe_phv_out_data_256,
  output [7:0]  io_pipe_phv_out_data_257,
  output [7:0]  io_pipe_phv_out_data_258,
  output [7:0]  io_pipe_phv_out_data_259,
  output [7:0]  io_pipe_phv_out_data_260,
  output [7:0]  io_pipe_phv_out_data_261,
  output [7:0]  io_pipe_phv_out_data_262,
  output [7:0]  io_pipe_phv_out_data_263,
  output [7:0]  io_pipe_phv_out_data_264,
  output [7:0]  io_pipe_phv_out_data_265,
  output [7:0]  io_pipe_phv_out_data_266,
  output [7:0]  io_pipe_phv_out_data_267,
  output [7:0]  io_pipe_phv_out_data_268,
  output [7:0]  io_pipe_phv_out_data_269,
  output [7:0]  io_pipe_phv_out_data_270,
  output [7:0]  io_pipe_phv_out_data_271,
  output [7:0]  io_pipe_phv_out_data_272,
  output [7:0]  io_pipe_phv_out_data_273,
  output [7:0]  io_pipe_phv_out_data_274,
  output [7:0]  io_pipe_phv_out_data_275,
  output [7:0]  io_pipe_phv_out_data_276,
  output [7:0]  io_pipe_phv_out_data_277,
  output [7:0]  io_pipe_phv_out_data_278,
  output [7:0]  io_pipe_phv_out_data_279,
  output [7:0]  io_pipe_phv_out_data_280,
  output [7:0]  io_pipe_phv_out_data_281,
  output [7:0]  io_pipe_phv_out_data_282,
  output [7:0]  io_pipe_phv_out_data_283,
  output [7:0]  io_pipe_phv_out_data_284,
  output [7:0]  io_pipe_phv_out_data_285,
  output [7:0]  io_pipe_phv_out_data_286,
  output [7:0]  io_pipe_phv_out_data_287,
  output [7:0]  io_pipe_phv_out_data_288,
  output [7:0]  io_pipe_phv_out_data_289,
  output [7:0]  io_pipe_phv_out_data_290,
  output [7:0]  io_pipe_phv_out_data_291,
  output [7:0]  io_pipe_phv_out_data_292,
  output [7:0]  io_pipe_phv_out_data_293,
  output [7:0]  io_pipe_phv_out_data_294,
  output [7:0]  io_pipe_phv_out_data_295,
  output [7:0]  io_pipe_phv_out_data_296,
  output [7:0]  io_pipe_phv_out_data_297,
  output [7:0]  io_pipe_phv_out_data_298,
  output [7:0]  io_pipe_phv_out_data_299,
  output [7:0]  io_pipe_phv_out_data_300,
  output [7:0]  io_pipe_phv_out_data_301,
  output [7:0]  io_pipe_phv_out_data_302,
  output [7:0]  io_pipe_phv_out_data_303,
  output [7:0]  io_pipe_phv_out_data_304,
  output [7:0]  io_pipe_phv_out_data_305,
  output [7:0]  io_pipe_phv_out_data_306,
  output [7:0]  io_pipe_phv_out_data_307,
  output [7:0]  io_pipe_phv_out_data_308,
  output [7:0]  io_pipe_phv_out_data_309,
  output [7:0]  io_pipe_phv_out_data_310,
  output [7:0]  io_pipe_phv_out_data_311,
  output [7:0]  io_pipe_phv_out_data_312,
  output [7:0]  io_pipe_phv_out_data_313,
  output [7:0]  io_pipe_phv_out_data_314,
  output [7:0]  io_pipe_phv_out_data_315,
  output [7:0]  io_pipe_phv_out_data_316,
  output [7:0]  io_pipe_phv_out_data_317,
  output [7:0]  io_pipe_phv_out_data_318,
  output [7:0]  io_pipe_phv_out_data_319,
  output [7:0]  io_pipe_phv_out_data_320,
  output [7:0]  io_pipe_phv_out_data_321,
  output [7:0]  io_pipe_phv_out_data_322,
  output [7:0]  io_pipe_phv_out_data_323,
  output [7:0]  io_pipe_phv_out_data_324,
  output [7:0]  io_pipe_phv_out_data_325,
  output [7:0]  io_pipe_phv_out_data_326,
  output [7:0]  io_pipe_phv_out_data_327,
  output [7:0]  io_pipe_phv_out_data_328,
  output [7:0]  io_pipe_phv_out_data_329,
  output [7:0]  io_pipe_phv_out_data_330,
  output [7:0]  io_pipe_phv_out_data_331,
  output [7:0]  io_pipe_phv_out_data_332,
  output [7:0]  io_pipe_phv_out_data_333,
  output [7:0]  io_pipe_phv_out_data_334,
  output [7:0]  io_pipe_phv_out_data_335,
  output [7:0]  io_pipe_phv_out_data_336,
  output [7:0]  io_pipe_phv_out_data_337,
  output [7:0]  io_pipe_phv_out_data_338,
  output [7:0]  io_pipe_phv_out_data_339,
  output [7:0]  io_pipe_phv_out_data_340,
  output [7:0]  io_pipe_phv_out_data_341,
  output [7:0]  io_pipe_phv_out_data_342,
  output [7:0]  io_pipe_phv_out_data_343,
  output [7:0]  io_pipe_phv_out_data_344,
  output [7:0]  io_pipe_phv_out_data_345,
  output [7:0]  io_pipe_phv_out_data_346,
  output [7:0]  io_pipe_phv_out_data_347,
  output [7:0]  io_pipe_phv_out_data_348,
  output [7:0]  io_pipe_phv_out_data_349,
  output [7:0]  io_pipe_phv_out_data_350,
  output [7:0]  io_pipe_phv_out_data_351,
  output [7:0]  io_pipe_phv_out_data_352,
  output [7:0]  io_pipe_phv_out_data_353,
  output [7:0]  io_pipe_phv_out_data_354,
  output [7:0]  io_pipe_phv_out_data_355,
  output [7:0]  io_pipe_phv_out_data_356,
  output [7:0]  io_pipe_phv_out_data_357,
  output [7:0]  io_pipe_phv_out_data_358,
  output [7:0]  io_pipe_phv_out_data_359,
  output [7:0]  io_pipe_phv_out_data_360,
  output [7:0]  io_pipe_phv_out_data_361,
  output [7:0]  io_pipe_phv_out_data_362,
  output [7:0]  io_pipe_phv_out_data_363,
  output [7:0]  io_pipe_phv_out_data_364,
  output [7:0]  io_pipe_phv_out_data_365,
  output [7:0]  io_pipe_phv_out_data_366,
  output [7:0]  io_pipe_phv_out_data_367,
  output [7:0]  io_pipe_phv_out_data_368,
  output [7:0]  io_pipe_phv_out_data_369,
  output [7:0]  io_pipe_phv_out_data_370,
  output [7:0]  io_pipe_phv_out_data_371,
  output [7:0]  io_pipe_phv_out_data_372,
  output [7:0]  io_pipe_phv_out_data_373,
  output [7:0]  io_pipe_phv_out_data_374,
  output [7:0]  io_pipe_phv_out_data_375,
  output [7:0]  io_pipe_phv_out_data_376,
  output [7:0]  io_pipe_phv_out_data_377,
  output [7:0]  io_pipe_phv_out_data_378,
  output [7:0]  io_pipe_phv_out_data_379,
  output [7:0]  io_pipe_phv_out_data_380,
  output [7:0]  io_pipe_phv_out_data_381,
  output [7:0]  io_pipe_phv_out_data_382,
  output [7:0]  io_pipe_phv_out_data_383,
  output [7:0]  io_pipe_phv_out_data_384,
  output [7:0]  io_pipe_phv_out_data_385,
  output [7:0]  io_pipe_phv_out_data_386,
  output [7:0]  io_pipe_phv_out_data_387,
  output [7:0]  io_pipe_phv_out_data_388,
  output [7:0]  io_pipe_phv_out_data_389,
  output [7:0]  io_pipe_phv_out_data_390,
  output [7:0]  io_pipe_phv_out_data_391,
  output [7:0]  io_pipe_phv_out_data_392,
  output [7:0]  io_pipe_phv_out_data_393,
  output [7:0]  io_pipe_phv_out_data_394,
  output [7:0]  io_pipe_phv_out_data_395,
  output [7:0]  io_pipe_phv_out_data_396,
  output [7:0]  io_pipe_phv_out_data_397,
  output [7:0]  io_pipe_phv_out_data_398,
  output [7:0]  io_pipe_phv_out_data_399,
  output [7:0]  io_pipe_phv_out_data_400,
  output [7:0]  io_pipe_phv_out_data_401,
  output [7:0]  io_pipe_phv_out_data_402,
  output [7:0]  io_pipe_phv_out_data_403,
  output [7:0]  io_pipe_phv_out_data_404,
  output [7:0]  io_pipe_phv_out_data_405,
  output [7:0]  io_pipe_phv_out_data_406,
  output [7:0]  io_pipe_phv_out_data_407,
  output [7:0]  io_pipe_phv_out_data_408,
  output [7:0]  io_pipe_phv_out_data_409,
  output [7:0]  io_pipe_phv_out_data_410,
  output [7:0]  io_pipe_phv_out_data_411,
  output [7:0]  io_pipe_phv_out_data_412,
  output [7:0]  io_pipe_phv_out_data_413,
  output [7:0]  io_pipe_phv_out_data_414,
  output [7:0]  io_pipe_phv_out_data_415,
  output [7:0]  io_pipe_phv_out_data_416,
  output [7:0]  io_pipe_phv_out_data_417,
  output [7:0]  io_pipe_phv_out_data_418,
  output [7:0]  io_pipe_phv_out_data_419,
  output [7:0]  io_pipe_phv_out_data_420,
  output [7:0]  io_pipe_phv_out_data_421,
  output [7:0]  io_pipe_phv_out_data_422,
  output [7:0]  io_pipe_phv_out_data_423,
  output [7:0]  io_pipe_phv_out_data_424,
  output [7:0]  io_pipe_phv_out_data_425,
  output [7:0]  io_pipe_phv_out_data_426,
  output [7:0]  io_pipe_phv_out_data_427,
  output [7:0]  io_pipe_phv_out_data_428,
  output [7:0]  io_pipe_phv_out_data_429,
  output [7:0]  io_pipe_phv_out_data_430,
  output [7:0]  io_pipe_phv_out_data_431,
  output [7:0]  io_pipe_phv_out_data_432,
  output [7:0]  io_pipe_phv_out_data_433,
  output [7:0]  io_pipe_phv_out_data_434,
  output [7:0]  io_pipe_phv_out_data_435,
  output [7:0]  io_pipe_phv_out_data_436,
  output [7:0]  io_pipe_phv_out_data_437,
  output [7:0]  io_pipe_phv_out_data_438,
  output [7:0]  io_pipe_phv_out_data_439,
  output [7:0]  io_pipe_phv_out_data_440,
  output [7:0]  io_pipe_phv_out_data_441,
  output [7:0]  io_pipe_phv_out_data_442,
  output [7:0]  io_pipe_phv_out_data_443,
  output [7:0]  io_pipe_phv_out_data_444,
  output [7:0]  io_pipe_phv_out_data_445,
  output [7:0]  io_pipe_phv_out_data_446,
  output [7:0]  io_pipe_phv_out_data_447,
  output [7:0]  io_pipe_phv_out_data_448,
  output [7:0]  io_pipe_phv_out_data_449,
  output [7:0]  io_pipe_phv_out_data_450,
  output [7:0]  io_pipe_phv_out_data_451,
  output [7:0]  io_pipe_phv_out_data_452,
  output [7:0]  io_pipe_phv_out_data_453,
  output [7:0]  io_pipe_phv_out_data_454,
  output [7:0]  io_pipe_phv_out_data_455,
  output [7:0]  io_pipe_phv_out_data_456,
  output [7:0]  io_pipe_phv_out_data_457,
  output [7:0]  io_pipe_phv_out_data_458,
  output [7:0]  io_pipe_phv_out_data_459,
  output [7:0]  io_pipe_phv_out_data_460,
  output [7:0]  io_pipe_phv_out_data_461,
  output [7:0]  io_pipe_phv_out_data_462,
  output [7:0]  io_pipe_phv_out_data_463,
  output [7:0]  io_pipe_phv_out_data_464,
  output [7:0]  io_pipe_phv_out_data_465,
  output [7:0]  io_pipe_phv_out_data_466,
  output [7:0]  io_pipe_phv_out_data_467,
  output [7:0]  io_pipe_phv_out_data_468,
  output [7:0]  io_pipe_phv_out_data_469,
  output [7:0]  io_pipe_phv_out_data_470,
  output [7:0]  io_pipe_phv_out_data_471,
  output [7:0]  io_pipe_phv_out_data_472,
  output [7:0]  io_pipe_phv_out_data_473,
  output [7:0]  io_pipe_phv_out_data_474,
  output [7:0]  io_pipe_phv_out_data_475,
  output [7:0]  io_pipe_phv_out_data_476,
  output [7:0]  io_pipe_phv_out_data_477,
  output [7:0]  io_pipe_phv_out_data_478,
  output [7:0]  io_pipe_phv_out_data_479,
  output [7:0]  io_pipe_phv_out_data_480,
  output [7:0]  io_pipe_phv_out_data_481,
  output [7:0]  io_pipe_phv_out_data_482,
  output [7:0]  io_pipe_phv_out_data_483,
  output [7:0]  io_pipe_phv_out_data_484,
  output [7:0]  io_pipe_phv_out_data_485,
  output [7:0]  io_pipe_phv_out_data_486,
  output [7:0]  io_pipe_phv_out_data_487,
  output [7:0]  io_pipe_phv_out_data_488,
  output [7:0]  io_pipe_phv_out_data_489,
  output [7:0]  io_pipe_phv_out_data_490,
  output [7:0]  io_pipe_phv_out_data_491,
  output [7:0]  io_pipe_phv_out_data_492,
  output [7:0]  io_pipe_phv_out_data_493,
  output [7:0]  io_pipe_phv_out_data_494,
  output [7:0]  io_pipe_phv_out_data_495,
  output [7:0]  io_pipe_phv_out_data_496,
  output [7:0]  io_pipe_phv_out_data_497,
  output [7:0]  io_pipe_phv_out_data_498,
  output [7:0]  io_pipe_phv_out_data_499,
  output [7:0]  io_pipe_phv_out_data_500,
  output [7:0]  io_pipe_phv_out_data_501,
  output [7:0]  io_pipe_phv_out_data_502,
  output [7:0]  io_pipe_phv_out_data_503,
  output [7:0]  io_pipe_phv_out_data_504,
  output [7:0]  io_pipe_phv_out_data_505,
  output [7:0]  io_pipe_phv_out_data_506,
  output [7:0]  io_pipe_phv_out_data_507,
  output [7:0]  io_pipe_phv_out_data_508,
  output [7:0]  io_pipe_phv_out_data_509,
  output [7:0]  io_pipe_phv_out_data_510,
  output [7:0]  io_pipe_phv_out_data_511,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input         io_mod_en,
  input         io_mod_config_id,
  input  [7:0]  io_mod_key_mod_header_id,
  input  [7:0]  io_mod_key_mod_internal_offset,
  input  [7:0]  io_mod_key_mod_key_length,
  input  [4:0]  io_mod_table_mod_table_width,
  input  [4:0]  io_mod_table_mod_table_depth,
  output        io_hit,
  output [63:0] io_match_value,
  output        io_mem_cluster_0_en,
  output [7:0]  io_mem_cluster_0_addr,
  input  [63:0] io_mem_cluster_0_data,
  output        io_mem_cluster_1_en,
  output [7:0]  io_mem_cluster_1_addr,
  input  [63:0] io_mem_cluster_1_data,
  output        io_mem_cluster_2_en,
  output [7:0]  io_mem_cluster_2_addr,
  input  [63:0] io_mem_cluster_2_data,
  output        io_mem_cluster_3_en,
  output [7:0]  io_mem_cluster_3_addr,
  input  [63:0] io_mem_cluster_3_data,
  output        io_mem_cluster_4_en,
  output [7:0]  io_mem_cluster_4_addr,
  input  [63:0] io_mem_cluster_4_data,
  output        io_mem_cluster_5_en,
  output [7:0]  io_mem_cluster_5_addr,
  input  [63:0] io_mem_cluster_5_data,
  output        io_mem_cluster_6_en,
  output [7:0]  io_mem_cluster_6_addr,
  input  [63:0] io_mem_cluster_6_data,
  output        io_mem_cluster_7_en,
  output [7:0]  io_mem_cluster_7_addr,
  input  [63:0] io_mem_cluster_7_data,
  output        io_mem_cluster_8_en,
  output [7:0]  io_mem_cluster_8_addr,
  input  [63:0] io_mem_cluster_8_data,
  output        io_mem_cluster_9_en,
  output [7:0]  io_mem_cluster_9_addr,
  input  [63:0] io_mem_cluster_9_data,
  output        io_mem_cluster_10_en,
  output [7:0]  io_mem_cluster_10_addr,
  input  [63:0] io_mem_cluster_10_data,
  output        io_mem_cluster_11_en,
  output [7:0]  io_mem_cluster_11_addr,
  input  [63:0] io_mem_cluster_11_data,
  output        io_mem_cluster_12_en,
  output [7:0]  io_mem_cluster_12_addr,
  input  [63:0] io_mem_cluster_12_data,
  output        io_mem_cluster_13_en,
  output [7:0]  io_mem_cluster_13_addr,
  input  [63:0] io_mem_cluster_13_data,
  output        io_mem_cluster_14_en,
  output [7:0]  io_mem_cluster_14_addr,
  input  [63:0] io_mem_cluster_14_data,
  output        io_mem_cluster_15_en,
  output [7:0]  io_mem_cluster_15_addr,
  input  [63:0] io_mem_cluster_15_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  pipe1_clock; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_0; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_1; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_2; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_3; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_4; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_5; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_6; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_7; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_8; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_9; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_10; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_11; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_12; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_13; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_14; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_15; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_16; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_17; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_18; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_19; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_20; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_21; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_22; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_23; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_24; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_25; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_26; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_27; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_28; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_29; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_30; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_31; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_32; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_33; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_34; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_35; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_36; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_37; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_38; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_39; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_40; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_41; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_42; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_43; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_44; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_45; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_46; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_47; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_48; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_49; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_50; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_51; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_52; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_53; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_54; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_55; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_56; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_57; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_58; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_59; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_60; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_61; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_62; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_63; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_64; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_65; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_66; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_67; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_68; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_69; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_70; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_71; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_72; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_73; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_74; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_75; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_76; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_77; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_78; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_79; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_80; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_81; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_82; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_83; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_84; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_85; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_86; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_87; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_88; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_89; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_90; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_91; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_92; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_93; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_94; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_95; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_96; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_97; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_98; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_99; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_100; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_101; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_102; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_103; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_104; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_105; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_106; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_107; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_108; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_109; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_110; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_111; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_112; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_113; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_114; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_115; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_116; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_117; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_118; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_119; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_120; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_121; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_122; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_123; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_124; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_125; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_126; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_127; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_128; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_129; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_130; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_131; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_132; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_133; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_134; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_135; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_136; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_137; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_138; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_139; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_140; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_141; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_142; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_143; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_144; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_145; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_146; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_147; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_148; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_149; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_150; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_151; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_152; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_153; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_154; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_155; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_156; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_157; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_158; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_159; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_160; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_161; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_162; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_163; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_164; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_165; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_166; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_167; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_168; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_169; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_170; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_171; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_172; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_173; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_174; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_175; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_176; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_177; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_178; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_179; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_180; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_181; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_182; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_183; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_184; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_185; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_186; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_187; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_188; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_189; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_190; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_191; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_192; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_193; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_194; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_195; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_196; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_197; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_198; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_199; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_200; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_201; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_202; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_203; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_204; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_205; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_206; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_207; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_208; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_209; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_210; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_211; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_212; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_213; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_214; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_215; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_216; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_217; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_218; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_219; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_220; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_221; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_222; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_223; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_224; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_225; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_226; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_227; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_228; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_229; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_230; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_231; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_232; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_233; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_234; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_235; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_236; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_237; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_238; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_239; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_240; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_241; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_242; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_243; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_244; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_245; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_246; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_247; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_248; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_249; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_250; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_251; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_252; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_253; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_254; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_255; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_256; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_257; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_258; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_259; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_260; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_261; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_262; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_263; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_264; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_265; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_266; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_267; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_268; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_269; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_270; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_271; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_272; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_273; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_274; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_275; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_276; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_277; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_278; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_279; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_280; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_281; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_282; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_283; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_284; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_285; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_286; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_287; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_288; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_289; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_290; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_291; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_292; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_293; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_294; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_295; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_296; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_297; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_298; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_299; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_300; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_301; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_302; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_303; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_304; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_305; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_306; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_307; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_308; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_309; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_310; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_311; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_312; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_313; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_314; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_315; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_316; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_317; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_318; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_319; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_320; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_321; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_322; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_323; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_324; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_325; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_326; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_327; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_328; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_329; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_330; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_331; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_332; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_333; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_334; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_335; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_336; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_337; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_338; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_339; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_340; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_341; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_342; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_343; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_344; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_345; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_346; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_347; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_348; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_349; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_350; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_351; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_352; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_353; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_354; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_355; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_356; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_357; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_358; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_359; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_360; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_361; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_362; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_363; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_364; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_365; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_366; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_367; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_368; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_369; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_370; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_371; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_372; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_373; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_374; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_375; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_376; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_377; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_378; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_379; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_380; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_381; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_382; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_383; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_384; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_385; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_386; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_387; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_388; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_389; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_390; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_391; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_392; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_393; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_394; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_395; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_396; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_397; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_398; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_399; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_400; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_401; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_402; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_403; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_404; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_405; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_406; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_407; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_408; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_409; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_410; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_411; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_412; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_413; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_414; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_415; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_416; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_417; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_418; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_419; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_420; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_421; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_422; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_423; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_424; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_425; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_426; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_427; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_428; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_429; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_430; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_431; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_432; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_433; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_434; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_435; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_436; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_437; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_438; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_439; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_440; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_441; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_442; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_443; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_444; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_445; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_446; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_447; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_448; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_449; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_450; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_451; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_452; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_453; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_454; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_455; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_456; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_457; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_458; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_459; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_460; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_461; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_462; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_463; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_464; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_465; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_466; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_467; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_468; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_469; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_470; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_471; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_472; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_473; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_474; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_475; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_476; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_477; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_478; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_479; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_480; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_481; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_482; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_483; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_484; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_485; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_486; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_487; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_488; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_489; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_490; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_491; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_492; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_493; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_494; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_495; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_496; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_497; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_498; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_499; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_500; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_501; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_502; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_503; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_504; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_505; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_506; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_507; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_508; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_509; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_510; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_511; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_0; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_1; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_2; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_3; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_4; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_5; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_6; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_7; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_8; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_9; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_10; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_11; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_12; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_13; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_14; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_15; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_state; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 343:23]
  wire [3:0] pipe1_io_pipe_phv_in_next_processor_id; // @[matcher.scala 343:23]
  wire  pipe1_io_pipe_phv_in_next_config_id; // @[matcher.scala 343:23]
  wire  pipe1_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_0; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_1; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_2; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_3; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_4; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_5; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_6; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_7; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_8; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_9; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_10; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_11; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_12; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_13; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_14; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_15; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_16; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_17; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_18; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_19; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_20; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_21; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_22; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_23; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_24; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_25; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_26; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_27; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_28; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_29; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_30; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_31; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_32; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_33; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_34; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_35; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_36; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_37; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_38; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_39; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_40; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_41; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_42; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_43; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_44; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_45; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_46; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_47; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_48; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_49; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_50; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_51; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_52; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_53; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_54; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_55; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_56; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_57; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_58; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_59; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_60; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_61; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_62; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_63; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_64; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_65; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_66; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_67; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_68; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_69; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_70; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_71; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_72; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_73; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_74; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_75; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_76; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_77; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_78; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_79; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_80; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_81; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_82; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_83; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_84; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_85; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_86; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_87; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_88; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_89; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_90; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_91; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_92; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_93; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_94; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_95; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_96; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_97; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_98; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_99; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_100; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_101; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_102; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_103; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_104; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_105; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_106; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_107; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_108; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_109; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_110; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_111; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_112; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_113; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_114; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_115; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_116; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_117; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_118; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_119; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_120; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_121; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_122; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_123; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_124; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_125; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_126; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_127; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_128; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_129; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_130; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_131; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_132; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_133; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_134; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_135; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_136; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_137; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_138; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_139; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_140; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_141; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_142; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_143; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_144; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_145; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_146; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_147; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_148; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_149; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_150; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_151; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_152; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_153; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_154; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_155; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_156; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_157; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_158; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_159; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_160; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_161; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_162; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_163; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_164; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_165; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_166; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_167; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_168; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_169; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_170; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_171; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_172; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_173; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_174; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_175; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_176; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_177; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_178; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_179; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_180; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_181; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_182; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_183; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_184; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_185; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_186; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_187; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_188; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_189; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_190; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_191; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_192; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_193; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_194; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_195; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_196; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_197; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_198; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_199; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_200; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_201; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_202; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_203; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_204; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_205; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_206; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_207; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_208; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_209; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_210; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_211; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_212; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_213; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_214; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_215; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_216; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_217; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_218; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_219; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_220; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_221; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_222; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_223; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_224; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_225; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_226; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_227; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_228; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_229; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_230; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_231; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_232; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_233; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_234; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_235; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_236; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_237; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_238; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_239; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_240; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_241; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_242; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_243; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_244; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_245; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_246; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_247; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_248; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_249; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_250; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_251; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_252; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_253; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_254; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_255; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_256; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_257; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_258; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_259; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_260; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_261; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_262; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_263; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_264; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_265; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_266; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_267; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_268; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_269; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_270; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_271; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_272; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_273; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_274; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_275; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_276; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_277; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_278; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_279; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_280; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_281; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_282; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_283; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_284; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_285; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_286; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_287; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_288; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_289; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_290; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_291; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_292; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_293; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_294; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_295; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_296; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_297; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_298; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_299; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_300; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_301; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_302; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_303; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_304; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_305; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_306; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_307; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_308; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_309; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_310; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_311; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_312; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_313; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_314; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_315; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_316; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_317; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_318; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_319; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_320; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_321; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_322; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_323; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_324; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_325; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_326; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_327; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_328; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_329; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_330; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_331; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_332; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_333; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_334; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_335; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_336; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_337; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_338; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_339; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_340; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_341; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_342; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_343; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_344; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_345; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_346; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_347; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_348; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_349; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_350; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_351; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_352; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_353; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_354; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_355; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_356; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_357; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_358; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_359; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_360; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_361; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_362; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_363; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_364; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_365; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_366; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_367; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_368; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_369; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_370; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_371; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_372; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_373; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_374; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_375; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_376; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_377; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_378; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_379; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_380; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_381; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_382; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_383; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_384; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_385; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_386; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_387; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_388; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_389; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_390; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_391; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_392; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_393; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_394; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_395; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_396; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_397; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_398; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_399; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_400; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_401; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_402; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_403; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_404; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_405; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_406; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_407; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_408; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_409; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_410; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_411; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_412; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_413; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_414; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_415; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_416; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_417; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_418; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_419; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_420; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_421; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_422; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_423; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_424; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_425; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_426; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_427; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_428; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_429; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_430; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_431; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_432; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_433; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_434; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_435; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_436; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_437; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_438; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_439; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_440; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_441; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_442; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_443; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_444; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_445; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_446; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_447; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_448; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_449; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_450; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_451; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_452; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_453; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_454; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_455; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_456; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_457; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_458; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_459; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_460; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_461; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_462; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_463; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_464; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_465; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_466; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_467; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_468; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_469; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_470; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_471; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_472; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_473; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_474; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_475; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_476; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_477; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_478; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_479; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_480; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_481; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_482; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_483; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_484; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_485; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_486; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_487; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_488; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_489; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_490; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_491; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_492; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_493; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_494; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_495; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_496; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_497; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_498; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_499; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_500; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_501; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_502; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_503; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_504; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_505; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_506; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_507; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_508; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_509; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_510; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_511; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_0; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_1; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_2; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_3; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_4; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_5; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_6; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_7; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_8; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_9; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_10; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_11; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_12; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_13; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_14; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_15; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_state; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 343:23]
  wire [3:0] pipe1_io_pipe_phv_out_next_processor_id; // @[matcher.scala 343:23]
  wire  pipe1_io_pipe_phv_out_next_config_id; // @[matcher.scala 343:23]
  wire  pipe1_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_key_config_0_header_id; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_key_config_0_internal_offset; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_key_config_1_header_id; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_key_config_1_internal_offset; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_key_offset; // @[matcher.scala 343:23]
  wire  pipe2_clock; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_0; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_1; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_2; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_3; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_4; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_5; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_6; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_7; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_8; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_9; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_10; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_11; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_12; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_13; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_14; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_15; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_16; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_17; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_18; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_19; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_20; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_21; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_22; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_23; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_24; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_25; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_26; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_27; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_28; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_29; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_30; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_31; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_32; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_33; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_34; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_35; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_36; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_37; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_38; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_39; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_40; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_41; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_42; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_43; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_44; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_45; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_46; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_47; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_48; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_49; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_50; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_51; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_52; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_53; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_54; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_55; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_56; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_57; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_58; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_59; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_60; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_61; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_62; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_63; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_64; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_65; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_66; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_67; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_68; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_69; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_70; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_71; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_72; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_73; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_74; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_75; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_76; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_77; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_78; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_79; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_80; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_81; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_82; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_83; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_84; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_85; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_86; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_87; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_88; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_89; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_90; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_91; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_92; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_93; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_94; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_95; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_96; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_97; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_98; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_99; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_100; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_101; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_102; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_103; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_104; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_105; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_106; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_107; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_108; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_109; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_110; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_111; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_112; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_113; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_114; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_115; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_116; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_117; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_118; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_119; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_120; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_121; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_122; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_123; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_124; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_125; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_126; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_127; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_128; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_129; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_130; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_131; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_132; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_133; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_134; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_135; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_136; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_137; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_138; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_139; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_140; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_141; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_142; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_143; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_144; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_145; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_146; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_147; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_148; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_149; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_150; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_151; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_152; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_153; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_154; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_155; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_156; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_157; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_158; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_159; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_160; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_161; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_162; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_163; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_164; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_165; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_166; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_167; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_168; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_169; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_170; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_171; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_172; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_173; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_174; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_175; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_176; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_177; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_178; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_179; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_180; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_181; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_182; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_183; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_184; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_185; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_186; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_187; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_188; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_189; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_190; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_191; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_192; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_193; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_194; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_195; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_196; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_197; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_198; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_199; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_200; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_201; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_202; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_203; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_204; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_205; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_206; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_207; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_208; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_209; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_210; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_211; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_212; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_213; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_214; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_215; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_216; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_217; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_218; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_219; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_220; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_221; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_222; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_223; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_224; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_225; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_226; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_227; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_228; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_229; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_230; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_231; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_232; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_233; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_234; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_235; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_236; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_237; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_238; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_239; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_240; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_241; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_242; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_243; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_244; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_245; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_246; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_247; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_248; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_249; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_250; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_251; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_252; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_253; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_254; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_255; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_256; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_257; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_258; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_259; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_260; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_261; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_262; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_263; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_264; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_265; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_266; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_267; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_268; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_269; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_270; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_271; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_272; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_273; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_274; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_275; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_276; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_277; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_278; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_279; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_280; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_281; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_282; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_283; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_284; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_285; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_286; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_287; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_288; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_289; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_290; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_291; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_292; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_293; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_294; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_295; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_296; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_297; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_298; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_299; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_300; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_301; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_302; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_303; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_304; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_305; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_306; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_307; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_308; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_309; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_310; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_311; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_312; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_313; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_314; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_315; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_316; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_317; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_318; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_319; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_320; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_321; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_322; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_323; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_324; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_325; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_326; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_327; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_328; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_329; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_330; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_331; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_332; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_333; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_334; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_335; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_336; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_337; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_338; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_339; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_340; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_341; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_342; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_343; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_344; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_345; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_346; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_347; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_348; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_349; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_350; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_351; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_352; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_353; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_354; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_355; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_356; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_357; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_358; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_359; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_360; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_361; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_362; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_363; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_364; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_365; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_366; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_367; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_368; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_369; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_370; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_371; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_372; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_373; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_374; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_375; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_376; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_377; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_378; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_379; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_380; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_381; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_382; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_383; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_384; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_385; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_386; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_387; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_388; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_389; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_390; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_391; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_392; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_393; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_394; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_395; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_396; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_397; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_398; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_399; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_400; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_401; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_402; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_403; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_404; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_405; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_406; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_407; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_408; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_409; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_410; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_411; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_412; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_413; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_414; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_415; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_416; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_417; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_418; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_419; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_420; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_421; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_422; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_423; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_424; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_425; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_426; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_427; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_428; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_429; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_430; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_431; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_432; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_433; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_434; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_435; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_436; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_437; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_438; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_439; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_440; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_441; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_442; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_443; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_444; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_445; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_446; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_447; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_448; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_449; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_450; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_451; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_452; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_453; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_454; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_455; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_456; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_457; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_458; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_459; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_460; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_461; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_462; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_463; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_464; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_465; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_466; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_467; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_468; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_469; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_470; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_471; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_472; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_473; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_474; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_475; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_476; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_477; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_478; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_479; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_480; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_481; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_482; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_483; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_484; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_485; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_486; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_487; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_488; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_489; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_490; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_491; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_492; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_493; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_494; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_495; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_496; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_497; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_498; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_499; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_500; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_501; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_502; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_503; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_504; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_505; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_506; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_507; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_508; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_509; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_510; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_511; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_0; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_1; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_2; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_3; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_4; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_5; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_6; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_7; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_8; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_9; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_10; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_11; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_12; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_13; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_14; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_15; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_state; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 344:23]
  wire [3:0] pipe2_io_pipe_phv_in_next_processor_id; // @[matcher.scala 344:23]
  wire  pipe2_io_pipe_phv_in_next_config_id; // @[matcher.scala 344:23]
  wire  pipe2_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_0; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_1; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_2; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_3; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_4; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_5; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_6; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_7; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_8; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_9; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_10; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_11; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_12; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_13; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_14; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_15; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_16; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_17; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_18; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_19; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_20; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_21; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_22; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_23; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_24; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_25; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_26; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_27; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_28; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_29; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_30; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_31; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_32; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_33; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_34; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_35; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_36; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_37; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_38; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_39; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_40; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_41; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_42; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_43; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_44; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_45; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_46; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_47; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_48; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_49; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_50; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_51; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_52; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_53; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_54; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_55; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_56; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_57; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_58; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_59; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_60; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_61; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_62; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_63; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_64; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_65; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_66; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_67; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_68; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_69; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_70; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_71; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_72; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_73; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_74; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_75; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_76; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_77; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_78; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_79; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_80; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_81; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_82; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_83; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_84; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_85; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_86; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_87; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_88; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_89; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_90; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_91; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_92; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_93; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_94; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_95; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_96; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_97; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_98; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_99; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_100; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_101; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_102; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_103; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_104; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_105; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_106; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_107; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_108; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_109; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_110; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_111; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_112; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_113; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_114; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_115; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_116; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_117; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_118; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_119; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_120; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_121; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_122; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_123; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_124; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_125; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_126; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_127; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_128; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_129; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_130; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_131; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_132; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_133; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_134; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_135; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_136; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_137; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_138; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_139; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_140; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_141; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_142; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_143; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_144; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_145; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_146; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_147; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_148; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_149; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_150; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_151; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_152; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_153; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_154; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_155; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_156; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_157; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_158; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_159; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_160; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_161; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_162; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_163; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_164; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_165; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_166; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_167; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_168; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_169; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_170; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_171; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_172; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_173; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_174; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_175; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_176; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_177; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_178; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_179; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_180; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_181; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_182; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_183; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_184; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_185; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_186; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_187; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_188; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_189; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_190; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_191; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_192; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_193; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_194; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_195; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_196; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_197; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_198; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_199; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_200; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_201; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_202; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_203; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_204; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_205; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_206; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_207; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_208; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_209; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_210; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_211; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_212; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_213; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_214; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_215; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_216; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_217; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_218; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_219; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_220; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_221; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_222; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_223; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_224; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_225; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_226; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_227; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_228; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_229; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_230; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_231; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_232; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_233; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_234; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_235; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_236; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_237; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_238; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_239; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_240; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_241; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_242; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_243; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_244; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_245; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_246; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_247; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_248; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_249; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_250; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_251; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_252; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_253; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_254; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_255; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_256; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_257; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_258; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_259; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_260; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_261; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_262; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_263; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_264; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_265; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_266; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_267; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_268; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_269; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_270; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_271; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_272; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_273; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_274; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_275; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_276; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_277; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_278; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_279; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_280; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_281; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_282; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_283; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_284; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_285; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_286; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_287; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_288; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_289; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_290; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_291; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_292; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_293; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_294; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_295; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_296; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_297; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_298; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_299; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_300; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_301; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_302; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_303; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_304; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_305; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_306; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_307; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_308; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_309; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_310; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_311; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_312; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_313; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_314; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_315; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_316; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_317; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_318; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_319; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_320; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_321; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_322; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_323; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_324; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_325; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_326; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_327; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_328; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_329; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_330; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_331; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_332; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_333; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_334; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_335; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_336; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_337; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_338; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_339; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_340; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_341; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_342; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_343; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_344; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_345; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_346; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_347; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_348; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_349; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_350; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_351; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_352; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_353; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_354; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_355; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_356; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_357; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_358; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_359; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_360; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_361; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_362; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_363; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_364; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_365; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_366; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_367; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_368; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_369; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_370; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_371; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_372; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_373; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_374; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_375; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_376; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_377; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_378; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_379; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_380; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_381; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_382; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_383; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_384; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_385; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_386; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_387; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_388; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_389; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_390; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_391; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_392; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_393; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_394; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_395; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_396; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_397; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_398; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_399; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_400; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_401; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_402; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_403; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_404; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_405; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_406; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_407; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_408; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_409; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_410; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_411; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_412; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_413; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_414; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_415; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_416; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_417; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_418; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_419; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_420; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_421; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_422; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_423; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_424; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_425; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_426; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_427; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_428; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_429; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_430; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_431; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_432; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_433; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_434; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_435; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_436; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_437; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_438; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_439; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_440; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_441; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_442; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_443; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_444; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_445; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_446; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_447; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_448; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_449; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_450; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_451; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_452; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_453; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_454; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_455; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_456; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_457; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_458; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_459; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_460; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_461; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_462; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_463; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_464; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_465; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_466; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_467; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_468; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_469; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_470; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_471; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_472; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_473; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_474; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_475; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_476; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_477; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_478; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_479; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_480; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_481; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_482; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_483; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_484; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_485; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_486; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_487; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_488; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_489; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_490; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_491; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_492; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_493; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_494; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_495; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_496; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_497; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_498; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_499; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_500; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_501; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_502; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_503; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_504; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_505; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_506; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_507; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_508; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_509; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_510; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_511; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_0; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_1; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_2; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_3; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_4; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_5; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_6; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_7; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_8; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_9; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_10; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_11; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_12; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_13; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_14; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_15; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_state; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 344:23]
  wire [3:0] pipe2_io_pipe_phv_out_next_processor_id; // @[matcher.scala 344:23]
  wire  pipe2_io_pipe_phv_out_next_config_id; // @[matcher.scala 344:23]
  wire  pipe2_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_key_config_0_key_length; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_key_config_1_key_length; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_key_offset; // @[matcher.scala 344:23]
  wire [191:0] pipe2_io_match_key; // @[matcher.scala 344:23]
  wire  pipe3to8_clock; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_0; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_1; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_2; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_3; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_4; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_5; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_6; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_7; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_8; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_9; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_10; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_11; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_12; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_13; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_14; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_15; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_16; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_17; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_18; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_19; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_20; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_21; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_22; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_23; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_24; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_25; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_26; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_27; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_28; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_29; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_30; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_31; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_32; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_33; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_34; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_35; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_36; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_37; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_38; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_39; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_40; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_41; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_42; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_43; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_44; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_45; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_46; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_47; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_48; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_49; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_50; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_51; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_52; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_53; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_54; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_55; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_56; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_57; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_58; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_59; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_60; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_61; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_62; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_63; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_64; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_65; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_66; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_67; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_68; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_69; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_70; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_71; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_72; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_73; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_74; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_75; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_76; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_77; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_78; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_79; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_80; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_81; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_82; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_83; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_84; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_85; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_86; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_87; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_88; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_89; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_90; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_91; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_92; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_93; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_94; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_95; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_96; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_97; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_98; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_99; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_100; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_101; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_102; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_103; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_104; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_105; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_106; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_107; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_108; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_109; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_110; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_111; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_112; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_113; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_114; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_115; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_116; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_117; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_118; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_119; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_120; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_121; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_122; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_123; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_124; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_125; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_126; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_127; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_128; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_129; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_130; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_131; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_132; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_133; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_134; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_135; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_136; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_137; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_138; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_139; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_140; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_141; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_142; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_143; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_144; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_145; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_146; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_147; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_148; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_149; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_150; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_151; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_152; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_153; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_154; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_155; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_156; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_157; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_158; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_159; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_160; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_161; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_162; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_163; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_164; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_165; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_166; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_167; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_168; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_169; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_170; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_171; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_172; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_173; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_174; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_175; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_176; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_177; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_178; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_179; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_180; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_181; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_182; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_183; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_184; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_185; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_186; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_187; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_188; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_189; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_190; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_191; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_192; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_193; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_194; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_195; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_196; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_197; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_198; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_199; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_200; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_201; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_202; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_203; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_204; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_205; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_206; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_207; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_208; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_209; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_210; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_211; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_212; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_213; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_214; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_215; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_216; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_217; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_218; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_219; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_220; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_221; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_222; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_223; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_224; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_225; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_226; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_227; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_228; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_229; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_230; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_231; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_232; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_233; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_234; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_235; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_236; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_237; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_238; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_239; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_240; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_241; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_242; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_243; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_244; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_245; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_246; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_247; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_248; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_249; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_250; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_251; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_252; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_253; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_254; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_255; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_256; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_257; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_258; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_259; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_260; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_261; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_262; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_263; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_264; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_265; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_266; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_267; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_268; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_269; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_270; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_271; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_272; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_273; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_274; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_275; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_276; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_277; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_278; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_279; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_280; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_281; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_282; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_283; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_284; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_285; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_286; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_287; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_288; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_289; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_290; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_291; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_292; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_293; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_294; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_295; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_296; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_297; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_298; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_299; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_300; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_301; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_302; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_303; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_304; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_305; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_306; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_307; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_308; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_309; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_310; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_311; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_312; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_313; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_314; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_315; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_316; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_317; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_318; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_319; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_320; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_321; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_322; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_323; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_324; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_325; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_326; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_327; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_328; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_329; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_330; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_331; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_332; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_333; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_334; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_335; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_336; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_337; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_338; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_339; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_340; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_341; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_342; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_343; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_344; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_345; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_346; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_347; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_348; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_349; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_350; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_351; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_352; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_353; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_354; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_355; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_356; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_357; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_358; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_359; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_360; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_361; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_362; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_363; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_364; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_365; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_366; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_367; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_368; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_369; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_370; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_371; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_372; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_373; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_374; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_375; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_376; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_377; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_378; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_379; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_380; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_381; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_382; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_383; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_384; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_385; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_386; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_387; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_388; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_389; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_390; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_391; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_392; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_393; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_394; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_395; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_396; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_397; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_398; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_399; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_400; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_401; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_402; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_403; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_404; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_405; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_406; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_407; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_408; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_409; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_410; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_411; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_412; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_413; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_414; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_415; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_416; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_417; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_418; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_419; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_420; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_421; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_422; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_423; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_424; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_425; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_426; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_427; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_428; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_429; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_430; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_431; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_432; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_433; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_434; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_435; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_436; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_437; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_438; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_439; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_440; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_441; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_442; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_443; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_444; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_445; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_446; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_447; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_448; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_449; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_450; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_451; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_452; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_453; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_454; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_455; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_456; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_457; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_458; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_459; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_460; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_461; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_462; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_463; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_464; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_465; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_466; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_467; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_468; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_469; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_470; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_471; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_472; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_473; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_474; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_475; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_476; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_477; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_478; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_479; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_480; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_481; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_482; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_483; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_484; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_485; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_486; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_487; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_488; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_489; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_490; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_491; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_492; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_493; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_494; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_495; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_496; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_497; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_498; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_499; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_500; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_501; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_502; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_503; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_504; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_505; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_506; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_507; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_508; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_509; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_510; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_511; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_0; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_1; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_2; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_3; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_4; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_5; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_6; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_7; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_8; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_9; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_10; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_11; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_12; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_13; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_14; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_15; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_parse_current_state; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 345:26]
  wire [3:0] pipe3to8_io_pipe_phv_in_next_processor_id; // @[matcher.scala 345:26]
  wire  pipe3to8_io_pipe_phv_in_next_config_id; // @[matcher.scala 345:26]
  wire  pipe3to8_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_0; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_1; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_2; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_3; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_4; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_5; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_6; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_7; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_8; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_9; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_10; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_11; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_12; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_13; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_14; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_15; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_16; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_17; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_18; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_19; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_20; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_21; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_22; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_23; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_24; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_25; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_26; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_27; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_28; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_29; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_30; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_31; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_32; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_33; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_34; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_35; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_36; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_37; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_38; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_39; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_40; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_41; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_42; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_43; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_44; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_45; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_46; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_47; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_48; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_49; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_50; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_51; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_52; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_53; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_54; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_55; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_56; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_57; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_58; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_59; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_60; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_61; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_62; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_63; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_64; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_65; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_66; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_67; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_68; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_69; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_70; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_71; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_72; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_73; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_74; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_75; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_76; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_77; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_78; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_79; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_80; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_81; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_82; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_83; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_84; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_85; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_86; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_87; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_88; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_89; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_90; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_91; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_92; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_93; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_94; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_95; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_96; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_97; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_98; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_99; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_100; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_101; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_102; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_103; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_104; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_105; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_106; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_107; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_108; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_109; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_110; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_111; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_112; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_113; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_114; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_115; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_116; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_117; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_118; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_119; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_120; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_121; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_122; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_123; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_124; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_125; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_126; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_127; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_128; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_129; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_130; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_131; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_132; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_133; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_134; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_135; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_136; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_137; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_138; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_139; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_140; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_141; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_142; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_143; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_144; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_145; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_146; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_147; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_148; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_149; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_150; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_151; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_152; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_153; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_154; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_155; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_156; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_157; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_158; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_159; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_160; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_161; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_162; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_163; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_164; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_165; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_166; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_167; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_168; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_169; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_170; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_171; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_172; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_173; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_174; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_175; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_176; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_177; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_178; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_179; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_180; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_181; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_182; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_183; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_184; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_185; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_186; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_187; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_188; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_189; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_190; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_191; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_192; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_193; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_194; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_195; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_196; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_197; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_198; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_199; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_200; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_201; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_202; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_203; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_204; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_205; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_206; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_207; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_208; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_209; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_210; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_211; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_212; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_213; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_214; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_215; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_216; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_217; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_218; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_219; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_220; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_221; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_222; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_223; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_224; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_225; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_226; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_227; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_228; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_229; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_230; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_231; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_232; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_233; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_234; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_235; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_236; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_237; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_238; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_239; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_240; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_241; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_242; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_243; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_244; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_245; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_246; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_247; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_248; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_249; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_250; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_251; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_252; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_253; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_254; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_255; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_256; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_257; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_258; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_259; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_260; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_261; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_262; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_263; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_264; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_265; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_266; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_267; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_268; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_269; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_270; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_271; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_272; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_273; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_274; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_275; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_276; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_277; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_278; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_279; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_280; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_281; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_282; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_283; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_284; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_285; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_286; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_287; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_288; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_289; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_290; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_291; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_292; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_293; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_294; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_295; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_296; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_297; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_298; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_299; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_300; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_301; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_302; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_303; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_304; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_305; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_306; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_307; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_308; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_309; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_310; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_311; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_312; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_313; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_314; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_315; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_316; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_317; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_318; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_319; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_320; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_321; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_322; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_323; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_324; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_325; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_326; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_327; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_328; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_329; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_330; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_331; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_332; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_333; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_334; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_335; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_336; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_337; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_338; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_339; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_340; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_341; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_342; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_343; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_344; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_345; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_346; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_347; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_348; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_349; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_350; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_351; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_352; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_353; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_354; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_355; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_356; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_357; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_358; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_359; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_360; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_361; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_362; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_363; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_364; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_365; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_366; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_367; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_368; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_369; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_370; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_371; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_372; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_373; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_374; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_375; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_376; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_377; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_378; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_379; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_380; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_381; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_382; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_383; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_384; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_385; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_386; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_387; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_388; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_389; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_390; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_391; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_392; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_393; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_394; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_395; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_396; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_397; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_398; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_399; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_400; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_401; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_402; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_403; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_404; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_405; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_406; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_407; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_408; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_409; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_410; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_411; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_412; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_413; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_414; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_415; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_416; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_417; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_418; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_419; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_420; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_421; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_422; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_423; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_424; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_425; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_426; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_427; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_428; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_429; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_430; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_431; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_432; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_433; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_434; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_435; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_436; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_437; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_438; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_439; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_440; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_441; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_442; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_443; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_444; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_445; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_446; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_447; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_448; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_449; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_450; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_451; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_452; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_453; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_454; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_455; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_456; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_457; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_458; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_459; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_460; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_461; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_462; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_463; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_464; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_465; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_466; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_467; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_468; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_469; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_470; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_471; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_472; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_473; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_474; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_475; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_476; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_477; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_478; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_479; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_480; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_481; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_482; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_483; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_484; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_485; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_486; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_487; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_488; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_489; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_490; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_491; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_492; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_493; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_494; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_495; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_496; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_497; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_498; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_499; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_500; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_501; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_502; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_503; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_504; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_505; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_506; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_507; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_508; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_509; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_510; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_511; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_0; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_1; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_2; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_3; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_4; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_5; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_6; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_7; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_8; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_9; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_10; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_11; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_12; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_13; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_14; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_15; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_parse_current_state; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 345:26]
  wire [3:0] pipe3to8_io_pipe_phv_out_next_processor_id; // @[matcher.scala 345:26]
  wire  pipe3to8_io_pipe_phv_out_next_config_id; // @[matcher.scala 345:26]
  wire  pipe3to8_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 345:26]
  wire  pipe3to8_io_mod_hash_depth_mod; // @[matcher.scala 345:26]
  wire  pipe3to8_io_mod_config_id; // @[matcher.scala 345:26]
  wire [3:0] pipe3to8_io_mod_hash_depth; // @[matcher.scala 345:26]
  wire [191:0] pipe3to8_io_key_in; // @[matcher.scala 345:26]
  wire [191:0] pipe3to8_io_key_out; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_hash_val; // @[matcher.scala 345:26]
  wire [3:0] pipe3to8_io_hash_val_cs; // @[matcher.scala 345:26]
  wire  pipe9_clock; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_0; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_1; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_2; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_3; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_4; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_5; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_6; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_7; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_8; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_9; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_10; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_11; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_12; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_13; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_14; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_15; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_16; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_17; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_18; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_19; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_20; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_21; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_22; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_23; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_24; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_25; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_26; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_27; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_28; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_29; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_30; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_31; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_32; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_33; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_34; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_35; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_36; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_37; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_38; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_39; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_40; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_41; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_42; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_43; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_44; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_45; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_46; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_47; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_48; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_49; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_50; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_51; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_52; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_53; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_54; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_55; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_56; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_57; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_58; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_59; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_60; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_61; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_62; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_63; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_64; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_65; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_66; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_67; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_68; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_69; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_70; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_71; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_72; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_73; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_74; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_75; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_76; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_77; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_78; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_79; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_80; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_81; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_82; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_83; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_84; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_85; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_86; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_87; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_88; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_89; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_90; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_91; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_92; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_93; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_94; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_95; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_96; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_97; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_98; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_99; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_100; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_101; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_102; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_103; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_104; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_105; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_106; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_107; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_108; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_109; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_110; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_111; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_112; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_113; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_114; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_115; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_116; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_117; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_118; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_119; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_120; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_121; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_122; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_123; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_124; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_125; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_126; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_127; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_128; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_129; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_130; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_131; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_132; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_133; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_134; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_135; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_136; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_137; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_138; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_139; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_140; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_141; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_142; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_143; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_144; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_145; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_146; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_147; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_148; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_149; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_150; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_151; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_152; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_153; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_154; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_155; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_156; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_157; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_158; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_159; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_160; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_161; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_162; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_163; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_164; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_165; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_166; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_167; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_168; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_169; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_170; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_171; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_172; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_173; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_174; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_175; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_176; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_177; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_178; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_179; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_180; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_181; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_182; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_183; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_184; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_185; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_186; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_187; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_188; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_189; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_190; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_191; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_192; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_193; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_194; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_195; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_196; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_197; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_198; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_199; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_200; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_201; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_202; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_203; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_204; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_205; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_206; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_207; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_208; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_209; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_210; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_211; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_212; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_213; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_214; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_215; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_216; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_217; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_218; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_219; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_220; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_221; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_222; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_223; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_224; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_225; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_226; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_227; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_228; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_229; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_230; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_231; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_232; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_233; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_234; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_235; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_236; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_237; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_238; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_239; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_240; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_241; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_242; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_243; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_244; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_245; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_246; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_247; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_248; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_249; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_250; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_251; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_252; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_253; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_254; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_255; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_256; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_257; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_258; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_259; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_260; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_261; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_262; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_263; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_264; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_265; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_266; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_267; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_268; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_269; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_270; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_271; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_272; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_273; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_274; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_275; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_276; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_277; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_278; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_279; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_280; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_281; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_282; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_283; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_284; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_285; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_286; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_287; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_288; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_289; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_290; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_291; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_292; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_293; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_294; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_295; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_296; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_297; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_298; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_299; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_300; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_301; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_302; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_303; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_304; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_305; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_306; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_307; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_308; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_309; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_310; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_311; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_312; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_313; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_314; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_315; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_316; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_317; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_318; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_319; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_320; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_321; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_322; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_323; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_324; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_325; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_326; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_327; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_328; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_329; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_330; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_331; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_332; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_333; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_334; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_335; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_336; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_337; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_338; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_339; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_340; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_341; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_342; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_343; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_344; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_345; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_346; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_347; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_348; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_349; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_350; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_351; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_352; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_353; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_354; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_355; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_356; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_357; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_358; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_359; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_360; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_361; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_362; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_363; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_364; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_365; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_366; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_367; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_368; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_369; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_370; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_371; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_372; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_373; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_374; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_375; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_376; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_377; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_378; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_379; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_380; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_381; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_382; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_383; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_384; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_385; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_386; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_387; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_388; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_389; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_390; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_391; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_392; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_393; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_394; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_395; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_396; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_397; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_398; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_399; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_400; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_401; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_402; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_403; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_404; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_405; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_406; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_407; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_408; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_409; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_410; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_411; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_412; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_413; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_414; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_415; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_416; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_417; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_418; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_419; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_420; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_421; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_422; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_423; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_424; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_425; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_426; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_427; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_428; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_429; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_430; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_431; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_432; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_433; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_434; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_435; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_436; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_437; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_438; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_439; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_440; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_441; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_442; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_443; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_444; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_445; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_446; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_447; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_448; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_449; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_450; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_451; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_452; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_453; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_454; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_455; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_456; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_457; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_458; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_459; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_460; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_461; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_462; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_463; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_464; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_465; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_466; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_467; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_468; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_469; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_470; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_471; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_472; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_473; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_474; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_475; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_476; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_477; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_478; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_479; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_480; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_481; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_482; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_483; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_484; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_485; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_486; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_487; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_488; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_489; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_490; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_491; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_492; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_493; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_494; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_495; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_496; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_497; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_498; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_499; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_500; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_501; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_502; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_503; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_504; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_505; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_506; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_507; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_508; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_509; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_510; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_511; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_0; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_1; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_2; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_3; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_4; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_5; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_6; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_7; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_8; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_9; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_10; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_11; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_12; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_13; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_14; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_15; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_parse_current_state; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 346:23]
  wire [3:0] pipe9_io_pipe_phv_in_next_processor_id; // @[matcher.scala 346:23]
  wire  pipe9_io_pipe_phv_in_next_config_id; // @[matcher.scala 346:23]
  wire  pipe9_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_0; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_1; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_2; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_3; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_4; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_5; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_6; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_7; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_8; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_9; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_10; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_11; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_12; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_13; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_14; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_15; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_16; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_17; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_18; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_19; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_20; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_21; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_22; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_23; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_24; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_25; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_26; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_27; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_28; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_29; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_30; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_31; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_32; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_33; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_34; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_35; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_36; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_37; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_38; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_39; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_40; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_41; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_42; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_43; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_44; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_45; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_46; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_47; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_48; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_49; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_50; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_51; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_52; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_53; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_54; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_55; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_56; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_57; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_58; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_59; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_60; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_61; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_62; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_63; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_64; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_65; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_66; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_67; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_68; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_69; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_70; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_71; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_72; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_73; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_74; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_75; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_76; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_77; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_78; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_79; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_80; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_81; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_82; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_83; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_84; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_85; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_86; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_87; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_88; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_89; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_90; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_91; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_92; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_93; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_94; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_95; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_96; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_97; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_98; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_99; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_100; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_101; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_102; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_103; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_104; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_105; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_106; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_107; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_108; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_109; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_110; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_111; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_112; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_113; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_114; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_115; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_116; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_117; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_118; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_119; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_120; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_121; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_122; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_123; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_124; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_125; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_126; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_127; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_128; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_129; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_130; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_131; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_132; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_133; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_134; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_135; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_136; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_137; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_138; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_139; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_140; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_141; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_142; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_143; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_144; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_145; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_146; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_147; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_148; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_149; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_150; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_151; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_152; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_153; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_154; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_155; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_156; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_157; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_158; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_159; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_160; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_161; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_162; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_163; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_164; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_165; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_166; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_167; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_168; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_169; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_170; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_171; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_172; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_173; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_174; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_175; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_176; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_177; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_178; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_179; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_180; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_181; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_182; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_183; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_184; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_185; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_186; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_187; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_188; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_189; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_190; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_191; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_192; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_193; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_194; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_195; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_196; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_197; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_198; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_199; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_200; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_201; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_202; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_203; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_204; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_205; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_206; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_207; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_208; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_209; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_210; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_211; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_212; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_213; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_214; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_215; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_216; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_217; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_218; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_219; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_220; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_221; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_222; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_223; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_224; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_225; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_226; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_227; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_228; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_229; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_230; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_231; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_232; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_233; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_234; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_235; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_236; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_237; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_238; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_239; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_240; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_241; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_242; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_243; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_244; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_245; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_246; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_247; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_248; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_249; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_250; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_251; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_252; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_253; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_254; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_255; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_256; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_257; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_258; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_259; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_260; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_261; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_262; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_263; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_264; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_265; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_266; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_267; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_268; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_269; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_270; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_271; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_272; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_273; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_274; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_275; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_276; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_277; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_278; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_279; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_280; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_281; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_282; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_283; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_284; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_285; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_286; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_287; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_288; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_289; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_290; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_291; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_292; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_293; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_294; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_295; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_296; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_297; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_298; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_299; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_300; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_301; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_302; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_303; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_304; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_305; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_306; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_307; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_308; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_309; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_310; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_311; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_312; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_313; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_314; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_315; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_316; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_317; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_318; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_319; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_320; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_321; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_322; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_323; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_324; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_325; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_326; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_327; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_328; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_329; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_330; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_331; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_332; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_333; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_334; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_335; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_336; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_337; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_338; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_339; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_340; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_341; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_342; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_343; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_344; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_345; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_346; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_347; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_348; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_349; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_350; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_351; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_352; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_353; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_354; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_355; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_356; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_357; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_358; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_359; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_360; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_361; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_362; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_363; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_364; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_365; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_366; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_367; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_368; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_369; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_370; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_371; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_372; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_373; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_374; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_375; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_376; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_377; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_378; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_379; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_380; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_381; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_382; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_383; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_384; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_385; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_386; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_387; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_388; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_389; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_390; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_391; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_392; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_393; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_394; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_395; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_396; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_397; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_398; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_399; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_400; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_401; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_402; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_403; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_404; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_405; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_406; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_407; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_408; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_409; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_410; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_411; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_412; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_413; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_414; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_415; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_416; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_417; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_418; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_419; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_420; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_421; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_422; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_423; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_424; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_425; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_426; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_427; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_428; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_429; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_430; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_431; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_432; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_433; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_434; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_435; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_436; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_437; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_438; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_439; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_440; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_441; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_442; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_443; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_444; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_445; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_446; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_447; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_448; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_449; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_450; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_451; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_452; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_453; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_454; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_455; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_456; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_457; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_458; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_459; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_460; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_461; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_462; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_463; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_464; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_465; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_466; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_467; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_468; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_469; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_470; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_471; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_472; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_473; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_474; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_475; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_476; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_477; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_478; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_479; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_480; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_481; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_482; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_483; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_484; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_485; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_486; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_487; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_488; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_489; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_490; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_491; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_492; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_493; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_494; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_495; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_496; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_497; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_498; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_499; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_500; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_501; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_502; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_503; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_504; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_505; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_506; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_507; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_508; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_509; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_510; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_511; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_0; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_1; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_2; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_3; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_4; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_5; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_6; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_7; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_8; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_9; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_10; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_11; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_12; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_13; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_14; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_15; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_parse_current_state; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 346:23]
  wire [3:0] pipe9_io_pipe_phv_out_next_processor_id; // @[matcher.scala 346:23]
  wire  pipe9_io_pipe_phv_out_next_config_id; // @[matcher.scala 346:23]
  wire  pipe9_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 346:23]
  wire [4:0] pipe9_io_table_config_0_table_width; // @[matcher.scala 346:23]
  wire [4:0] pipe9_io_table_config_0_table_depth; // @[matcher.scala 346:23]
  wire [4:0] pipe9_io_table_config_1_table_width; // @[matcher.scala 346:23]
  wire [4:0] pipe9_io_table_config_1_table_depth; // @[matcher.scala 346:23]
  wire [191:0] pipe9_io_key_in; // @[matcher.scala 346:23]
  wire [191:0] pipe9_io_key_out; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_addr_in; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_addr_out; // @[matcher.scala 346:23]
  wire [3:0] pipe9_io_cs_in; // @[matcher.scala 346:23]
  wire [3:0] pipe9_io_cs_out; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_0; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_1; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_2; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_3; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_4; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_5; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_6; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_7; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_8; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_9; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_10; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_11; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_12; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_13; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_14; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_15; // @[matcher.scala 346:23]
  wire  pipe10_clock; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_0; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_1; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_2; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_3; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_4; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_5; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_6; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_7; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_8; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_9; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_10; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_11; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_12; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_13; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_14; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_15; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_16; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_17; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_18; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_19; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_20; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_21; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_22; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_23; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_24; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_25; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_26; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_27; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_28; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_29; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_30; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_31; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_32; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_33; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_34; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_35; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_36; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_37; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_38; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_39; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_40; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_41; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_42; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_43; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_44; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_45; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_46; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_47; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_48; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_49; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_50; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_51; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_52; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_53; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_54; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_55; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_56; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_57; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_58; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_59; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_60; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_61; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_62; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_63; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_64; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_65; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_66; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_67; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_68; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_69; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_70; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_71; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_72; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_73; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_74; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_75; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_76; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_77; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_78; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_79; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_80; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_81; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_82; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_83; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_84; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_85; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_86; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_87; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_88; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_89; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_90; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_91; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_92; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_93; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_94; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_95; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_96; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_97; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_98; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_99; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_100; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_101; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_102; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_103; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_104; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_105; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_106; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_107; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_108; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_109; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_110; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_111; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_112; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_113; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_114; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_115; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_116; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_117; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_118; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_119; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_120; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_121; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_122; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_123; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_124; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_125; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_126; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_127; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_128; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_129; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_130; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_131; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_132; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_133; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_134; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_135; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_136; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_137; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_138; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_139; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_140; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_141; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_142; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_143; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_144; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_145; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_146; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_147; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_148; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_149; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_150; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_151; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_152; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_153; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_154; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_155; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_156; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_157; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_158; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_159; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_160; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_161; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_162; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_163; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_164; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_165; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_166; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_167; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_168; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_169; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_170; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_171; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_172; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_173; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_174; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_175; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_176; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_177; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_178; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_179; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_180; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_181; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_182; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_183; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_184; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_185; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_186; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_187; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_188; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_189; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_190; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_191; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_192; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_193; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_194; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_195; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_196; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_197; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_198; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_199; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_200; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_201; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_202; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_203; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_204; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_205; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_206; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_207; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_208; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_209; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_210; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_211; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_212; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_213; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_214; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_215; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_216; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_217; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_218; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_219; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_220; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_221; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_222; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_223; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_224; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_225; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_226; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_227; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_228; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_229; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_230; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_231; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_232; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_233; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_234; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_235; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_236; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_237; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_238; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_239; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_240; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_241; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_242; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_243; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_244; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_245; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_246; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_247; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_248; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_249; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_250; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_251; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_252; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_253; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_254; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_255; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_256; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_257; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_258; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_259; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_260; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_261; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_262; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_263; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_264; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_265; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_266; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_267; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_268; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_269; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_270; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_271; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_272; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_273; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_274; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_275; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_276; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_277; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_278; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_279; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_280; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_281; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_282; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_283; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_284; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_285; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_286; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_287; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_288; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_289; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_290; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_291; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_292; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_293; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_294; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_295; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_296; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_297; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_298; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_299; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_300; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_301; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_302; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_303; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_304; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_305; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_306; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_307; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_308; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_309; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_310; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_311; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_312; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_313; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_314; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_315; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_316; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_317; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_318; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_319; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_320; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_321; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_322; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_323; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_324; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_325; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_326; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_327; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_328; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_329; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_330; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_331; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_332; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_333; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_334; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_335; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_336; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_337; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_338; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_339; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_340; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_341; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_342; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_343; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_344; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_345; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_346; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_347; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_348; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_349; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_350; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_351; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_352; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_353; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_354; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_355; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_356; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_357; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_358; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_359; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_360; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_361; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_362; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_363; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_364; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_365; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_366; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_367; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_368; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_369; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_370; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_371; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_372; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_373; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_374; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_375; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_376; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_377; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_378; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_379; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_380; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_381; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_382; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_383; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_384; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_385; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_386; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_387; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_388; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_389; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_390; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_391; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_392; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_393; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_394; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_395; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_396; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_397; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_398; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_399; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_400; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_401; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_402; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_403; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_404; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_405; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_406; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_407; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_408; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_409; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_410; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_411; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_412; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_413; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_414; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_415; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_416; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_417; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_418; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_419; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_420; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_421; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_422; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_423; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_424; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_425; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_426; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_427; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_428; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_429; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_430; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_431; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_432; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_433; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_434; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_435; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_436; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_437; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_438; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_439; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_440; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_441; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_442; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_443; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_444; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_445; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_446; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_447; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_448; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_449; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_450; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_451; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_452; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_453; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_454; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_455; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_456; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_457; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_458; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_459; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_460; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_461; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_462; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_463; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_464; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_465; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_466; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_467; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_468; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_469; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_470; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_471; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_472; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_473; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_474; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_475; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_476; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_477; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_478; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_479; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_480; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_481; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_482; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_483; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_484; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_485; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_486; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_487; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_488; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_489; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_490; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_491; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_492; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_493; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_494; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_495; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_496; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_497; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_498; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_499; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_500; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_501; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_502; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_503; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_504; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_505; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_506; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_507; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_508; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_509; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_510; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_511; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_0; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_1; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_2; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_3; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_4; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_5; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_6; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_7; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_8; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_9; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_10; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_11; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_12; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_13; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_14; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_15; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_parse_current_state; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 347:24]
  wire [3:0] pipe10_io_pipe_phv_in_next_processor_id; // @[matcher.scala 347:24]
  wire  pipe10_io_pipe_phv_in_next_config_id; // @[matcher.scala 347:24]
  wire  pipe10_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_0; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_1; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_2; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_3; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_4; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_5; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_6; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_7; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_8; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_9; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_10; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_11; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_12; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_13; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_14; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_15; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_16; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_17; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_18; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_19; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_20; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_21; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_22; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_23; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_24; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_25; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_26; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_27; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_28; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_29; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_30; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_31; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_32; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_33; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_34; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_35; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_36; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_37; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_38; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_39; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_40; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_41; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_42; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_43; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_44; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_45; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_46; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_47; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_48; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_49; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_50; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_51; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_52; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_53; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_54; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_55; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_56; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_57; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_58; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_59; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_60; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_61; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_62; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_63; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_64; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_65; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_66; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_67; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_68; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_69; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_70; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_71; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_72; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_73; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_74; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_75; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_76; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_77; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_78; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_79; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_80; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_81; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_82; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_83; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_84; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_85; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_86; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_87; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_88; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_89; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_90; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_91; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_92; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_93; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_94; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_95; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_96; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_97; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_98; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_99; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_100; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_101; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_102; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_103; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_104; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_105; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_106; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_107; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_108; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_109; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_110; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_111; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_112; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_113; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_114; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_115; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_116; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_117; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_118; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_119; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_120; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_121; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_122; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_123; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_124; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_125; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_126; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_127; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_128; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_129; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_130; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_131; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_132; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_133; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_134; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_135; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_136; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_137; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_138; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_139; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_140; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_141; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_142; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_143; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_144; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_145; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_146; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_147; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_148; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_149; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_150; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_151; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_152; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_153; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_154; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_155; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_156; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_157; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_158; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_159; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_160; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_161; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_162; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_163; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_164; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_165; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_166; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_167; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_168; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_169; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_170; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_171; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_172; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_173; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_174; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_175; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_176; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_177; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_178; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_179; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_180; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_181; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_182; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_183; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_184; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_185; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_186; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_187; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_188; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_189; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_190; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_191; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_192; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_193; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_194; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_195; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_196; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_197; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_198; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_199; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_200; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_201; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_202; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_203; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_204; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_205; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_206; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_207; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_208; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_209; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_210; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_211; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_212; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_213; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_214; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_215; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_216; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_217; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_218; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_219; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_220; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_221; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_222; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_223; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_224; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_225; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_226; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_227; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_228; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_229; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_230; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_231; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_232; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_233; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_234; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_235; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_236; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_237; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_238; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_239; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_240; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_241; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_242; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_243; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_244; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_245; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_246; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_247; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_248; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_249; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_250; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_251; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_252; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_253; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_254; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_255; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_256; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_257; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_258; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_259; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_260; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_261; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_262; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_263; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_264; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_265; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_266; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_267; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_268; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_269; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_270; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_271; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_272; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_273; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_274; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_275; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_276; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_277; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_278; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_279; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_280; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_281; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_282; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_283; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_284; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_285; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_286; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_287; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_288; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_289; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_290; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_291; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_292; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_293; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_294; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_295; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_296; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_297; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_298; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_299; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_300; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_301; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_302; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_303; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_304; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_305; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_306; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_307; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_308; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_309; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_310; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_311; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_312; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_313; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_314; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_315; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_316; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_317; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_318; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_319; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_320; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_321; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_322; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_323; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_324; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_325; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_326; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_327; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_328; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_329; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_330; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_331; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_332; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_333; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_334; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_335; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_336; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_337; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_338; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_339; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_340; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_341; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_342; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_343; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_344; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_345; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_346; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_347; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_348; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_349; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_350; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_351; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_352; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_353; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_354; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_355; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_356; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_357; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_358; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_359; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_360; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_361; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_362; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_363; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_364; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_365; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_366; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_367; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_368; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_369; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_370; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_371; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_372; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_373; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_374; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_375; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_376; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_377; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_378; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_379; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_380; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_381; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_382; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_383; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_384; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_385; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_386; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_387; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_388; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_389; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_390; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_391; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_392; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_393; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_394; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_395; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_396; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_397; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_398; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_399; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_400; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_401; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_402; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_403; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_404; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_405; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_406; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_407; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_408; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_409; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_410; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_411; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_412; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_413; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_414; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_415; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_416; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_417; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_418; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_419; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_420; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_421; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_422; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_423; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_424; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_425; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_426; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_427; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_428; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_429; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_430; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_431; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_432; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_433; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_434; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_435; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_436; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_437; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_438; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_439; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_440; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_441; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_442; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_443; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_444; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_445; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_446; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_447; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_448; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_449; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_450; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_451; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_452; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_453; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_454; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_455; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_456; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_457; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_458; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_459; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_460; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_461; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_462; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_463; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_464; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_465; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_466; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_467; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_468; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_469; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_470; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_471; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_472; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_473; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_474; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_475; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_476; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_477; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_478; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_479; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_480; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_481; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_482; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_483; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_484; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_485; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_486; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_487; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_488; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_489; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_490; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_491; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_492; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_493; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_494; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_495; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_496; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_497; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_498; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_499; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_500; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_501; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_502; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_503; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_504; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_505; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_506; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_507; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_508; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_509; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_510; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_511; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_0; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_1; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_2; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_3; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_4; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_5; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_6; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_7; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_8; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_9; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_10; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_11; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_12; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_13; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_14; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_15; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_parse_current_state; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 347:24]
  wire [3:0] pipe10_io_pipe_phv_out_next_processor_id; // @[matcher.scala 347:24]
  wire  pipe10_io_pipe_phv_out_next_config_id; // @[matcher.scala 347:24]
  wire  pipe10_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 347:24]
  wire [191:0] pipe10_io_key_in; // @[matcher.scala 347:24]
  wire [191:0] pipe10_io_key_out; // @[matcher.scala 347:24]
  wire [3:0] pipe10_io_cs_in; // @[matcher.scala 347:24]
  wire [3:0] pipe10_io_cs_out; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_addr_in; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_0; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_1; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_2; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_3; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_4; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_5; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_6; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_7; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_8; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_9; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_10; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_11; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_12; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_13; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_14; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_15; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_0; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_1; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_2; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_3; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_4; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_5; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_6; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_7; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_8; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_9; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_10; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_11; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_12; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_13; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_14; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_15; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_0_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_0_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_0_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_1_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_1_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_1_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_2_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_2_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_2_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_3_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_3_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_3_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_4_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_4_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_4_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_5_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_5_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_5_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_6_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_6_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_6_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_7_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_7_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_7_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_8_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_8_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_8_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_9_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_9_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_9_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_10_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_10_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_10_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_11_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_11_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_11_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_12_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_12_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_12_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_13_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_13_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_13_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_14_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_14_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_14_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_15_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_15_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_15_data; // @[matcher.scala 347:24]
  wire  pipe11_clock; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_0; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_1; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_2; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_3; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_4; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_5; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_6; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_7; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_8; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_9; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_10; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_11; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_12; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_13; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_14; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_15; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_16; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_17; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_18; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_19; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_20; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_21; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_22; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_23; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_24; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_25; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_26; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_27; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_28; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_29; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_30; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_31; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_32; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_33; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_34; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_35; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_36; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_37; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_38; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_39; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_40; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_41; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_42; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_43; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_44; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_45; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_46; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_47; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_48; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_49; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_50; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_51; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_52; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_53; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_54; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_55; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_56; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_57; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_58; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_59; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_60; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_61; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_62; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_63; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_64; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_65; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_66; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_67; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_68; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_69; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_70; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_71; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_72; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_73; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_74; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_75; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_76; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_77; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_78; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_79; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_80; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_81; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_82; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_83; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_84; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_85; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_86; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_87; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_88; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_89; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_90; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_91; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_92; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_93; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_94; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_95; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_96; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_97; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_98; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_99; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_100; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_101; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_102; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_103; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_104; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_105; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_106; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_107; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_108; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_109; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_110; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_111; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_112; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_113; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_114; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_115; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_116; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_117; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_118; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_119; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_120; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_121; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_122; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_123; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_124; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_125; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_126; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_127; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_128; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_129; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_130; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_131; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_132; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_133; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_134; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_135; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_136; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_137; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_138; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_139; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_140; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_141; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_142; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_143; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_144; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_145; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_146; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_147; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_148; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_149; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_150; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_151; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_152; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_153; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_154; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_155; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_156; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_157; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_158; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_159; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_160; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_161; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_162; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_163; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_164; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_165; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_166; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_167; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_168; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_169; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_170; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_171; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_172; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_173; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_174; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_175; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_176; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_177; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_178; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_179; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_180; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_181; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_182; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_183; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_184; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_185; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_186; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_187; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_188; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_189; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_190; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_191; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_192; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_193; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_194; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_195; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_196; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_197; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_198; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_199; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_200; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_201; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_202; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_203; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_204; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_205; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_206; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_207; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_208; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_209; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_210; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_211; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_212; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_213; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_214; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_215; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_216; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_217; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_218; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_219; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_220; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_221; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_222; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_223; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_224; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_225; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_226; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_227; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_228; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_229; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_230; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_231; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_232; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_233; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_234; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_235; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_236; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_237; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_238; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_239; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_240; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_241; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_242; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_243; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_244; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_245; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_246; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_247; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_248; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_249; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_250; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_251; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_252; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_253; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_254; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_255; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_256; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_257; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_258; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_259; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_260; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_261; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_262; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_263; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_264; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_265; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_266; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_267; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_268; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_269; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_270; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_271; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_272; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_273; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_274; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_275; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_276; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_277; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_278; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_279; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_280; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_281; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_282; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_283; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_284; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_285; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_286; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_287; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_288; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_289; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_290; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_291; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_292; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_293; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_294; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_295; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_296; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_297; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_298; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_299; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_300; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_301; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_302; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_303; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_304; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_305; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_306; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_307; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_308; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_309; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_310; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_311; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_312; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_313; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_314; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_315; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_316; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_317; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_318; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_319; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_320; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_321; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_322; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_323; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_324; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_325; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_326; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_327; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_328; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_329; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_330; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_331; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_332; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_333; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_334; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_335; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_336; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_337; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_338; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_339; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_340; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_341; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_342; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_343; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_344; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_345; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_346; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_347; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_348; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_349; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_350; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_351; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_352; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_353; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_354; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_355; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_356; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_357; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_358; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_359; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_360; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_361; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_362; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_363; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_364; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_365; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_366; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_367; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_368; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_369; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_370; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_371; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_372; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_373; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_374; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_375; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_376; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_377; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_378; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_379; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_380; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_381; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_382; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_383; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_384; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_385; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_386; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_387; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_388; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_389; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_390; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_391; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_392; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_393; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_394; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_395; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_396; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_397; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_398; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_399; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_400; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_401; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_402; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_403; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_404; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_405; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_406; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_407; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_408; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_409; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_410; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_411; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_412; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_413; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_414; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_415; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_416; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_417; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_418; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_419; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_420; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_421; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_422; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_423; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_424; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_425; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_426; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_427; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_428; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_429; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_430; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_431; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_432; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_433; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_434; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_435; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_436; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_437; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_438; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_439; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_440; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_441; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_442; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_443; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_444; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_445; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_446; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_447; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_448; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_449; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_450; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_451; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_452; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_453; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_454; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_455; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_456; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_457; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_458; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_459; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_460; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_461; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_462; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_463; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_464; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_465; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_466; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_467; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_468; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_469; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_470; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_471; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_472; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_473; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_474; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_475; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_476; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_477; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_478; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_479; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_480; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_481; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_482; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_483; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_484; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_485; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_486; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_487; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_488; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_489; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_490; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_491; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_492; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_493; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_494; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_495; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_496; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_497; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_498; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_499; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_500; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_501; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_502; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_503; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_504; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_505; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_506; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_507; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_508; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_509; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_510; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_511; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_0; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_1; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_2; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_3; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_4; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_5; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_6; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_7; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_8; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_9; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_10; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_11; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_12; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_13; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_14; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_15; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_parse_current_state; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 348:24]
  wire [3:0] pipe11_io_pipe_phv_in_next_processor_id; // @[matcher.scala 348:24]
  wire  pipe11_io_pipe_phv_in_next_config_id; // @[matcher.scala 348:24]
  wire  pipe11_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_0; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_1; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_2; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_3; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_4; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_5; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_6; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_7; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_8; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_9; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_10; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_11; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_12; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_13; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_14; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_15; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_16; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_17; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_18; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_19; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_20; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_21; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_22; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_23; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_24; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_25; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_26; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_27; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_28; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_29; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_30; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_31; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_32; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_33; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_34; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_35; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_36; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_37; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_38; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_39; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_40; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_41; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_42; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_43; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_44; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_45; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_46; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_47; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_48; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_49; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_50; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_51; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_52; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_53; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_54; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_55; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_56; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_57; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_58; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_59; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_60; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_61; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_62; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_63; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_64; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_65; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_66; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_67; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_68; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_69; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_70; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_71; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_72; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_73; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_74; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_75; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_76; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_77; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_78; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_79; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_80; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_81; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_82; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_83; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_84; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_85; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_86; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_87; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_88; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_89; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_90; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_91; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_92; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_93; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_94; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_95; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_96; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_97; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_98; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_99; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_100; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_101; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_102; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_103; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_104; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_105; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_106; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_107; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_108; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_109; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_110; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_111; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_112; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_113; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_114; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_115; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_116; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_117; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_118; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_119; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_120; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_121; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_122; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_123; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_124; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_125; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_126; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_127; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_128; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_129; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_130; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_131; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_132; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_133; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_134; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_135; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_136; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_137; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_138; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_139; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_140; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_141; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_142; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_143; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_144; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_145; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_146; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_147; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_148; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_149; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_150; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_151; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_152; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_153; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_154; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_155; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_156; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_157; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_158; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_159; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_160; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_161; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_162; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_163; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_164; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_165; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_166; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_167; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_168; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_169; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_170; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_171; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_172; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_173; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_174; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_175; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_176; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_177; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_178; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_179; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_180; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_181; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_182; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_183; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_184; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_185; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_186; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_187; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_188; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_189; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_190; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_191; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_192; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_193; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_194; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_195; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_196; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_197; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_198; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_199; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_200; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_201; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_202; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_203; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_204; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_205; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_206; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_207; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_208; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_209; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_210; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_211; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_212; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_213; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_214; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_215; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_216; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_217; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_218; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_219; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_220; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_221; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_222; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_223; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_224; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_225; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_226; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_227; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_228; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_229; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_230; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_231; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_232; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_233; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_234; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_235; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_236; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_237; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_238; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_239; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_240; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_241; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_242; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_243; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_244; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_245; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_246; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_247; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_248; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_249; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_250; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_251; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_252; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_253; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_254; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_255; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_256; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_257; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_258; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_259; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_260; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_261; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_262; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_263; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_264; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_265; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_266; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_267; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_268; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_269; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_270; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_271; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_272; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_273; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_274; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_275; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_276; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_277; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_278; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_279; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_280; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_281; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_282; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_283; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_284; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_285; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_286; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_287; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_288; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_289; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_290; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_291; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_292; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_293; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_294; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_295; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_296; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_297; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_298; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_299; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_300; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_301; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_302; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_303; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_304; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_305; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_306; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_307; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_308; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_309; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_310; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_311; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_312; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_313; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_314; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_315; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_316; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_317; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_318; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_319; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_320; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_321; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_322; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_323; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_324; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_325; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_326; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_327; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_328; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_329; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_330; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_331; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_332; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_333; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_334; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_335; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_336; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_337; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_338; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_339; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_340; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_341; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_342; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_343; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_344; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_345; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_346; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_347; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_348; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_349; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_350; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_351; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_352; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_353; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_354; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_355; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_356; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_357; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_358; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_359; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_360; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_361; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_362; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_363; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_364; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_365; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_366; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_367; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_368; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_369; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_370; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_371; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_372; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_373; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_374; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_375; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_376; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_377; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_378; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_379; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_380; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_381; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_382; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_383; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_384; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_385; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_386; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_387; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_388; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_389; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_390; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_391; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_392; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_393; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_394; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_395; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_396; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_397; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_398; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_399; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_400; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_401; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_402; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_403; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_404; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_405; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_406; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_407; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_408; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_409; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_410; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_411; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_412; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_413; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_414; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_415; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_416; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_417; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_418; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_419; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_420; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_421; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_422; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_423; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_424; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_425; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_426; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_427; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_428; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_429; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_430; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_431; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_432; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_433; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_434; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_435; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_436; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_437; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_438; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_439; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_440; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_441; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_442; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_443; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_444; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_445; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_446; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_447; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_448; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_449; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_450; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_451; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_452; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_453; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_454; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_455; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_456; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_457; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_458; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_459; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_460; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_461; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_462; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_463; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_464; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_465; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_466; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_467; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_468; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_469; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_470; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_471; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_472; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_473; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_474; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_475; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_476; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_477; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_478; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_479; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_480; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_481; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_482; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_483; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_484; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_485; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_486; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_487; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_488; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_489; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_490; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_491; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_492; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_493; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_494; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_495; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_496; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_497; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_498; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_499; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_500; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_501; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_502; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_503; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_504; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_505; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_506; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_507; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_508; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_509; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_510; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_511; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_0; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_1; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_2; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_3; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_4; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_5; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_6; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_7; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_8; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_9; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_10; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_11; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_12; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_13; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_14; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_15; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_parse_current_state; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 348:24]
  wire [3:0] pipe11_io_pipe_phv_out_next_processor_id; // @[matcher.scala 348:24]
  wire  pipe11_io_pipe_phv_out_next_config_id; // @[matcher.scala 348:24]
  wire  pipe11_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 348:24]
  wire [4:0] pipe11_io_table_config_0_table_width; // @[matcher.scala 348:24]
  wire [4:0] pipe11_io_table_config_0_table_depth; // @[matcher.scala 348:24]
  wire [4:0] pipe11_io_table_config_1_table_width; // @[matcher.scala 348:24]
  wire [4:0] pipe11_io_table_config_1_table_depth; // @[matcher.scala 348:24]
  wire [191:0] pipe11_io_key_in; // @[matcher.scala 348:24]
  wire [191:0] pipe11_io_key_out; // @[matcher.scala 348:24]
  wire [3:0] pipe11_io_cs_in; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_0; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_1; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_2; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_3; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_4; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_5; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_6; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_7; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_8; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_9; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_10; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_11; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_12; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_13; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_14; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_15; // @[matcher.scala 348:24]
  wire [255:0] pipe11_io_data_out; // @[matcher.scala 348:24]
  wire  pipe12_clock; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_0; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_1; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_2; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_3; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_4; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_5; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_6; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_7; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_8; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_9; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_10; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_11; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_12; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_13; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_14; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_15; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_16; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_17; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_18; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_19; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_20; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_21; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_22; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_23; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_24; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_25; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_26; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_27; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_28; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_29; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_30; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_31; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_32; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_33; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_34; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_35; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_36; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_37; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_38; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_39; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_40; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_41; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_42; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_43; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_44; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_45; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_46; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_47; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_48; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_49; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_50; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_51; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_52; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_53; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_54; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_55; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_56; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_57; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_58; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_59; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_60; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_61; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_62; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_63; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_64; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_65; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_66; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_67; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_68; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_69; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_70; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_71; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_72; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_73; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_74; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_75; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_76; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_77; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_78; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_79; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_80; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_81; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_82; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_83; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_84; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_85; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_86; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_87; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_88; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_89; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_90; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_91; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_92; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_93; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_94; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_95; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_96; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_97; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_98; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_99; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_100; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_101; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_102; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_103; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_104; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_105; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_106; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_107; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_108; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_109; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_110; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_111; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_112; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_113; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_114; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_115; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_116; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_117; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_118; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_119; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_120; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_121; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_122; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_123; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_124; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_125; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_126; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_127; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_128; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_129; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_130; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_131; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_132; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_133; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_134; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_135; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_136; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_137; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_138; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_139; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_140; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_141; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_142; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_143; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_144; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_145; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_146; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_147; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_148; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_149; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_150; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_151; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_152; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_153; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_154; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_155; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_156; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_157; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_158; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_159; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_160; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_161; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_162; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_163; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_164; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_165; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_166; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_167; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_168; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_169; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_170; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_171; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_172; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_173; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_174; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_175; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_176; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_177; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_178; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_179; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_180; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_181; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_182; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_183; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_184; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_185; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_186; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_187; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_188; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_189; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_190; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_191; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_192; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_193; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_194; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_195; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_196; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_197; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_198; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_199; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_200; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_201; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_202; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_203; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_204; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_205; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_206; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_207; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_208; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_209; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_210; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_211; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_212; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_213; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_214; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_215; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_216; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_217; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_218; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_219; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_220; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_221; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_222; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_223; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_224; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_225; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_226; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_227; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_228; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_229; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_230; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_231; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_232; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_233; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_234; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_235; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_236; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_237; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_238; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_239; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_240; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_241; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_242; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_243; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_244; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_245; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_246; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_247; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_248; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_249; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_250; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_251; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_252; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_253; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_254; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_255; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_256; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_257; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_258; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_259; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_260; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_261; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_262; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_263; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_264; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_265; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_266; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_267; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_268; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_269; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_270; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_271; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_272; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_273; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_274; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_275; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_276; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_277; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_278; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_279; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_280; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_281; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_282; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_283; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_284; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_285; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_286; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_287; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_288; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_289; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_290; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_291; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_292; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_293; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_294; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_295; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_296; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_297; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_298; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_299; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_300; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_301; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_302; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_303; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_304; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_305; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_306; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_307; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_308; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_309; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_310; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_311; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_312; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_313; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_314; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_315; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_316; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_317; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_318; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_319; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_320; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_321; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_322; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_323; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_324; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_325; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_326; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_327; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_328; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_329; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_330; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_331; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_332; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_333; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_334; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_335; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_336; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_337; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_338; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_339; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_340; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_341; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_342; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_343; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_344; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_345; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_346; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_347; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_348; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_349; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_350; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_351; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_352; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_353; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_354; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_355; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_356; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_357; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_358; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_359; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_360; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_361; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_362; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_363; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_364; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_365; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_366; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_367; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_368; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_369; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_370; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_371; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_372; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_373; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_374; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_375; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_376; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_377; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_378; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_379; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_380; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_381; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_382; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_383; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_384; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_385; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_386; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_387; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_388; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_389; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_390; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_391; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_392; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_393; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_394; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_395; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_396; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_397; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_398; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_399; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_400; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_401; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_402; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_403; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_404; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_405; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_406; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_407; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_408; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_409; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_410; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_411; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_412; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_413; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_414; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_415; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_416; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_417; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_418; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_419; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_420; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_421; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_422; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_423; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_424; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_425; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_426; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_427; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_428; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_429; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_430; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_431; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_432; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_433; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_434; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_435; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_436; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_437; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_438; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_439; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_440; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_441; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_442; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_443; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_444; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_445; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_446; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_447; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_448; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_449; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_450; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_451; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_452; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_453; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_454; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_455; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_456; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_457; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_458; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_459; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_460; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_461; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_462; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_463; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_464; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_465; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_466; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_467; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_468; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_469; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_470; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_471; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_472; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_473; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_474; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_475; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_476; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_477; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_478; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_479; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_480; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_481; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_482; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_483; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_484; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_485; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_486; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_487; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_488; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_489; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_490; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_491; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_492; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_493; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_494; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_495; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_496; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_497; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_498; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_499; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_500; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_501; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_502; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_503; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_504; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_505; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_506; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_507; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_508; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_509; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_510; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_511; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_0; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_1; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_2; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_3; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_4; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_5; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_6; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_7; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_8; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_9; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_10; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_11; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_12; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_13; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_14; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_15; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_parse_current_state; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 349:24]
  wire [3:0] pipe12_io_pipe_phv_in_next_processor_id; // @[matcher.scala 349:24]
  wire  pipe12_io_pipe_phv_in_next_config_id; // @[matcher.scala 349:24]
  wire  pipe12_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_0; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_1; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_2; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_3; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_4; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_5; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_6; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_7; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_8; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_9; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_10; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_11; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_12; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_13; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_14; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_15; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_16; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_17; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_18; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_19; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_20; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_21; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_22; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_23; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_24; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_25; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_26; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_27; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_28; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_29; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_30; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_31; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_32; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_33; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_34; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_35; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_36; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_37; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_38; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_39; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_40; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_41; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_42; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_43; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_44; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_45; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_46; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_47; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_48; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_49; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_50; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_51; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_52; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_53; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_54; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_55; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_56; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_57; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_58; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_59; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_60; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_61; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_62; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_63; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_64; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_65; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_66; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_67; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_68; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_69; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_70; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_71; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_72; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_73; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_74; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_75; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_76; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_77; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_78; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_79; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_80; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_81; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_82; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_83; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_84; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_85; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_86; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_87; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_88; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_89; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_90; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_91; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_92; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_93; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_94; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_95; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_96; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_97; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_98; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_99; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_100; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_101; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_102; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_103; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_104; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_105; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_106; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_107; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_108; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_109; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_110; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_111; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_112; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_113; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_114; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_115; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_116; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_117; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_118; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_119; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_120; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_121; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_122; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_123; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_124; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_125; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_126; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_127; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_128; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_129; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_130; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_131; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_132; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_133; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_134; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_135; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_136; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_137; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_138; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_139; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_140; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_141; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_142; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_143; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_144; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_145; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_146; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_147; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_148; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_149; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_150; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_151; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_152; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_153; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_154; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_155; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_156; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_157; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_158; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_159; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_160; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_161; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_162; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_163; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_164; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_165; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_166; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_167; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_168; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_169; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_170; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_171; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_172; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_173; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_174; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_175; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_176; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_177; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_178; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_179; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_180; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_181; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_182; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_183; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_184; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_185; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_186; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_187; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_188; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_189; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_190; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_191; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_192; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_193; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_194; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_195; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_196; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_197; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_198; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_199; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_200; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_201; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_202; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_203; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_204; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_205; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_206; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_207; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_208; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_209; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_210; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_211; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_212; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_213; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_214; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_215; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_216; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_217; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_218; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_219; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_220; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_221; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_222; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_223; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_224; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_225; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_226; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_227; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_228; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_229; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_230; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_231; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_232; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_233; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_234; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_235; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_236; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_237; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_238; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_239; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_240; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_241; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_242; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_243; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_244; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_245; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_246; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_247; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_248; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_249; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_250; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_251; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_252; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_253; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_254; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_255; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_256; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_257; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_258; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_259; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_260; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_261; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_262; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_263; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_264; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_265; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_266; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_267; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_268; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_269; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_270; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_271; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_272; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_273; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_274; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_275; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_276; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_277; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_278; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_279; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_280; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_281; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_282; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_283; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_284; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_285; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_286; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_287; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_288; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_289; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_290; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_291; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_292; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_293; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_294; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_295; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_296; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_297; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_298; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_299; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_300; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_301; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_302; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_303; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_304; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_305; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_306; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_307; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_308; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_309; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_310; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_311; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_312; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_313; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_314; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_315; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_316; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_317; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_318; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_319; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_320; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_321; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_322; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_323; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_324; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_325; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_326; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_327; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_328; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_329; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_330; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_331; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_332; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_333; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_334; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_335; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_336; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_337; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_338; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_339; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_340; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_341; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_342; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_343; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_344; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_345; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_346; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_347; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_348; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_349; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_350; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_351; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_352; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_353; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_354; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_355; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_356; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_357; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_358; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_359; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_360; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_361; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_362; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_363; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_364; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_365; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_366; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_367; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_368; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_369; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_370; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_371; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_372; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_373; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_374; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_375; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_376; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_377; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_378; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_379; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_380; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_381; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_382; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_383; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_384; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_385; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_386; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_387; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_388; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_389; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_390; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_391; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_392; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_393; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_394; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_395; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_396; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_397; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_398; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_399; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_400; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_401; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_402; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_403; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_404; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_405; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_406; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_407; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_408; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_409; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_410; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_411; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_412; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_413; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_414; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_415; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_416; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_417; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_418; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_419; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_420; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_421; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_422; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_423; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_424; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_425; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_426; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_427; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_428; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_429; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_430; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_431; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_432; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_433; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_434; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_435; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_436; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_437; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_438; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_439; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_440; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_441; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_442; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_443; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_444; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_445; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_446; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_447; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_448; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_449; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_450; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_451; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_452; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_453; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_454; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_455; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_456; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_457; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_458; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_459; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_460; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_461; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_462; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_463; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_464; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_465; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_466; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_467; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_468; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_469; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_470; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_471; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_472; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_473; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_474; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_475; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_476; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_477; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_478; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_479; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_480; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_481; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_482; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_483; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_484; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_485; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_486; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_487; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_488; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_489; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_490; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_491; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_492; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_493; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_494; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_495; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_496; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_497; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_498; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_499; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_500; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_501; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_502; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_503; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_504; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_505; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_506; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_507; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_508; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_509; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_510; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_511; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_0; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_1; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_2; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_3; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_4; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_5; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_6; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_7; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_8; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_9; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_10; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_11; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_12; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_13; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_14; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_15; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_parse_current_state; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 349:24]
  wire [3:0] pipe12_io_pipe_phv_out_next_processor_id; // @[matcher.scala 349:24]
  wire  pipe12_io_pipe_phv_out_next_config_id; // @[matcher.scala 349:24]
  wire  pipe12_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_key_config_0_key_length; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_key_config_1_key_length; // @[matcher.scala 349:24]
  wire [191:0] pipe12_io_key_in; // @[matcher.scala 349:24]
  wire [255:0] pipe12_io_data_in; // @[matcher.scala 349:24]
  wire  pipe12_io_hit; // @[matcher.scala 349:24]
  wire [63:0] pipe12_io_match_value; // @[matcher.scala 349:24]
  reg [7:0] key_config_0_header_id; // @[matcher.scala 17:25]
  reg [7:0] key_config_0_internal_offset; // @[matcher.scala 17:25]
  reg [7:0] key_config_0_key_length; // @[matcher.scala 17:25]
  reg [7:0] key_config_1_header_id; // @[matcher.scala 17:25]
  reg [7:0] key_config_1_internal_offset; // @[matcher.scala 17:25]
  reg [7:0] key_config_1_key_length; // @[matcher.scala 17:25]
  reg [4:0] table_config_0_table_width; // @[matcher.scala 18:27]
  reg [4:0] table_config_0_table_depth; // @[matcher.scala 18:27]
  reg [4:0] table_config_1_table_width; // @[matcher.scala 18:27]
  reg [4:0] table_config_1_table_depth; // @[matcher.scala 18:27]
  MatchGetOffset pipe1 ( // @[matcher.scala 343:23]
    .clock(pipe1_clock),
    .io_pipe_phv_in_data_0(pipe1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe1_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe1_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe1_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe1_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe1_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe1_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe1_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe1_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe1_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe1_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe1_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe1_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe1_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe1_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe1_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe1_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe1_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe1_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe1_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe1_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe1_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe1_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe1_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe1_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe1_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe1_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe1_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe1_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe1_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe1_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe1_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe1_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe1_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe1_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe1_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe1_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe1_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe1_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe1_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe1_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe1_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe1_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe1_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe1_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe1_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe1_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe1_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe1_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe1_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe1_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe1_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe1_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe1_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe1_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe1_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe1_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe1_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe1_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe1_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe1_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe1_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe1_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe1_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe1_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe1_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe1_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe1_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe1_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe1_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe1_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe1_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe1_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe1_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe1_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe1_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe1_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe1_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe1_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe1_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe1_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe1_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe1_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe1_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe1_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe1_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe1_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe1_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe1_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe1_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe1_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe1_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe1_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe1_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe1_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe1_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe1_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe1_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe1_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe1_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe1_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe1_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe1_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe1_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe1_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe1_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe1_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe1_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe1_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe1_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe1_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe1_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe1_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe1_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe1_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe1_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe1_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe1_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe1_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe1_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe1_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe1_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe1_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe1_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe1_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe1_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe1_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe1_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe1_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe1_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe1_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe1_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe1_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe1_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe1_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe1_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe1_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe1_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe1_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe1_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe1_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe1_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe1_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe1_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe1_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe1_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe1_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe1_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe1_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe1_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe1_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe1_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe1_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe1_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe1_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe1_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe1_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe1_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe1_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe1_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe1_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe1_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe1_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe1_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe1_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe1_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe1_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe1_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe1_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe1_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe1_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe1_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe1_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe1_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe1_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe1_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe1_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe1_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe1_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe1_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe1_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe1_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe1_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe1_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe1_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe1_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe1_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe1_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe1_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe1_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe1_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe1_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe1_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe1_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe1_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe1_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe1_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe1_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe1_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe1_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe1_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe1_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe1_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe1_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe1_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe1_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe1_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe1_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe1_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe1_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe1_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe1_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe1_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe1_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe1_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe1_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe1_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe1_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe1_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe1_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe1_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe1_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe1_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe1_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe1_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe1_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe1_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe1_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe1_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe1_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe1_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe1_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe1_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe1_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe1_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe1_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe1_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe1_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe1_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe1_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe1_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe1_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe1_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe1_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe1_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe1_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe1_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe1_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe1_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe1_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe1_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe1_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe1_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe1_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe1_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe1_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe1_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe1_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe1_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe1_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe1_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe1_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe1_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe1_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe1_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe1_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe1_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe1_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe1_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe1_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe1_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe1_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe1_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe1_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe1_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe1_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe1_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe1_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe1_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe1_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe1_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe1_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe1_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe1_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe1_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe1_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe1_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe1_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe1_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe1_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe1_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe1_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe1_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe1_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe1_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe1_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe1_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe1_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe1_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe1_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe1_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe1_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe1_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe1_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe1_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe1_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe1_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe1_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe1_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe1_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe1_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe1_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe1_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe1_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe1_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe1_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe1_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe1_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe1_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe1_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe1_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe1_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe1_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe1_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe1_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe1_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe1_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe1_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe1_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe1_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe1_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe1_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe1_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe1_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe1_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe1_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe1_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe1_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe1_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe1_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe1_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe1_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe1_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe1_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe1_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe1_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe1_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe1_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe1_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe1_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe1_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe1_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe1_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe1_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe1_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe1_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe1_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe1_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe1_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe1_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe1_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe1_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe1_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe1_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe1_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe1_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe1_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe1_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe1_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe1_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe1_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe1_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe1_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe1_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe1_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe1_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe1_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe1_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe1_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe1_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe1_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe1_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe1_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe1_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe1_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe1_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe1_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe1_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe1_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe1_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe1_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe1_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe1_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe1_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe1_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe1_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe1_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe1_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe1_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe1_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe1_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe1_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe1_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe1_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe1_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe1_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe1_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe1_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe1_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe1_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe1_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe1_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe1_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe1_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe1_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe1_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe1_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe1_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe1_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe1_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe1_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe1_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe1_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe1_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe1_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe1_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe1_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe1_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe1_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe1_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe1_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe1_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe1_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe1_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe1_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe1_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe1_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe1_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe1_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe1_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe1_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe1_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe1_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe1_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe1_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe1_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe1_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe1_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe1_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe1_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe1_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe1_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe1_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe1_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe1_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe1_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe1_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe1_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe1_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe1_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe1_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe1_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe1_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe1_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe1_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe1_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe1_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe1_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe1_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe1_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe1_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe1_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe1_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe1_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe1_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe1_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe1_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe1_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe1_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe1_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe1_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe1_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe1_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe1_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe1_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe1_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe1_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe1_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe1_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe1_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe1_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe1_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe1_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe1_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe1_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe1_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe1_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe1_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe1_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe1_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe1_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe1_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe1_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe1_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe1_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe1_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe1_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe1_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe1_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe1_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe1_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe1_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe1_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe1_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe1_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe1_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe1_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe1_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe1_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe1_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe1_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe1_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe1_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe1_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe1_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe1_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe1_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe1_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe1_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe1_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe1_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe1_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe1_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe1_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe1_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe1_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe1_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe1_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe1_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe1_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe1_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe1_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe1_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe1_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe1_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe1_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe1_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe1_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe1_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe1_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe1_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe1_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe1_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe1_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe1_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe1_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe1_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe1_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe1_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe1_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe1_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe1_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe1_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe1_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe1_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe1_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe1_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe1_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe1_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe1_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe1_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe1_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe1_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe1_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe1_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe1_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe1_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe1_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe1_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe1_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe1_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe1_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe1_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe1_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe1_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe1_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe1_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe1_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe1_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe1_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe1_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe1_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe1_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe1_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe1_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe1_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe1_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe1_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe1_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe1_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe1_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe1_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe1_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe1_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe1_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe1_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe1_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe1_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe1_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe1_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe1_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe1_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe1_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe1_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe1_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe1_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe1_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe1_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe1_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe1_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe1_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe1_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe1_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe1_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe1_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe1_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe1_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe1_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe1_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe1_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe1_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe1_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe1_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe1_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe1_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe1_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe1_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe1_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe1_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe1_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe1_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe1_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe1_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe1_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe1_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe1_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe1_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe1_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe1_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe1_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe1_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe1_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe1_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe1_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe1_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe1_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe1_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe1_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe1_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe1_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe1_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe1_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe1_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe1_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe1_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe1_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe1_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe1_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe1_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe1_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe1_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe1_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe1_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe1_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe1_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe1_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe1_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe1_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe1_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe1_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe1_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe1_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe1_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe1_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe1_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe1_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe1_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe1_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe1_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe1_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe1_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe1_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe1_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe1_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe1_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe1_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe1_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe1_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe1_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe1_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe1_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe1_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe1_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe1_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe1_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe1_io_pipe_phv_out_is_valid_processor),
    .io_key_config_0_header_id(pipe1_io_key_config_0_header_id),
    .io_key_config_0_internal_offset(pipe1_io_key_config_0_internal_offset),
    .io_key_config_1_header_id(pipe1_io_key_config_1_header_id),
    .io_key_config_1_internal_offset(pipe1_io_key_config_1_internal_offset),
    .io_key_offset(pipe1_io_key_offset)
  );
  MatchGetKey pipe2 ( // @[matcher.scala 344:23]
    .clock(pipe2_clock),
    .io_pipe_phv_in_data_0(pipe2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe2_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe2_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe2_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe2_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe2_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe2_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe2_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe2_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe2_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe2_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe2_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe2_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe2_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe2_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe2_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe2_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe2_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe2_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe2_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe2_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe2_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe2_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe2_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe2_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe2_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe2_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe2_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe2_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe2_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe2_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe2_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe2_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe2_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe2_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe2_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe2_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe2_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe2_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe2_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe2_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe2_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe2_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe2_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe2_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe2_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe2_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe2_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe2_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe2_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe2_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe2_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe2_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe2_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe2_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe2_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe2_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe2_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe2_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe2_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe2_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe2_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe2_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe2_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe2_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe2_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe2_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe2_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe2_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe2_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe2_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe2_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe2_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe2_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe2_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe2_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe2_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe2_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe2_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe2_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe2_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe2_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe2_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe2_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe2_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe2_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe2_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe2_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe2_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe2_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe2_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe2_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe2_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe2_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe2_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe2_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe2_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe2_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe2_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe2_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe2_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe2_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe2_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe2_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe2_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe2_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe2_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe2_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe2_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe2_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe2_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe2_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe2_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe2_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe2_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe2_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe2_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe2_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe2_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe2_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe2_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe2_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe2_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe2_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe2_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe2_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe2_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe2_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe2_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe2_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe2_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe2_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe2_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe2_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe2_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe2_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe2_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe2_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe2_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe2_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe2_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe2_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe2_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe2_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe2_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe2_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe2_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe2_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe2_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe2_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe2_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe2_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe2_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe2_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe2_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe2_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe2_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe2_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe2_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe2_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe2_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe2_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe2_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe2_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe2_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe2_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe2_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe2_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe2_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe2_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe2_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe2_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe2_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe2_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe2_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe2_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe2_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe2_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe2_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe2_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe2_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe2_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe2_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe2_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe2_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe2_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe2_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe2_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe2_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe2_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe2_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe2_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe2_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe2_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe2_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe2_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe2_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe2_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe2_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe2_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe2_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe2_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe2_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe2_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe2_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe2_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe2_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe2_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe2_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe2_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe2_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe2_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe2_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe2_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe2_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe2_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe2_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe2_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe2_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe2_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe2_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe2_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe2_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe2_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe2_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe2_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe2_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe2_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe2_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe2_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe2_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe2_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe2_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe2_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe2_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe2_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe2_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe2_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe2_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe2_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe2_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe2_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe2_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe2_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe2_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe2_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe2_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe2_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe2_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe2_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe2_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe2_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe2_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe2_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe2_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe2_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe2_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe2_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe2_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe2_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe2_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe2_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe2_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe2_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe2_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe2_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe2_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe2_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe2_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe2_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe2_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe2_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe2_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe2_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe2_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe2_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe2_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe2_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe2_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe2_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe2_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe2_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe2_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe2_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe2_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe2_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe2_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe2_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe2_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe2_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe2_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe2_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe2_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe2_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe2_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe2_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe2_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe2_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe2_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe2_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe2_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe2_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe2_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe2_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe2_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe2_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe2_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe2_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe2_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe2_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe2_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe2_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe2_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe2_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe2_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe2_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe2_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe2_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe2_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe2_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe2_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe2_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe2_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe2_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe2_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe2_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe2_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe2_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe2_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe2_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe2_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe2_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe2_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe2_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe2_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe2_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe2_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe2_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe2_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe2_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe2_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe2_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe2_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe2_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe2_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe2_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe2_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe2_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe2_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe2_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe2_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe2_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe2_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe2_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe2_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe2_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe2_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe2_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe2_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe2_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe2_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe2_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe2_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe2_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe2_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe2_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe2_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe2_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe2_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe2_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe2_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe2_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe2_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe2_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe2_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe2_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe2_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe2_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe2_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe2_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe2_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe2_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe2_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe2_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe2_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe2_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe2_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe2_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe2_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe2_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe2_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe2_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe2_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe2_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe2_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe2_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe2_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe2_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe2_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe2_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe2_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe2_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe2_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe2_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe2_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe2_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe2_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe2_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe2_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe2_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe2_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe2_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe2_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe2_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe2_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe2_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe2_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe2_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe2_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe2_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe2_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe2_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe2_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe2_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe2_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe2_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe2_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe2_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe2_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe2_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe2_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe2_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe2_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe2_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe2_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe2_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe2_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe2_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe2_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe2_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe2_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe2_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe2_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe2_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe2_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe2_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe2_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe2_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe2_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe2_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe2_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe2_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe2_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe2_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe2_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe2_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe2_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe2_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe2_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe2_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe2_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe2_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe2_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe2_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe2_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe2_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe2_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe2_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe2_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe2_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe2_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe2_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe2_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe2_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe2_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe2_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe2_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe2_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe2_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe2_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe2_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe2_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe2_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe2_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe2_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe2_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe2_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe2_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe2_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe2_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe2_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe2_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe2_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe2_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe2_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe2_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe2_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe2_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe2_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe2_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe2_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe2_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe2_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe2_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe2_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe2_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe2_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe2_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe2_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe2_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe2_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe2_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe2_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe2_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe2_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe2_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe2_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe2_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe2_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe2_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe2_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe2_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe2_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe2_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe2_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe2_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe2_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe2_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe2_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe2_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe2_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe2_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe2_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe2_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe2_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe2_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe2_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe2_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe2_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe2_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe2_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe2_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe2_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe2_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe2_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe2_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe2_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe2_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe2_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe2_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe2_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe2_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe2_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe2_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe2_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe2_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe2_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe2_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe2_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe2_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe2_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe2_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe2_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe2_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe2_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe2_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe2_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe2_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe2_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe2_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe2_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe2_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe2_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe2_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe2_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe2_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe2_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe2_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe2_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe2_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe2_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe2_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe2_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe2_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe2_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe2_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe2_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe2_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe2_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe2_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe2_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe2_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe2_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe2_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe2_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe2_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe2_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe2_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe2_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe2_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe2_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe2_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe2_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe2_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe2_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe2_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe2_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe2_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe2_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe2_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe2_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe2_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe2_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe2_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe2_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe2_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe2_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe2_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe2_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe2_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe2_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe2_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe2_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe2_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe2_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe2_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe2_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe2_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe2_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe2_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe2_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe2_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe2_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe2_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe2_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe2_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe2_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe2_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe2_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe2_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe2_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe2_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe2_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe2_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe2_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe2_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe2_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe2_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe2_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe2_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe2_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe2_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe2_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe2_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe2_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe2_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe2_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe2_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe2_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe2_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe2_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe2_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe2_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe2_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe2_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe2_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe2_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe2_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe2_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe2_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe2_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe2_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe2_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe2_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe2_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe2_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe2_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe2_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe2_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe2_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe2_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe2_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe2_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe2_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe2_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe2_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe2_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe2_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe2_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe2_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe2_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe2_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe2_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe2_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe2_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe2_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe2_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe2_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe2_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe2_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe2_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe2_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe2_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe2_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe2_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe2_io_pipe_phv_out_is_valid_processor),
    .io_key_config_0_key_length(pipe2_io_key_config_0_key_length),
    .io_key_config_1_key_length(pipe2_io_key_config_1_key_length),
    .io_key_offset(pipe2_io_key_offset),
    .io_match_key(pipe2_io_match_key)
  );
  Hash pipe3to8 ( // @[matcher.scala 345:26]
    .clock(pipe3to8_clock),
    .io_pipe_phv_in_data_0(pipe3to8_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe3to8_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe3to8_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe3to8_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe3to8_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe3to8_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe3to8_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe3to8_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe3to8_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe3to8_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe3to8_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe3to8_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe3to8_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe3to8_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe3to8_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe3to8_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe3to8_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe3to8_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe3to8_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe3to8_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe3to8_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe3to8_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe3to8_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe3to8_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe3to8_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe3to8_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe3to8_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe3to8_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe3to8_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe3to8_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe3to8_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe3to8_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe3to8_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe3to8_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe3to8_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe3to8_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe3to8_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe3to8_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe3to8_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe3to8_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe3to8_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe3to8_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe3to8_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe3to8_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe3to8_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe3to8_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe3to8_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe3to8_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe3to8_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe3to8_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe3to8_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe3to8_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe3to8_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe3to8_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe3to8_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe3to8_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe3to8_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe3to8_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe3to8_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe3to8_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe3to8_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe3to8_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe3to8_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe3to8_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe3to8_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe3to8_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe3to8_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe3to8_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe3to8_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe3to8_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe3to8_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe3to8_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe3to8_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe3to8_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe3to8_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe3to8_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe3to8_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe3to8_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe3to8_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe3to8_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe3to8_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe3to8_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe3to8_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe3to8_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe3to8_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe3to8_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe3to8_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe3to8_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe3to8_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe3to8_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe3to8_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe3to8_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe3to8_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe3to8_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe3to8_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe3to8_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe3to8_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe3to8_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe3to8_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe3to8_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe3to8_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe3to8_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe3to8_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe3to8_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe3to8_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe3to8_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe3to8_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe3to8_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe3to8_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe3to8_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe3to8_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe3to8_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe3to8_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe3to8_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe3to8_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe3to8_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe3to8_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe3to8_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe3to8_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe3to8_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe3to8_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe3to8_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe3to8_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe3to8_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe3to8_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe3to8_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe3to8_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe3to8_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe3to8_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe3to8_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe3to8_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe3to8_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe3to8_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe3to8_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe3to8_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe3to8_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe3to8_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe3to8_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe3to8_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe3to8_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe3to8_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe3to8_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe3to8_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe3to8_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe3to8_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe3to8_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe3to8_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe3to8_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe3to8_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe3to8_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe3to8_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe3to8_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe3to8_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe3to8_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe3to8_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe3to8_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe3to8_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe3to8_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe3to8_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe3to8_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe3to8_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe3to8_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe3to8_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe3to8_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe3to8_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe3to8_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe3to8_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe3to8_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe3to8_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe3to8_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe3to8_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe3to8_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe3to8_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe3to8_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe3to8_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe3to8_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe3to8_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe3to8_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe3to8_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe3to8_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe3to8_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe3to8_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe3to8_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe3to8_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe3to8_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe3to8_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe3to8_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe3to8_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe3to8_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe3to8_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe3to8_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe3to8_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe3to8_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe3to8_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe3to8_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe3to8_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe3to8_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe3to8_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe3to8_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe3to8_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe3to8_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe3to8_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe3to8_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe3to8_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe3to8_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe3to8_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe3to8_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe3to8_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe3to8_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe3to8_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe3to8_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe3to8_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe3to8_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe3to8_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe3to8_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe3to8_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe3to8_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe3to8_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe3to8_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe3to8_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe3to8_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe3to8_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe3to8_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe3to8_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe3to8_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe3to8_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe3to8_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe3to8_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe3to8_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe3to8_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe3to8_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe3to8_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe3to8_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe3to8_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe3to8_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe3to8_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe3to8_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe3to8_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe3to8_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe3to8_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe3to8_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe3to8_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe3to8_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe3to8_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe3to8_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe3to8_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe3to8_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe3to8_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe3to8_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe3to8_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe3to8_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe3to8_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe3to8_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe3to8_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe3to8_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe3to8_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe3to8_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe3to8_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe3to8_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe3to8_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe3to8_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe3to8_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe3to8_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe3to8_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe3to8_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe3to8_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe3to8_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe3to8_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe3to8_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe3to8_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe3to8_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe3to8_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe3to8_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe3to8_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe3to8_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe3to8_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe3to8_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe3to8_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe3to8_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe3to8_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe3to8_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe3to8_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe3to8_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe3to8_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe3to8_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe3to8_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe3to8_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe3to8_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe3to8_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe3to8_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe3to8_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe3to8_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe3to8_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe3to8_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe3to8_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe3to8_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe3to8_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe3to8_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe3to8_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe3to8_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe3to8_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe3to8_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe3to8_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe3to8_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe3to8_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe3to8_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe3to8_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe3to8_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe3to8_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe3to8_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe3to8_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe3to8_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe3to8_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe3to8_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe3to8_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe3to8_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe3to8_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe3to8_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe3to8_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe3to8_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe3to8_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe3to8_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe3to8_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe3to8_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe3to8_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe3to8_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe3to8_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe3to8_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe3to8_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe3to8_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe3to8_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe3to8_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe3to8_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe3to8_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe3to8_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe3to8_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe3to8_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe3to8_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe3to8_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe3to8_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe3to8_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe3to8_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe3to8_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe3to8_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe3to8_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe3to8_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe3to8_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe3to8_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe3to8_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe3to8_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe3to8_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe3to8_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe3to8_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe3to8_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe3to8_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe3to8_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe3to8_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe3to8_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe3to8_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe3to8_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe3to8_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe3to8_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe3to8_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe3to8_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe3to8_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe3to8_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe3to8_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe3to8_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe3to8_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe3to8_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe3to8_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe3to8_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe3to8_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe3to8_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe3to8_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe3to8_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe3to8_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe3to8_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe3to8_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe3to8_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe3to8_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe3to8_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe3to8_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe3to8_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe3to8_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe3to8_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe3to8_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe3to8_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe3to8_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe3to8_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe3to8_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe3to8_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe3to8_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe3to8_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe3to8_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe3to8_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe3to8_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe3to8_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe3to8_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe3to8_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe3to8_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe3to8_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe3to8_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe3to8_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe3to8_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe3to8_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe3to8_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe3to8_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe3to8_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe3to8_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe3to8_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe3to8_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe3to8_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe3to8_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe3to8_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe3to8_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe3to8_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe3to8_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe3to8_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe3to8_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe3to8_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe3to8_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe3to8_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe3to8_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe3to8_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe3to8_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe3to8_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe3to8_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe3to8_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe3to8_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe3to8_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe3to8_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe3to8_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe3to8_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe3to8_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe3to8_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe3to8_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe3to8_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe3to8_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe3to8_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe3to8_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe3to8_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe3to8_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe3to8_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe3to8_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe3to8_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe3to8_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe3to8_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe3to8_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe3to8_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe3to8_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe3to8_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe3to8_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe3to8_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe3to8_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe3to8_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe3to8_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe3to8_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe3to8_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe3to8_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe3to8_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe3to8_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe3to8_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe3to8_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe3to8_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe3to8_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe3to8_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe3to8_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe3to8_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe3to8_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe3to8_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe3to8_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe3to8_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe3to8_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe3to8_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe3to8_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe3to8_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe3to8_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe3to8_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe3to8_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe3to8_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe3to8_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe3to8_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe3to8_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe3to8_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe3to8_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe3to8_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe3to8_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe3to8_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe3to8_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe3to8_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe3to8_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe3to8_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe3to8_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe3to8_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe3to8_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe3to8_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe3to8_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe3to8_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe3to8_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe3to8_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe3to8_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe3to8_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe3to8_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe3to8_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe3to8_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe3to8_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe3to8_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe3to8_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe3to8_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe3to8_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe3to8_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe3to8_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe3to8_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe3to8_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe3to8_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe3to8_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe3to8_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe3to8_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe3to8_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe3to8_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe3to8_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe3to8_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe3to8_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe3to8_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe3to8_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe3to8_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe3to8_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe3to8_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe3to8_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe3to8_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe3to8_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe3to8_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe3to8_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe3to8_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe3to8_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe3to8_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe3to8_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe3to8_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe3to8_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe3to8_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe3to8_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe3to8_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe3to8_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe3to8_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe3to8_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe3to8_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe3to8_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe3to8_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe3to8_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe3to8_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe3to8_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe3to8_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe3to8_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe3to8_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe3to8_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe3to8_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe3to8_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe3to8_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe3to8_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe3to8_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe3to8_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe3to8_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe3to8_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe3to8_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe3to8_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe3to8_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe3to8_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe3to8_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe3to8_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe3to8_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe3to8_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe3to8_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe3to8_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe3to8_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe3to8_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe3to8_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe3to8_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe3to8_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe3to8_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe3to8_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe3to8_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe3to8_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe3to8_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe3to8_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe3to8_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe3to8_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe3to8_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe3to8_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe3to8_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe3to8_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe3to8_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe3to8_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe3to8_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe3to8_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe3to8_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe3to8_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe3to8_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe3to8_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe3to8_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe3to8_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe3to8_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe3to8_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe3to8_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe3to8_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe3to8_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe3to8_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe3to8_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe3to8_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe3to8_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe3to8_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe3to8_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe3to8_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe3to8_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe3to8_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe3to8_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe3to8_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe3to8_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe3to8_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe3to8_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe3to8_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe3to8_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe3to8_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe3to8_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe3to8_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe3to8_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe3to8_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe3to8_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe3to8_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe3to8_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe3to8_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe3to8_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe3to8_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe3to8_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe3to8_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe3to8_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe3to8_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe3to8_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe3to8_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe3to8_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe3to8_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe3to8_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe3to8_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe3to8_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe3to8_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe3to8_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe3to8_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe3to8_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe3to8_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe3to8_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe3to8_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe3to8_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe3to8_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe3to8_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe3to8_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe3to8_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe3to8_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe3to8_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe3to8_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe3to8_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe3to8_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe3to8_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe3to8_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe3to8_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe3to8_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe3to8_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe3to8_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe3to8_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe3to8_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe3to8_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe3to8_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe3to8_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe3to8_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe3to8_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe3to8_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe3to8_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe3to8_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe3to8_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe3to8_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe3to8_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe3to8_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe3to8_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe3to8_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe3to8_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe3to8_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe3to8_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe3to8_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe3to8_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe3to8_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe3to8_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe3to8_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe3to8_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe3to8_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe3to8_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe3to8_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe3to8_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe3to8_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe3to8_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe3to8_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe3to8_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe3to8_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe3to8_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe3to8_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe3to8_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe3to8_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe3to8_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe3to8_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe3to8_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe3to8_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe3to8_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe3to8_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe3to8_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe3to8_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe3to8_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe3to8_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe3to8_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe3to8_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe3to8_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe3to8_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe3to8_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe3to8_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe3to8_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe3to8_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe3to8_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe3to8_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe3to8_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe3to8_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe3to8_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe3to8_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe3to8_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe3to8_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe3to8_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe3to8_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe3to8_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe3to8_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe3to8_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe3to8_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe3to8_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe3to8_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe3to8_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe3to8_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe3to8_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe3to8_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe3to8_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe3to8_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe3to8_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe3to8_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe3to8_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe3to8_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe3to8_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe3to8_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe3to8_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe3to8_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe3to8_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe3to8_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe3to8_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe3to8_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe3to8_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe3to8_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe3to8_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe3to8_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe3to8_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe3to8_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe3to8_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe3to8_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe3to8_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe3to8_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe3to8_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe3to8_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe3to8_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe3to8_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe3to8_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe3to8_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe3to8_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe3to8_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe3to8_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe3to8_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe3to8_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe3to8_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe3to8_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe3to8_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe3to8_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe3to8_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe3to8_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe3to8_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe3to8_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe3to8_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe3to8_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe3to8_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe3to8_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe3to8_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe3to8_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe3to8_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe3to8_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe3to8_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe3to8_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe3to8_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe3to8_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe3to8_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe3to8_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe3to8_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe3to8_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe3to8_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe3to8_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe3to8_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe3to8_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe3to8_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe3to8_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe3to8_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe3to8_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe3to8_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe3to8_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe3to8_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe3to8_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe3to8_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe3to8_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe3to8_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe3to8_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe3to8_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe3to8_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe3to8_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe3to8_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe3to8_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe3to8_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe3to8_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe3to8_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe3to8_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe3to8_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe3to8_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe3to8_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe3to8_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe3to8_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe3to8_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe3to8_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe3to8_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe3to8_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe3to8_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe3to8_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe3to8_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe3to8_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe3to8_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe3to8_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe3to8_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe3to8_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe3to8_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe3to8_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe3to8_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe3to8_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe3to8_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe3to8_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe3to8_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe3to8_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe3to8_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe3to8_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe3to8_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe3to8_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe3to8_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe3to8_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe3to8_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe3to8_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe3to8_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe3to8_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe3to8_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe3to8_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe3to8_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe3to8_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe3to8_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe3to8_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe3to8_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe3to8_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe3to8_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe3to8_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe3to8_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe3to8_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe3to8_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe3to8_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe3to8_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe3to8_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe3to8_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe3to8_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe3to8_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe3to8_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe3to8_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe3to8_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe3to8_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe3to8_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe3to8_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe3to8_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe3to8_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe3to8_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe3to8_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe3to8_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe3to8_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe3to8_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe3to8_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe3to8_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe3to8_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe3to8_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe3to8_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe3to8_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe3to8_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe3to8_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe3to8_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe3to8_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe3to8_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe3to8_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe3to8_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe3to8_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe3to8_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe3to8_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe3to8_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe3to8_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe3to8_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe3to8_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe3to8_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe3to8_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe3to8_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe3to8_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe3to8_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe3to8_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe3to8_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe3to8_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe3to8_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe3to8_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe3to8_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe3to8_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe3to8_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe3to8_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe3to8_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe3to8_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe3to8_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe3to8_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe3to8_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe3to8_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe3to8_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe3to8_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe3to8_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe3to8_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe3to8_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe3to8_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe3to8_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe3to8_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe3to8_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe3to8_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe3to8_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe3to8_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe3to8_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe3to8_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe3to8_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe3to8_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe3to8_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe3to8_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe3to8_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe3to8_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe3to8_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe3to8_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe3to8_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe3to8_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe3to8_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe3to8_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe3to8_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe3to8_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe3to8_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe3to8_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe3to8_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe3to8_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe3to8_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe3to8_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe3to8_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe3to8_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe3to8_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe3to8_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe3to8_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe3to8_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe3to8_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe3to8_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe3to8_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe3to8_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe3to8_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe3to8_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe3to8_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe3to8_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe3to8_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe3to8_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe3to8_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe3to8_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe3to8_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe3to8_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe3to8_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe3to8_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe3to8_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe3to8_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe3to8_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe3to8_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe3to8_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe3to8_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe3to8_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe3to8_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe3to8_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe3to8_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe3to8_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe3to8_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe3to8_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe3to8_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe3to8_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe3to8_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe3to8_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe3to8_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe3to8_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe3to8_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe3to8_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe3to8_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe3to8_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe3to8_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe3to8_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe3to8_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe3to8_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe3to8_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe3to8_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe3to8_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe3to8_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe3to8_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe3to8_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe3to8_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe3to8_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe3to8_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe3to8_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe3to8_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe3to8_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe3to8_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe3to8_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe3to8_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe3to8_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe3to8_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe3to8_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe3to8_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe3to8_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe3to8_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe3to8_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe3to8_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe3to8_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe3to8_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe3to8_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe3to8_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe3to8_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe3to8_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe3to8_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe3to8_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe3to8_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe3to8_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe3to8_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe3to8_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe3to8_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe3to8_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe3to8_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe3to8_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe3to8_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe3to8_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe3to8_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe3to8_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe3to8_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe3to8_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe3to8_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe3to8_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe3to8_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe3to8_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe3to8_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe3to8_io_pipe_phv_out_is_valid_processor),
    .io_mod_hash_depth_mod(pipe3to8_io_mod_hash_depth_mod),
    .io_mod_config_id(pipe3to8_io_mod_config_id),
    .io_mod_hash_depth(pipe3to8_io_mod_hash_depth),
    .io_key_in(pipe3to8_io_key_in),
    .io_key_out(pipe3to8_io_key_out),
    .io_hash_val(pipe3to8_io_hash_val),
    .io_hash_val_cs(pipe3to8_io_hash_val_cs)
  );
  MatchGetCs pipe9 ( // @[matcher.scala 346:23]
    .clock(pipe9_clock),
    .io_pipe_phv_in_data_0(pipe9_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe9_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe9_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe9_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe9_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe9_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe9_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe9_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe9_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe9_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe9_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe9_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe9_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe9_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe9_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe9_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe9_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe9_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe9_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe9_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe9_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe9_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe9_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe9_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe9_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe9_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe9_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe9_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe9_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe9_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe9_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe9_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe9_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe9_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe9_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe9_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe9_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe9_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe9_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe9_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe9_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe9_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe9_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe9_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe9_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe9_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe9_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe9_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe9_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe9_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe9_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe9_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe9_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe9_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe9_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe9_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe9_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe9_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe9_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe9_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe9_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe9_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe9_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe9_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe9_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe9_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe9_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe9_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe9_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe9_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe9_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe9_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe9_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe9_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe9_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe9_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe9_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe9_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe9_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe9_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe9_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe9_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe9_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe9_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe9_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe9_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe9_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe9_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe9_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe9_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe9_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe9_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe9_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe9_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe9_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe9_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe9_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe9_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe9_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe9_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe9_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe9_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe9_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe9_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe9_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe9_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe9_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe9_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe9_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe9_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe9_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe9_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe9_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe9_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe9_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe9_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe9_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe9_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe9_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe9_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe9_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe9_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe9_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe9_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe9_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe9_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe9_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe9_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe9_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe9_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe9_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe9_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe9_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe9_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe9_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe9_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe9_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe9_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe9_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe9_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe9_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe9_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe9_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe9_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe9_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe9_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe9_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe9_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe9_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe9_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe9_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe9_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe9_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe9_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe9_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe9_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe9_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe9_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe9_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe9_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe9_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe9_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe9_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe9_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe9_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe9_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe9_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe9_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe9_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe9_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe9_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe9_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe9_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe9_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe9_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe9_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe9_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe9_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe9_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe9_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe9_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe9_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe9_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe9_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe9_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe9_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe9_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe9_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe9_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe9_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe9_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe9_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe9_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe9_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe9_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe9_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe9_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe9_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe9_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe9_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe9_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe9_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe9_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe9_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe9_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe9_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe9_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe9_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe9_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe9_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe9_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe9_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe9_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe9_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe9_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe9_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe9_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe9_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe9_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe9_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe9_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe9_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe9_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe9_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe9_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe9_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe9_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe9_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe9_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe9_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe9_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe9_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe9_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe9_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe9_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe9_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe9_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe9_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe9_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe9_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe9_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe9_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe9_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe9_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe9_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe9_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe9_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe9_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe9_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe9_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe9_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe9_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe9_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe9_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe9_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe9_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe9_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe9_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe9_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe9_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe9_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe9_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe9_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe9_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe9_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe9_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe9_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe9_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe9_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe9_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe9_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe9_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe9_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe9_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe9_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe9_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe9_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe9_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe9_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe9_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe9_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe9_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe9_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe9_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe9_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe9_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe9_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe9_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe9_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe9_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe9_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe9_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe9_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe9_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe9_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe9_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe9_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe9_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe9_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe9_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe9_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe9_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe9_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe9_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe9_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe9_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe9_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe9_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe9_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe9_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe9_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe9_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe9_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe9_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe9_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe9_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe9_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe9_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe9_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe9_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe9_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe9_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe9_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe9_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe9_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe9_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe9_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe9_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe9_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe9_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe9_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe9_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe9_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe9_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe9_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe9_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe9_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe9_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe9_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe9_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe9_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe9_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe9_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe9_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe9_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe9_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe9_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe9_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe9_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe9_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe9_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe9_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe9_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe9_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe9_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe9_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe9_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe9_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe9_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe9_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe9_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe9_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe9_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe9_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe9_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe9_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe9_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe9_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe9_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe9_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe9_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe9_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe9_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe9_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe9_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe9_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe9_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe9_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe9_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe9_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe9_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe9_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe9_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe9_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe9_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe9_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe9_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe9_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe9_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe9_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe9_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe9_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe9_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe9_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe9_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe9_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe9_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe9_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe9_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe9_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe9_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe9_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe9_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe9_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe9_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe9_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe9_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe9_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe9_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe9_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe9_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe9_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe9_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe9_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe9_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe9_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe9_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe9_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe9_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe9_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe9_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe9_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe9_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe9_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe9_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe9_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe9_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe9_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe9_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe9_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe9_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe9_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe9_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe9_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe9_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe9_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe9_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe9_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe9_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe9_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe9_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe9_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe9_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe9_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe9_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe9_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe9_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe9_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe9_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe9_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe9_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe9_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe9_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe9_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe9_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe9_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe9_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe9_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe9_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe9_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe9_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe9_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe9_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe9_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe9_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe9_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe9_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe9_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe9_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe9_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe9_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe9_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe9_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe9_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe9_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe9_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe9_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe9_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe9_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe9_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe9_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe9_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe9_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe9_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe9_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe9_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe9_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe9_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe9_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe9_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe9_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe9_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe9_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe9_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe9_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe9_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe9_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe9_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe9_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe9_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe9_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe9_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe9_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe9_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe9_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe9_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe9_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe9_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe9_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe9_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe9_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe9_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe9_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe9_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe9_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe9_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe9_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe9_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe9_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe9_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe9_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe9_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe9_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe9_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe9_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe9_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe9_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe9_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe9_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe9_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe9_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe9_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe9_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe9_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe9_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe9_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe9_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe9_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe9_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe9_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe9_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe9_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe9_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe9_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe9_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe9_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe9_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe9_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe9_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe9_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe9_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe9_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe9_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe9_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe9_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe9_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe9_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe9_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe9_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe9_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe9_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe9_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe9_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe9_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe9_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe9_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe9_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe9_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe9_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe9_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe9_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe9_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe9_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe9_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe9_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe9_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe9_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe9_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe9_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe9_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe9_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe9_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe9_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe9_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe9_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe9_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe9_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe9_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe9_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe9_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe9_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe9_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe9_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe9_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe9_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe9_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe9_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe9_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe9_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe9_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe9_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe9_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe9_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe9_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe9_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe9_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe9_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe9_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe9_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe9_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe9_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe9_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe9_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe9_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe9_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe9_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe9_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe9_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe9_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe9_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe9_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe9_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe9_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe9_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe9_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe9_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe9_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe9_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe9_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe9_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe9_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe9_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe9_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe9_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe9_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe9_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe9_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe9_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe9_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe9_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe9_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe9_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe9_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe9_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe9_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe9_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe9_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe9_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe9_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe9_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe9_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe9_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe9_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe9_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe9_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe9_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe9_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe9_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe9_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe9_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe9_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe9_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe9_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe9_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe9_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe9_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe9_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe9_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe9_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe9_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe9_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe9_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe9_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe9_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe9_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe9_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe9_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe9_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe9_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe9_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe9_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe9_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe9_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe9_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe9_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe9_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe9_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe9_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe9_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe9_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe9_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe9_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe9_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe9_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe9_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe9_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe9_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe9_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe9_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe9_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe9_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe9_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe9_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe9_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe9_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe9_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe9_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe9_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe9_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe9_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe9_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe9_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe9_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe9_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe9_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe9_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe9_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe9_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe9_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe9_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe9_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe9_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe9_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe9_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe9_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe9_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe9_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe9_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe9_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe9_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe9_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe9_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe9_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe9_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe9_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe9_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe9_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe9_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe9_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe9_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe9_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe9_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe9_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe9_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe9_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe9_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe9_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe9_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe9_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe9_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe9_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe9_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe9_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe9_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe9_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe9_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe9_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe9_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe9_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe9_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe9_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe9_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe9_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe9_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe9_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe9_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe9_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe9_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe9_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe9_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe9_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe9_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe9_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe9_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe9_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe9_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe9_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe9_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe9_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe9_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe9_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe9_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe9_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe9_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe9_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe9_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe9_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe9_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe9_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe9_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe9_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe9_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe9_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe9_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe9_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe9_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe9_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe9_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe9_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe9_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe9_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe9_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe9_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe9_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe9_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe9_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe9_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe9_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe9_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe9_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe9_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe9_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe9_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe9_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe9_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe9_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe9_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe9_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe9_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe9_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe9_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe9_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe9_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe9_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe9_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe9_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe9_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe9_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe9_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe9_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe9_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe9_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe9_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe9_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe9_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe9_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe9_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe9_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe9_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe9_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe9_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe9_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe9_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe9_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe9_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe9_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe9_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe9_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe9_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe9_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe9_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe9_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe9_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe9_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe9_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe9_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe9_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe9_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe9_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe9_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe9_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe9_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe9_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe9_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe9_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe9_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe9_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe9_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe9_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe9_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe9_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe9_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe9_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe9_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe9_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe9_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe9_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe9_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe9_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe9_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe9_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe9_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe9_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe9_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe9_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe9_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe9_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe9_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe9_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe9_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe9_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe9_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe9_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe9_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe9_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe9_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe9_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe9_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe9_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe9_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe9_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe9_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe9_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe9_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe9_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe9_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe9_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe9_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe9_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe9_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe9_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe9_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe9_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe9_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe9_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe9_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe9_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe9_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe9_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe9_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe9_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe9_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe9_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe9_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe9_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe9_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe9_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe9_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe9_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe9_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe9_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe9_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe9_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe9_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe9_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe9_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe9_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe9_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe9_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe9_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe9_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe9_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe9_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe9_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe9_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe9_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe9_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe9_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe9_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe9_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe9_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe9_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe9_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe9_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe9_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe9_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe9_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe9_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe9_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe9_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe9_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe9_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe9_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe9_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe9_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe9_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe9_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe9_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe9_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe9_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe9_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe9_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe9_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe9_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe9_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe9_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe9_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe9_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe9_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe9_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe9_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe9_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe9_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe9_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe9_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe9_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe9_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe9_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe9_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe9_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe9_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe9_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe9_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe9_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe9_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe9_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe9_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe9_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe9_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe9_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe9_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe9_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe9_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe9_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe9_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe9_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe9_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe9_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe9_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe9_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe9_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe9_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe9_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe9_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe9_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe9_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe9_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe9_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe9_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe9_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe9_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe9_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe9_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe9_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe9_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe9_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe9_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe9_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe9_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe9_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe9_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe9_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe9_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe9_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe9_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe9_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe9_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe9_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe9_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe9_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe9_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe9_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe9_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe9_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe9_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe9_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe9_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe9_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe9_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe9_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe9_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe9_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe9_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe9_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe9_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe9_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe9_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe9_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe9_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe9_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe9_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe9_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe9_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe9_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe9_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe9_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe9_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe9_io_pipe_phv_out_is_valid_processor),
    .io_table_config_0_table_width(pipe9_io_table_config_0_table_width),
    .io_table_config_0_table_depth(pipe9_io_table_config_0_table_depth),
    .io_table_config_1_table_width(pipe9_io_table_config_1_table_width),
    .io_table_config_1_table_depth(pipe9_io_table_config_1_table_depth),
    .io_key_in(pipe9_io_key_in),
    .io_key_out(pipe9_io_key_out),
    .io_addr_in(pipe9_io_addr_in),
    .io_addr_out(pipe9_io_addr_out),
    .io_cs_in(pipe9_io_cs_in),
    .io_cs_out(pipe9_io_cs_out),
    .io_cs_vec_out_0(pipe9_io_cs_vec_out_0),
    .io_cs_vec_out_1(pipe9_io_cs_vec_out_1),
    .io_cs_vec_out_2(pipe9_io_cs_vec_out_2),
    .io_cs_vec_out_3(pipe9_io_cs_vec_out_3),
    .io_cs_vec_out_4(pipe9_io_cs_vec_out_4),
    .io_cs_vec_out_5(pipe9_io_cs_vec_out_5),
    .io_cs_vec_out_6(pipe9_io_cs_vec_out_6),
    .io_cs_vec_out_7(pipe9_io_cs_vec_out_7),
    .io_cs_vec_out_8(pipe9_io_cs_vec_out_8),
    .io_cs_vec_out_9(pipe9_io_cs_vec_out_9),
    .io_cs_vec_out_10(pipe9_io_cs_vec_out_10),
    .io_cs_vec_out_11(pipe9_io_cs_vec_out_11),
    .io_cs_vec_out_12(pipe9_io_cs_vec_out_12),
    .io_cs_vec_out_13(pipe9_io_cs_vec_out_13),
    .io_cs_vec_out_14(pipe9_io_cs_vec_out_14),
    .io_cs_vec_out_15(pipe9_io_cs_vec_out_15)
  );
  MatchReadData pipe10 ( // @[matcher.scala 347:24]
    .clock(pipe10_clock),
    .io_pipe_phv_in_data_0(pipe10_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe10_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe10_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe10_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe10_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe10_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe10_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe10_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe10_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe10_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe10_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe10_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe10_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe10_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe10_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe10_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe10_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe10_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe10_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe10_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe10_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe10_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe10_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe10_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe10_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe10_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe10_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe10_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe10_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe10_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe10_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe10_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe10_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe10_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe10_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe10_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe10_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe10_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe10_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe10_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe10_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe10_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe10_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe10_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe10_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe10_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe10_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe10_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe10_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe10_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe10_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe10_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe10_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe10_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe10_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe10_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe10_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe10_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe10_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe10_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe10_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe10_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe10_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe10_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe10_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe10_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe10_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe10_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe10_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe10_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe10_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe10_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe10_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe10_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe10_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe10_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe10_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe10_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe10_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe10_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe10_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe10_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe10_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe10_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe10_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe10_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe10_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe10_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe10_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe10_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe10_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe10_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe10_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe10_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe10_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe10_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe10_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe10_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe10_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe10_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe10_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe10_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe10_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe10_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe10_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe10_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe10_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe10_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe10_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe10_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe10_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe10_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe10_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe10_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe10_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe10_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe10_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe10_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe10_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe10_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe10_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe10_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe10_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe10_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe10_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe10_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe10_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe10_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe10_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe10_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe10_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe10_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe10_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe10_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe10_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe10_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe10_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe10_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe10_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe10_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe10_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe10_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe10_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe10_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe10_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe10_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe10_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe10_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe10_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe10_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe10_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe10_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe10_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe10_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe10_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe10_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe10_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe10_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe10_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe10_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe10_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe10_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe10_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe10_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe10_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe10_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe10_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe10_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe10_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe10_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe10_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe10_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe10_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe10_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe10_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe10_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe10_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe10_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe10_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe10_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe10_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe10_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe10_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe10_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe10_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe10_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe10_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe10_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe10_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe10_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe10_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe10_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe10_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe10_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe10_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe10_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe10_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe10_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe10_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe10_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe10_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe10_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe10_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe10_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe10_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe10_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe10_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe10_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe10_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe10_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe10_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe10_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe10_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe10_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe10_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe10_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe10_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe10_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe10_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe10_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe10_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe10_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe10_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe10_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe10_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe10_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe10_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe10_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe10_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe10_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe10_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe10_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe10_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe10_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe10_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe10_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe10_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe10_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe10_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe10_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe10_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe10_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe10_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe10_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe10_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe10_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe10_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe10_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe10_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe10_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe10_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe10_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe10_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe10_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe10_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe10_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe10_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe10_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe10_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe10_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe10_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe10_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe10_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe10_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe10_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe10_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe10_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe10_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe10_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe10_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe10_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe10_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe10_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe10_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe10_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe10_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe10_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe10_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe10_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe10_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe10_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe10_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe10_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe10_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe10_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe10_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe10_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe10_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe10_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe10_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe10_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe10_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe10_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe10_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe10_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe10_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe10_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe10_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe10_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe10_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe10_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe10_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe10_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe10_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe10_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe10_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe10_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe10_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe10_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe10_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe10_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe10_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe10_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe10_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe10_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe10_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe10_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe10_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe10_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe10_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe10_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe10_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe10_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe10_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe10_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe10_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe10_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe10_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe10_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe10_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe10_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe10_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe10_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe10_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe10_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe10_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe10_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe10_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe10_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe10_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe10_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe10_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe10_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe10_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe10_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe10_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe10_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe10_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe10_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe10_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe10_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe10_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe10_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe10_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe10_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe10_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe10_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe10_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe10_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe10_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe10_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe10_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe10_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe10_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe10_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe10_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe10_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe10_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe10_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe10_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe10_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe10_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe10_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe10_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe10_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe10_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe10_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe10_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe10_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe10_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe10_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe10_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe10_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe10_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe10_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe10_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe10_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe10_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe10_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe10_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe10_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe10_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe10_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe10_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe10_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe10_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe10_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe10_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe10_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe10_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe10_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe10_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe10_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe10_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe10_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe10_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe10_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe10_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe10_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe10_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe10_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe10_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe10_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe10_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe10_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe10_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe10_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe10_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe10_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe10_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe10_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe10_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe10_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe10_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe10_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe10_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe10_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe10_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe10_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe10_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe10_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe10_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe10_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe10_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe10_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe10_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe10_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe10_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe10_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe10_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe10_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe10_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe10_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe10_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe10_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe10_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe10_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe10_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe10_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe10_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe10_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe10_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe10_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe10_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe10_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe10_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe10_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe10_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe10_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe10_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe10_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe10_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe10_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe10_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe10_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe10_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe10_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe10_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe10_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe10_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe10_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe10_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe10_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe10_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe10_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe10_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe10_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe10_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe10_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe10_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe10_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe10_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe10_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe10_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe10_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe10_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe10_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe10_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe10_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe10_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe10_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe10_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe10_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe10_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe10_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe10_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe10_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe10_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe10_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe10_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe10_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe10_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe10_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe10_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe10_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe10_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe10_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe10_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe10_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe10_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe10_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe10_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe10_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe10_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe10_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe10_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe10_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe10_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe10_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe10_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe10_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe10_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe10_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe10_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe10_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe10_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe10_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe10_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe10_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe10_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe10_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe10_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe10_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe10_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe10_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe10_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe10_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe10_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe10_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe10_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe10_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe10_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe10_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe10_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe10_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe10_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe10_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe10_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe10_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe10_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe10_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe10_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe10_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe10_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe10_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe10_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe10_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe10_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe10_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe10_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe10_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe10_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe10_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe10_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe10_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe10_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe10_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe10_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe10_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe10_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe10_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe10_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe10_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe10_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe10_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe10_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe10_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe10_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe10_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe10_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe10_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe10_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe10_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe10_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe10_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe10_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe10_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe10_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe10_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe10_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe10_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe10_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe10_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe10_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe10_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe10_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe10_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe10_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe10_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe10_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe10_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe10_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe10_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe10_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe10_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe10_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe10_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe10_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe10_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe10_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe10_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe10_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe10_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe10_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe10_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe10_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe10_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe10_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe10_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe10_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe10_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe10_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe10_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe10_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe10_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe10_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe10_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe10_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe10_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe10_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe10_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe10_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe10_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe10_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe10_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe10_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe10_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe10_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe10_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe10_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe10_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe10_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe10_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe10_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe10_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe10_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe10_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe10_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe10_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe10_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe10_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe10_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe10_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe10_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe10_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe10_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe10_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe10_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe10_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe10_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe10_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe10_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe10_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe10_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe10_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe10_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe10_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe10_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe10_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe10_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe10_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe10_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe10_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe10_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe10_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe10_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe10_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe10_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe10_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe10_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe10_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe10_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe10_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe10_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe10_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe10_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe10_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe10_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe10_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe10_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe10_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe10_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe10_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe10_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe10_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe10_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe10_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe10_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe10_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe10_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe10_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe10_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe10_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe10_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe10_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe10_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe10_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe10_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe10_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe10_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe10_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe10_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe10_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe10_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe10_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe10_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe10_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe10_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe10_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe10_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe10_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe10_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe10_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe10_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe10_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe10_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe10_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe10_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe10_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe10_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe10_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe10_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe10_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe10_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe10_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe10_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe10_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe10_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe10_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe10_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe10_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe10_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe10_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe10_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe10_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe10_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe10_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe10_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe10_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe10_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe10_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe10_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe10_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe10_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe10_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe10_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe10_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe10_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe10_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe10_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe10_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe10_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe10_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe10_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe10_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe10_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe10_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe10_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe10_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe10_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe10_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe10_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe10_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe10_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe10_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe10_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe10_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe10_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe10_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe10_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe10_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe10_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe10_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe10_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe10_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe10_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe10_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe10_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe10_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe10_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe10_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe10_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe10_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe10_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe10_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe10_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe10_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe10_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe10_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe10_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe10_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe10_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe10_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe10_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe10_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe10_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe10_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe10_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe10_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe10_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe10_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe10_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe10_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe10_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe10_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe10_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe10_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe10_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe10_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe10_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe10_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe10_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe10_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe10_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe10_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe10_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe10_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe10_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe10_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe10_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe10_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe10_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe10_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe10_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe10_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe10_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe10_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe10_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe10_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe10_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe10_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe10_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe10_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe10_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe10_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe10_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe10_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe10_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe10_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe10_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe10_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe10_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe10_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe10_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe10_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe10_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe10_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe10_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe10_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe10_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe10_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe10_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe10_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe10_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe10_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe10_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe10_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe10_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe10_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe10_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe10_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe10_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe10_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe10_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe10_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe10_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe10_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe10_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe10_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe10_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe10_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe10_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe10_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe10_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe10_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe10_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe10_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe10_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe10_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe10_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe10_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe10_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe10_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe10_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe10_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe10_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe10_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe10_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe10_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe10_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe10_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe10_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe10_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe10_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe10_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe10_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe10_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe10_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe10_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe10_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe10_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe10_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe10_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe10_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe10_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe10_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe10_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe10_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe10_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe10_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe10_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe10_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe10_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe10_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe10_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe10_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe10_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe10_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe10_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe10_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe10_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe10_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe10_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe10_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe10_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe10_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe10_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe10_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe10_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe10_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe10_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe10_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe10_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe10_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe10_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe10_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe10_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe10_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe10_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe10_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe10_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe10_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe10_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe10_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe10_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe10_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe10_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe10_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe10_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe10_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe10_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe10_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe10_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe10_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe10_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe10_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe10_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe10_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe10_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe10_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe10_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe10_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe10_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe10_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe10_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe10_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe10_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe10_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe10_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe10_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe10_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe10_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe10_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe10_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe10_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe10_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe10_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe10_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe10_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe10_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe10_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe10_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe10_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe10_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe10_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe10_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe10_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe10_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe10_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe10_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe10_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe10_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe10_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe10_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe10_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe10_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe10_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe10_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe10_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe10_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe10_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe10_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe10_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe10_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe10_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe10_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe10_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe10_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe10_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe10_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe10_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe10_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe10_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe10_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe10_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe10_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe10_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe10_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe10_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe10_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe10_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe10_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe10_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe10_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe10_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe10_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe10_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe10_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe10_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe10_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe10_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe10_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe10_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe10_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe10_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe10_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe10_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe10_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe10_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe10_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe10_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe10_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe10_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe10_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe10_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe10_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe10_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe10_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe10_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe10_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe10_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe10_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe10_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe10_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe10_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe10_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe10_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe10_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe10_io_key_in),
    .io_key_out(pipe10_io_key_out),
    .io_cs_in(pipe10_io_cs_in),
    .io_cs_out(pipe10_io_cs_out),
    .io_addr_in(pipe10_io_addr_in),
    .io_cs_vec_in_0(pipe10_io_cs_vec_in_0),
    .io_cs_vec_in_1(pipe10_io_cs_vec_in_1),
    .io_cs_vec_in_2(pipe10_io_cs_vec_in_2),
    .io_cs_vec_in_3(pipe10_io_cs_vec_in_3),
    .io_cs_vec_in_4(pipe10_io_cs_vec_in_4),
    .io_cs_vec_in_5(pipe10_io_cs_vec_in_5),
    .io_cs_vec_in_6(pipe10_io_cs_vec_in_6),
    .io_cs_vec_in_7(pipe10_io_cs_vec_in_7),
    .io_cs_vec_in_8(pipe10_io_cs_vec_in_8),
    .io_cs_vec_in_9(pipe10_io_cs_vec_in_9),
    .io_cs_vec_in_10(pipe10_io_cs_vec_in_10),
    .io_cs_vec_in_11(pipe10_io_cs_vec_in_11),
    .io_cs_vec_in_12(pipe10_io_cs_vec_in_12),
    .io_cs_vec_in_13(pipe10_io_cs_vec_in_13),
    .io_cs_vec_in_14(pipe10_io_cs_vec_in_14),
    .io_cs_vec_in_15(pipe10_io_cs_vec_in_15),
    .io_data_out_0(pipe10_io_data_out_0),
    .io_data_out_1(pipe10_io_data_out_1),
    .io_data_out_2(pipe10_io_data_out_2),
    .io_data_out_3(pipe10_io_data_out_3),
    .io_data_out_4(pipe10_io_data_out_4),
    .io_data_out_5(pipe10_io_data_out_5),
    .io_data_out_6(pipe10_io_data_out_6),
    .io_data_out_7(pipe10_io_data_out_7),
    .io_data_out_8(pipe10_io_data_out_8),
    .io_data_out_9(pipe10_io_data_out_9),
    .io_data_out_10(pipe10_io_data_out_10),
    .io_data_out_11(pipe10_io_data_out_11),
    .io_data_out_12(pipe10_io_data_out_12),
    .io_data_out_13(pipe10_io_data_out_13),
    .io_data_out_14(pipe10_io_data_out_14),
    .io_data_out_15(pipe10_io_data_out_15),
    .io_mem_cluster_0_en(pipe10_io_mem_cluster_0_en),
    .io_mem_cluster_0_addr(pipe10_io_mem_cluster_0_addr),
    .io_mem_cluster_0_data(pipe10_io_mem_cluster_0_data),
    .io_mem_cluster_1_en(pipe10_io_mem_cluster_1_en),
    .io_mem_cluster_1_addr(pipe10_io_mem_cluster_1_addr),
    .io_mem_cluster_1_data(pipe10_io_mem_cluster_1_data),
    .io_mem_cluster_2_en(pipe10_io_mem_cluster_2_en),
    .io_mem_cluster_2_addr(pipe10_io_mem_cluster_2_addr),
    .io_mem_cluster_2_data(pipe10_io_mem_cluster_2_data),
    .io_mem_cluster_3_en(pipe10_io_mem_cluster_3_en),
    .io_mem_cluster_3_addr(pipe10_io_mem_cluster_3_addr),
    .io_mem_cluster_3_data(pipe10_io_mem_cluster_3_data),
    .io_mem_cluster_4_en(pipe10_io_mem_cluster_4_en),
    .io_mem_cluster_4_addr(pipe10_io_mem_cluster_4_addr),
    .io_mem_cluster_4_data(pipe10_io_mem_cluster_4_data),
    .io_mem_cluster_5_en(pipe10_io_mem_cluster_5_en),
    .io_mem_cluster_5_addr(pipe10_io_mem_cluster_5_addr),
    .io_mem_cluster_5_data(pipe10_io_mem_cluster_5_data),
    .io_mem_cluster_6_en(pipe10_io_mem_cluster_6_en),
    .io_mem_cluster_6_addr(pipe10_io_mem_cluster_6_addr),
    .io_mem_cluster_6_data(pipe10_io_mem_cluster_6_data),
    .io_mem_cluster_7_en(pipe10_io_mem_cluster_7_en),
    .io_mem_cluster_7_addr(pipe10_io_mem_cluster_7_addr),
    .io_mem_cluster_7_data(pipe10_io_mem_cluster_7_data),
    .io_mem_cluster_8_en(pipe10_io_mem_cluster_8_en),
    .io_mem_cluster_8_addr(pipe10_io_mem_cluster_8_addr),
    .io_mem_cluster_8_data(pipe10_io_mem_cluster_8_data),
    .io_mem_cluster_9_en(pipe10_io_mem_cluster_9_en),
    .io_mem_cluster_9_addr(pipe10_io_mem_cluster_9_addr),
    .io_mem_cluster_9_data(pipe10_io_mem_cluster_9_data),
    .io_mem_cluster_10_en(pipe10_io_mem_cluster_10_en),
    .io_mem_cluster_10_addr(pipe10_io_mem_cluster_10_addr),
    .io_mem_cluster_10_data(pipe10_io_mem_cluster_10_data),
    .io_mem_cluster_11_en(pipe10_io_mem_cluster_11_en),
    .io_mem_cluster_11_addr(pipe10_io_mem_cluster_11_addr),
    .io_mem_cluster_11_data(pipe10_io_mem_cluster_11_data),
    .io_mem_cluster_12_en(pipe10_io_mem_cluster_12_en),
    .io_mem_cluster_12_addr(pipe10_io_mem_cluster_12_addr),
    .io_mem_cluster_12_data(pipe10_io_mem_cluster_12_data),
    .io_mem_cluster_13_en(pipe10_io_mem_cluster_13_en),
    .io_mem_cluster_13_addr(pipe10_io_mem_cluster_13_addr),
    .io_mem_cluster_13_data(pipe10_io_mem_cluster_13_data),
    .io_mem_cluster_14_en(pipe10_io_mem_cluster_14_en),
    .io_mem_cluster_14_addr(pipe10_io_mem_cluster_14_addr),
    .io_mem_cluster_14_data(pipe10_io_mem_cluster_14_data),
    .io_mem_cluster_15_en(pipe10_io_mem_cluster_15_en),
    .io_mem_cluster_15_addr(pipe10_io_mem_cluster_15_addr),
    .io_mem_cluster_15_data(pipe10_io_mem_cluster_15_data)
  );
  MatchDataReshape pipe11 ( // @[matcher.scala 348:24]
    .clock(pipe11_clock),
    .io_pipe_phv_in_data_0(pipe11_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe11_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe11_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe11_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe11_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe11_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe11_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe11_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe11_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe11_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe11_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe11_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe11_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe11_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe11_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe11_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe11_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe11_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe11_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe11_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe11_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe11_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe11_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe11_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe11_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe11_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe11_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe11_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe11_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe11_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe11_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe11_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe11_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe11_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe11_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe11_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe11_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe11_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe11_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe11_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe11_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe11_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe11_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe11_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe11_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe11_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe11_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe11_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe11_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe11_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe11_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe11_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe11_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe11_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe11_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe11_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe11_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe11_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe11_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe11_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe11_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe11_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe11_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe11_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe11_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe11_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe11_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe11_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe11_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe11_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe11_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe11_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe11_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe11_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe11_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe11_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe11_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe11_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe11_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe11_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe11_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe11_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe11_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe11_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe11_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe11_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe11_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe11_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe11_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe11_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe11_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe11_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe11_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe11_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe11_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe11_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe11_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe11_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe11_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe11_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe11_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe11_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe11_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe11_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe11_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe11_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe11_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe11_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe11_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe11_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe11_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe11_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe11_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe11_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe11_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe11_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe11_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe11_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe11_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe11_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe11_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe11_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe11_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe11_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe11_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe11_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe11_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe11_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe11_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe11_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe11_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe11_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe11_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe11_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe11_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe11_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe11_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe11_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe11_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe11_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe11_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe11_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe11_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe11_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe11_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe11_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe11_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe11_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe11_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe11_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe11_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe11_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe11_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe11_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe11_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe11_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe11_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe11_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe11_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe11_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe11_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe11_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe11_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe11_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe11_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe11_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe11_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe11_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe11_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe11_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe11_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe11_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe11_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe11_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe11_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe11_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe11_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe11_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe11_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe11_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe11_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe11_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe11_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe11_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe11_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe11_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe11_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe11_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe11_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe11_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe11_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe11_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe11_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe11_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe11_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe11_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe11_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe11_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe11_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe11_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe11_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe11_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe11_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe11_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe11_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe11_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe11_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe11_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe11_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe11_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe11_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe11_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe11_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe11_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe11_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe11_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe11_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe11_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe11_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe11_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe11_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe11_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe11_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe11_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe11_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe11_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe11_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe11_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe11_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe11_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe11_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe11_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe11_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe11_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe11_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe11_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe11_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe11_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe11_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe11_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe11_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe11_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe11_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe11_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe11_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe11_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe11_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe11_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe11_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe11_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe11_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe11_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe11_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe11_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe11_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe11_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe11_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe11_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe11_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe11_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe11_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe11_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe11_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe11_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe11_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe11_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe11_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe11_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe11_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe11_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe11_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe11_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe11_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe11_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe11_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe11_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe11_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe11_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe11_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe11_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe11_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe11_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe11_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe11_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe11_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe11_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe11_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe11_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe11_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe11_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe11_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe11_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe11_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe11_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe11_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe11_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe11_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe11_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe11_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe11_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe11_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe11_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe11_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe11_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe11_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe11_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe11_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe11_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe11_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe11_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe11_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe11_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe11_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe11_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe11_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe11_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe11_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe11_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe11_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe11_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe11_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe11_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe11_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe11_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe11_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe11_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe11_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe11_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe11_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe11_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe11_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe11_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe11_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe11_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe11_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe11_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe11_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe11_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe11_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe11_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe11_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe11_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe11_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe11_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe11_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe11_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe11_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe11_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe11_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe11_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe11_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe11_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe11_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe11_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe11_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe11_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe11_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe11_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe11_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe11_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe11_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe11_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe11_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe11_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe11_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe11_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe11_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe11_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe11_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe11_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe11_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe11_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe11_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe11_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe11_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe11_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe11_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe11_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe11_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe11_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe11_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe11_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe11_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe11_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe11_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe11_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe11_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe11_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe11_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe11_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe11_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe11_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe11_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe11_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe11_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe11_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe11_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe11_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe11_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe11_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe11_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe11_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe11_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe11_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe11_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe11_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe11_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe11_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe11_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe11_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe11_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe11_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe11_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe11_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe11_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe11_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe11_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe11_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe11_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe11_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe11_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe11_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe11_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe11_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe11_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe11_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe11_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe11_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe11_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe11_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe11_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe11_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe11_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe11_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe11_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe11_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe11_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe11_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe11_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe11_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe11_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe11_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe11_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe11_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe11_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe11_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe11_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe11_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe11_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe11_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe11_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe11_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe11_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe11_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe11_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe11_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe11_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe11_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe11_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe11_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe11_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe11_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe11_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe11_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe11_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe11_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe11_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe11_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe11_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe11_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe11_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe11_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe11_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe11_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe11_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe11_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe11_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe11_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe11_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe11_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe11_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe11_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe11_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe11_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe11_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe11_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe11_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe11_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe11_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe11_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe11_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe11_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe11_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe11_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe11_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe11_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe11_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe11_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe11_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe11_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe11_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe11_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe11_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe11_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe11_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe11_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe11_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe11_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe11_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe11_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe11_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe11_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe11_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe11_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe11_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe11_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe11_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe11_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe11_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe11_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe11_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe11_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe11_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe11_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe11_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe11_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe11_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe11_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe11_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe11_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe11_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe11_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe11_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe11_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe11_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe11_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe11_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe11_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe11_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe11_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe11_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe11_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe11_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe11_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe11_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe11_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe11_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe11_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe11_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe11_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe11_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe11_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe11_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe11_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe11_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe11_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe11_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe11_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe11_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe11_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe11_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe11_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe11_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe11_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe11_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe11_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe11_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe11_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe11_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe11_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe11_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe11_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe11_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe11_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe11_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe11_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe11_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe11_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe11_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe11_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe11_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe11_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe11_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe11_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe11_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe11_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe11_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe11_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe11_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe11_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe11_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe11_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe11_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe11_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe11_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe11_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe11_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe11_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe11_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe11_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe11_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe11_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe11_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe11_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe11_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe11_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe11_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe11_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe11_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe11_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe11_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe11_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe11_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe11_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe11_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe11_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe11_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe11_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe11_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe11_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe11_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe11_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe11_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe11_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe11_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe11_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe11_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe11_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe11_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe11_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe11_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe11_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe11_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe11_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe11_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe11_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe11_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe11_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe11_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe11_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe11_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe11_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe11_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe11_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe11_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe11_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe11_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe11_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe11_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe11_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe11_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe11_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe11_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe11_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe11_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe11_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe11_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe11_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe11_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe11_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe11_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe11_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe11_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe11_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe11_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe11_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe11_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe11_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe11_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe11_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe11_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe11_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe11_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe11_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe11_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe11_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe11_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe11_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe11_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe11_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe11_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe11_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe11_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe11_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe11_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe11_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe11_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe11_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe11_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe11_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe11_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe11_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe11_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe11_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe11_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe11_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe11_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe11_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe11_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe11_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe11_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe11_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe11_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe11_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe11_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe11_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe11_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe11_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe11_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe11_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe11_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe11_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe11_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe11_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe11_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe11_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe11_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe11_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe11_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe11_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe11_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe11_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe11_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe11_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe11_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe11_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe11_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe11_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe11_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe11_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe11_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe11_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe11_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe11_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe11_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe11_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe11_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe11_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe11_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe11_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe11_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe11_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe11_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe11_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe11_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe11_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe11_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe11_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe11_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe11_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe11_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe11_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe11_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe11_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe11_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe11_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe11_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe11_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe11_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe11_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe11_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe11_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe11_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe11_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe11_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe11_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe11_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe11_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe11_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe11_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe11_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe11_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe11_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe11_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe11_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe11_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe11_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe11_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe11_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe11_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe11_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe11_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe11_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe11_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe11_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe11_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe11_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe11_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe11_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe11_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe11_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe11_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe11_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe11_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe11_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe11_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe11_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe11_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe11_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe11_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe11_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe11_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe11_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe11_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe11_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe11_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe11_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe11_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe11_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe11_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe11_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe11_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe11_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe11_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe11_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe11_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe11_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe11_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe11_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe11_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe11_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe11_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe11_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe11_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe11_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe11_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe11_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe11_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe11_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe11_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe11_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe11_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe11_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe11_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe11_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe11_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe11_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe11_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe11_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe11_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe11_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe11_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe11_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe11_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe11_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe11_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe11_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe11_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe11_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe11_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe11_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe11_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe11_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe11_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe11_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe11_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe11_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe11_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe11_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe11_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe11_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe11_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe11_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe11_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe11_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe11_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe11_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe11_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe11_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe11_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe11_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe11_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe11_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe11_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe11_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe11_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe11_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe11_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe11_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe11_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe11_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe11_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe11_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe11_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe11_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe11_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe11_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe11_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe11_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe11_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe11_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe11_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe11_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe11_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe11_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe11_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe11_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe11_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe11_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe11_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe11_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe11_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe11_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe11_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe11_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe11_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe11_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe11_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe11_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe11_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe11_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe11_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe11_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe11_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe11_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe11_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe11_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe11_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe11_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe11_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe11_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe11_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe11_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe11_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe11_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe11_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe11_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe11_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe11_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe11_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe11_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe11_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe11_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe11_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe11_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe11_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe11_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe11_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe11_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe11_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe11_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe11_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe11_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe11_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe11_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe11_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe11_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe11_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe11_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe11_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe11_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe11_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe11_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe11_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe11_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe11_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe11_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe11_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe11_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe11_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe11_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe11_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe11_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe11_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe11_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe11_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe11_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe11_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe11_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe11_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe11_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe11_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe11_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe11_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe11_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe11_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe11_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe11_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe11_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe11_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe11_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe11_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe11_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe11_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe11_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe11_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe11_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe11_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe11_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe11_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe11_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe11_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe11_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe11_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe11_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe11_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe11_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe11_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe11_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe11_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe11_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe11_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe11_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe11_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe11_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe11_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe11_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe11_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe11_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe11_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe11_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe11_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe11_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe11_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe11_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe11_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe11_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe11_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe11_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe11_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe11_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe11_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe11_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe11_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe11_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe11_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe11_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe11_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe11_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe11_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe11_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe11_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe11_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe11_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe11_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe11_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe11_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe11_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe11_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe11_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe11_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe11_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe11_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe11_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe11_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe11_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe11_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe11_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe11_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe11_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe11_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe11_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe11_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe11_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe11_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe11_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe11_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe11_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe11_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe11_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe11_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe11_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe11_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe11_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe11_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe11_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe11_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe11_io_pipe_phv_out_is_valid_processor),
    .io_table_config_0_table_width(pipe11_io_table_config_0_table_width),
    .io_table_config_0_table_depth(pipe11_io_table_config_0_table_depth),
    .io_table_config_1_table_width(pipe11_io_table_config_1_table_width),
    .io_table_config_1_table_depth(pipe11_io_table_config_1_table_depth),
    .io_key_in(pipe11_io_key_in),
    .io_key_out(pipe11_io_key_out),
    .io_cs_in(pipe11_io_cs_in),
    .io_data_in_0(pipe11_io_data_in_0),
    .io_data_in_1(pipe11_io_data_in_1),
    .io_data_in_2(pipe11_io_data_in_2),
    .io_data_in_3(pipe11_io_data_in_3),
    .io_data_in_4(pipe11_io_data_in_4),
    .io_data_in_5(pipe11_io_data_in_5),
    .io_data_in_6(pipe11_io_data_in_6),
    .io_data_in_7(pipe11_io_data_in_7),
    .io_data_in_8(pipe11_io_data_in_8),
    .io_data_in_9(pipe11_io_data_in_9),
    .io_data_in_10(pipe11_io_data_in_10),
    .io_data_in_11(pipe11_io_data_in_11),
    .io_data_in_12(pipe11_io_data_in_12),
    .io_data_in_13(pipe11_io_data_in_13),
    .io_data_in_14(pipe11_io_data_in_14),
    .io_data_in_15(pipe11_io_data_in_15),
    .io_data_out(pipe11_io_data_out)
  );
  MatchResult pipe12 ( // @[matcher.scala 349:24]
    .clock(pipe12_clock),
    .io_pipe_phv_in_data_0(pipe12_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe12_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe12_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe12_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe12_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe12_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe12_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe12_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe12_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe12_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe12_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe12_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe12_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe12_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe12_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe12_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe12_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe12_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe12_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe12_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe12_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe12_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe12_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe12_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe12_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe12_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe12_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe12_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe12_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe12_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe12_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe12_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe12_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe12_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe12_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe12_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe12_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe12_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe12_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe12_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe12_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe12_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe12_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe12_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe12_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe12_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe12_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe12_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe12_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe12_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe12_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe12_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe12_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe12_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe12_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe12_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe12_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe12_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe12_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe12_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe12_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe12_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe12_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe12_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe12_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe12_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe12_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe12_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe12_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe12_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe12_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe12_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe12_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe12_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe12_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe12_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe12_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe12_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe12_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe12_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe12_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe12_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe12_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe12_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe12_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe12_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe12_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe12_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe12_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe12_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe12_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe12_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe12_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe12_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe12_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe12_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe12_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe12_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe12_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe12_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe12_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe12_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe12_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe12_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe12_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe12_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe12_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe12_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe12_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe12_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe12_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe12_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe12_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe12_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe12_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe12_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe12_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe12_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe12_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe12_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe12_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe12_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe12_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe12_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe12_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe12_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe12_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe12_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe12_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe12_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe12_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe12_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe12_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe12_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe12_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe12_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe12_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe12_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe12_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe12_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe12_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe12_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe12_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe12_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe12_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe12_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe12_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe12_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe12_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe12_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe12_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe12_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe12_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe12_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe12_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe12_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe12_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe12_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe12_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe12_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe12_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe12_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe12_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe12_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe12_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe12_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe12_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe12_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe12_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe12_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe12_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe12_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe12_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe12_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe12_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe12_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe12_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe12_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe12_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe12_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe12_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe12_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe12_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe12_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe12_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe12_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe12_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe12_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe12_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe12_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe12_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe12_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe12_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe12_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe12_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe12_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe12_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe12_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe12_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe12_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe12_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe12_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe12_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe12_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe12_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe12_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe12_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe12_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe12_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe12_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe12_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe12_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe12_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe12_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe12_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe12_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe12_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe12_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe12_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe12_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe12_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe12_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe12_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe12_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe12_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe12_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe12_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe12_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe12_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe12_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe12_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe12_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe12_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe12_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe12_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe12_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe12_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe12_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe12_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe12_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe12_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe12_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe12_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe12_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe12_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe12_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe12_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe12_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe12_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe12_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe12_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe12_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe12_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe12_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe12_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe12_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe12_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe12_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe12_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe12_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe12_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe12_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe12_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe12_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe12_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe12_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe12_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe12_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe12_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe12_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe12_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe12_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe12_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe12_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe12_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe12_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe12_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe12_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe12_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe12_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe12_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe12_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe12_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe12_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe12_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe12_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe12_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe12_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe12_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe12_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe12_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe12_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe12_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe12_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe12_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe12_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe12_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe12_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe12_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe12_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe12_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe12_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe12_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe12_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe12_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe12_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe12_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe12_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe12_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe12_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe12_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe12_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe12_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe12_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe12_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe12_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe12_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe12_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe12_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe12_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe12_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe12_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe12_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe12_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe12_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe12_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe12_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe12_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe12_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe12_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe12_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe12_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe12_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe12_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe12_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe12_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe12_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe12_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe12_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe12_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe12_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe12_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe12_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe12_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe12_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe12_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe12_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe12_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe12_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe12_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe12_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe12_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe12_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe12_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe12_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe12_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe12_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe12_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe12_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe12_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe12_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe12_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe12_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe12_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe12_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe12_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe12_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe12_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe12_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe12_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe12_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe12_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe12_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe12_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe12_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe12_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe12_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe12_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe12_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe12_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe12_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe12_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe12_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe12_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe12_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe12_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe12_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe12_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe12_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe12_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe12_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe12_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe12_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe12_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe12_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe12_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe12_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe12_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe12_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe12_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe12_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe12_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe12_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe12_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe12_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe12_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe12_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe12_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe12_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe12_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe12_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe12_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe12_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe12_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe12_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe12_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe12_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe12_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe12_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe12_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe12_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe12_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe12_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe12_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe12_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe12_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe12_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe12_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe12_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe12_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe12_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe12_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe12_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe12_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe12_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe12_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe12_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe12_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe12_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe12_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe12_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe12_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe12_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe12_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe12_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe12_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe12_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe12_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe12_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe12_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe12_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe12_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe12_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe12_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe12_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe12_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe12_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe12_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe12_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe12_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe12_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe12_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe12_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe12_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe12_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe12_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe12_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe12_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe12_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe12_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe12_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe12_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe12_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe12_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe12_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe12_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe12_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe12_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe12_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe12_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe12_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe12_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe12_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe12_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe12_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe12_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe12_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe12_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe12_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe12_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe12_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe12_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe12_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe12_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe12_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe12_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe12_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe12_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe12_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe12_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe12_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe12_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe12_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe12_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe12_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe12_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe12_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe12_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe12_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe12_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe12_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe12_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe12_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe12_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe12_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe12_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe12_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe12_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe12_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe12_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe12_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe12_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe12_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe12_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe12_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe12_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe12_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe12_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe12_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe12_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe12_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe12_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe12_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe12_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe12_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe12_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe12_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe12_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe12_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe12_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe12_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe12_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe12_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe12_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe12_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe12_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe12_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe12_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe12_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe12_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe12_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe12_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe12_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe12_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe12_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe12_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe12_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe12_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe12_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe12_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe12_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe12_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe12_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe12_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe12_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe12_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe12_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe12_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe12_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe12_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe12_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe12_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe12_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe12_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe12_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe12_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe12_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe12_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe12_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe12_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe12_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe12_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe12_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe12_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe12_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe12_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe12_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe12_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe12_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe12_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe12_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe12_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe12_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe12_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe12_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe12_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe12_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe12_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe12_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe12_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe12_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe12_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe12_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe12_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe12_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe12_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe12_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe12_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe12_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe12_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe12_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe12_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe12_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe12_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe12_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe12_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe12_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe12_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe12_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe12_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe12_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe12_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe12_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe12_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe12_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe12_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe12_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe12_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe12_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe12_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe12_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe12_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe12_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe12_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe12_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe12_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe12_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe12_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe12_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe12_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe12_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe12_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe12_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe12_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe12_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe12_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe12_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe12_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe12_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe12_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe12_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe12_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe12_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe12_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe12_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe12_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe12_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe12_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe12_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe12_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe12_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe12_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe12_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe12_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe12_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe12_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe12_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe12_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe12_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe12_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe12_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe12_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe12_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe12_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe12_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe12_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe12_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe12_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe12_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe12_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe12_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe12_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe12_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe12_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe12_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe12_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe12_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe12_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe12_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe12_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe12_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe12_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe12_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe12_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe12_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe12_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe12_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe12_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe12_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe12_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe12_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe12_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe12_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe12_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe12_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe12_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe12_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe12_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe12_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe12_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe12_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe12_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe12_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe12_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe12_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe12_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe12_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe12_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe12_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe12_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe12_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe12_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe12_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe12_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe12_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe12_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe12_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe12_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe12_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe12_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe12_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe12_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe12_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe12_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe12_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe12_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe12_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe12_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe12_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe12_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe12_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe12_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe12_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe12_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe12_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe12_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe12_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe12_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe12_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe12_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe12_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe12_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe12_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe12_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe12_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe12_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe12_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe12_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe12_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe12_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe12_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe12_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe12_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe12_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe12_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe12_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe12_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe12_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe12_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe12_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe12_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe12_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe12_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe12_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe12_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe12_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe12_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe12_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe12_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe12_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe12_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe12_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe12_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe12_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe12_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe12_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe12_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe12_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe12_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe12_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe12_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe12_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe12_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe12_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe12_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe12_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe12_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe12_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe12_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe12_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe12_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe12_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe12_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe12_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe12_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe12_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe12_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe12_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe12_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe12_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe12_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe12_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe12_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe12_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe12_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe12_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe12_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe12_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe12_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe12_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe12_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe12_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe12_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe12_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe12_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe12_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe12_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe12_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe12_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe12_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe12_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe12_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe12_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe12_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe12_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe12_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe12_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe12_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe12_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe12_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe12_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe12_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe12_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe12_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe12_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe12_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe12_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe12_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe12_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe12_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe12_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe12_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe12_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe12_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe12_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe12_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe12_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe12_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe12_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe12_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe12_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe12_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe12_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe12_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe12_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe12_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe12_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe12_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe12_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe12_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe12_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe12_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe12_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe12_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe12_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe12_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe12_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe12_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe12_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe12_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe12_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe12_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe12_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe12_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe12_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe12_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe12_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe12_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe12_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe12_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe12_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe12_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe12_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe12_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe12_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe12_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe12_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe12_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe12_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe12_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe12_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe12_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe12_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe12_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe12_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe12_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe12_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe12_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe12_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe12_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe12_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe12_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe12_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe12_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe12_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe12_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe12_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe12_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe12_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe12_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe12_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe12_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe12_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe12_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe12_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe12_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe12_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe12_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe12_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe12_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe12_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe12_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe12_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe12_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe12_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe12_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe12_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe12_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe12_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe12_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe12_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe12_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe12_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe12_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe12_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe12_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe12_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe12_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe12_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe12_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe12_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe12_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe12_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe12_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe12_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe12_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe12_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe12_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe12_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe12_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe12_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe12_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe12_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe12_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe12_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe12_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe12_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe12_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe12_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe12_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe12_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe12_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe12_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe12_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe12_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe12_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe12_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe12_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe12_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe12_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe12_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe12_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe12_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe12_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe12_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe12_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe12_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe12_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe12_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe12_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe12_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe12_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe12_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe12_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe12_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe12_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe12_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe12_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe12_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe12_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe12_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe12_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe12_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe12_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe12_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe12_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe12_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe12_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe12_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe12_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe12_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe12_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe12_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe12_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe12_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe12_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe12_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe12_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe12_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe12_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe12_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe12_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe12_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe12_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe12_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe12_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe12_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe12_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe12_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe12_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe12_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe12_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe12_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe12_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe12_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe12_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe12_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe12_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe12_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe12_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe12_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe12_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe12_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe12_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe12_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe12_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe12_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe12_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe12_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe12_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe12_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe12_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe12_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe12_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe12_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe12_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe12_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe12_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe12_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe12_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe12_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe12_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe12_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe12_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe12_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe12_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe12_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe12_io_pipe_phv_out_is_valid_processor),
    .io_key_config_0_key_length(pipe12_io_key_config_0_key_length),
    .io_key_config_1_key_length(pipe12_io_key_config_1_key_length),
    .io_key_in(pipe12_io_key_in),
    .io_data_in(pipe12_io_data_in),
    .io_hit(pipe12_io_hit),
    .io_match_value(pipe12_io_match_value)
  );
  assign io_pipe_phv_out_data_0 = pipe12_io_pipe_phv_out_data_0; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_1 = pipe12_io_pipe_phv_out_data_1; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_2 = pipe12_io_pipe_phv_out_data_2; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_3 = pipe12_io_pipe_phv_out_data_3; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_4 = pipe12_io_pipe_phv_out_data_4; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_5 = pipe12_io_pipe_phv_out_data_5; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_6 = pipe12_io_pipe_phv_out_data_6; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_7 = pipe12_io_pipe_phv_out_data_7; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_8 = pipe12_io_pipe_phv_out_data_8; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_9 = pipe12_io_pipe_phv_out_data_9; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_10 = pipe12_io_pipe_phv_out_data_10; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_11 = pipe12_io_pipe_phv_out_data_11; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_12 = pipe12_io_pipe_phv_out_data_12; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_13 = pipe12_io_pipe_phv_out_data_13; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_14 = pipe12_io_pipe_phv_out_data_14; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_15 = pipe12_io_pipe_phv_out_data_15; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_16 = pipe12_io_pipe_phv_out_data_16; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_17 = pipe12_io_pipe_phv_out_data_17; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_18 = pipe12_io_pipe_phv_out_data_18; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_19 = pipe12_io_pipe_phv_out_data_19; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_20 = pipe12_io_pipe_phv_out_data_20; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_21 = pipe12_io_pipe_phv_out_data_21; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_22 = pipe12_io_pipe_phv_out_data_22; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_23 = pipe12_io_pipe_phv_out_data_23; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_24 = pipe12_io_pipe_phv_out_data_24; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_25 = pipe12_io_pipe_phv_out_data_25; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_26 = pipe12_io_pipe_phv_out_data_26; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_27 = pipe12_io_pipe_phv_out_data_27; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_28 = pipe12_io_pipe_phv_out_data_28; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_29 = pipe12_io_pipe_phv_out_data_29; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_30 = pipe12_io_pipe_phv_out_data_30; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_31 = pipe12_io_pipe_phv_out_data_31; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_32 = pipe12_io_pipe_phv_out_data_32; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_33 = pipe12_io_pipe_phv_out_data_33; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_34 = pipe12_io_pipe_phv_out_data_34; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_35 = pipe12_io_pipe_phv_out_data_35; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_36 = pipe12_io_pipe_phv_out_data_36; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_37 = pipe12_io_pipe_phv_out_data_37; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_38 = pipe12_io_pipe_phv_out_data_38; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_39 = pipe12_io_pipe_phv_out_data_39; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_40 = pipe12_io_pipe_phv_out_data_40; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_41 = pipe12_io_pipe_phv_out_data_41; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_42 = pipe12_io_pipe_phv_out_data_42; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_43 = pipe12_io_pipe_phv_out_data_43; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_44 = pipe12_io_pipe_phv_out_data_44; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_45 = pipe12_io_pipe_phv_out_data_45; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_46 = pipe12_io_pipe_phv_out_data_46; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_47 = pipe12_io_pipe_phv_out_data_47; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_48 = pipe12_io_pipe_phv_out_data_48; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_49 = pipe12_io_pipe_phv_out_data_49; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_50 = pipe12_io_pipe_phv_out_data_50; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_51 = pipe12_io_pipe_phv_out_data_51; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_52 = pipe12_io_pipe_phv_out_data_52; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_53 = pipe12_io_pipe_phv_out_data_53; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_54 = pipe12_io_pipe_phv_out_data_54; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_55 = pipe12_io_pipe_phv_out_data_55; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_56 = pipe12_io_pipe_phv_out_data_56; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_57 = pipe12_io_pipe_phv_out_data_57; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_58 = pipe12_io_pipe_phv_out_data_58; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_59 = pipe12_io_pipe_phv_out_data_59; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_60 = pipe12_io_pipe_phv_out_data_60; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_61 = pipe12_io_pipe_phv_out_data_61; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_62 = pipe12_io_pipe_phv_out_data_62; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_63 = pipe12_io_pipe_phv_out_data_63; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_64 = pipe12_io_pipe_phv_out_data_64; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_65 = pipe12_io_pipe_phv_out_data_65; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_66 = pipe12_io_pipe_phv_out_data_66; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_67 = pipe12_io_pipe_phv_out_data_67; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_68 = pipe12_io_pipe_phv_out_data_68; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_69 = pipe12_io_pipe_phv_out_data_69; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_70 = pipe12_io_pipe_phv_out_data_70; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_71 = pipe12_io_pipe_phv_out_data_71; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_72 = pipe12_io_pipe_phv_out_data_72; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_73 = pipe12_io_pipe_phv_out_data_73; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_74 = pipe12_io_pipe_phv_out_data_74; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_75 = pipe12_io_pipe_phv_out_data_75; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_76 = pipe12_io_pipe_phv_out_data_76; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_77 = pipe12_io_pipe_phv_out_data_77; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_78 = pipe12_io_pipe_phv_out_data_78; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_79 = pipe12_io_pipe_phv_out_data_79; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_80 = pipe12_io_pipe_phv_out_data_80; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_81 = pipe12_io_pipe_phv_out_data_81; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_82 = pipe12_io_pipe_phv_out_data_82; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_83 = pipe12_io_pipe_phv_out_data_83; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_84 = pipe12_io_pipe_phv_out_data_84; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_85 = pipe12_io_pipe_phv_out_data_85; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_86 = pipe12_io_pipe_phv_out_data_86; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_87 = pipe12_io_pipe_phv_out_data_87; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_88 = pipe12_io_pipe_phv_out_data_88; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_89 = pipe12_io_pipe_phv_out_data_89; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_90 = pipe12_io_pipe_phv_out_data_90; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_91 = pipe12_io_pipe_phv_out_data_91; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_92 = pipe12_io_pipe_phv_out_data_92; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_93 = pipe12_io_pipe_phv_out_data_93; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_94 = pipe12_io_pipe_phv_out_data_94; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_95 = pipe12_io_pipe_phv_out_data_95; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_96 = pipe12_io_pipe_phv_out_data_96; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_97 = pipe12_io_pipe_phv_out_data_97; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_98 = pipe12_io_pipe_phv_out_data_98; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_99 = pipe12_io_pipe_phv_out_data_99; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_100 = pipe12_io_pipe_phv_out_data_100; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_101 = pipe12_io_pipe_phv_out_data_101; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_102 = pipe12_io_pipe_phv_out_data_102; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_103 = pipe12_io_pipe_phv_out_data_103; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_104 = pipe12_io_pipe_phv_out_data_104; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_105 = pipe12_io_pipe_phv_out_data_105; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_106 = pipe12_io_pipe_phv_out_data_106; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_107 = pipe12_io_pipe_phv_out_data_107; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_108 = pipe12_io_pipe_phv_out_data_108; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_109 = pipe12_io_pipe_phv_out_data_109; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_110 = pipe12_io_pipe_phv_out_data_110; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_111 = pipe12_io_pipe_phv_out_data_111; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_112 = pipe12_io_pipe_phv_out_data_112; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_113 = pipe12_io_pipe_phv_out_data_113; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_114 = pipe12_io_pipe_phv_out_data_114; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_115 = pipe12_io_pipe_phv_out_data_115; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_116 = pipe12_io_pipe_phv_out_data_116; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_117 = pipe12_io_pipe_phv_out_data_117; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_118 = pipe12_io_pipe_phv_out_data_118; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_119 = pipe12_io_pipe_phv_out_data_119; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_120 = pipe12_io_pipe_phv_out_data_120; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_121 = pipe12_io_pipe_phv_out_data_121; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_122 = pipe12_io_pipe_phv_out_data_122; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_123 = pipe12_io_pipe_phv_out_data_123; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_124 = pipe12_io_pipe_phv_out_data_124; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_125 = pipe12_io_pipe_phv_out_data_125; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_126 = pipe12_io_pipe_phv_out_data_126; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_127 = pipe12_io_pipe_phv_out_data_127; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_128 = pipe12_io_pipe_phv_out_data_128; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_129 = pipe12_io_pipe_phv_out_data_129; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_130 = pipe12_io_pipe_phv_out_data_130; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_131 = pipe12_io_pipe_phv_out_data_131; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_132 = pipe12_io_pipe_phv_out_data_132; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_133 = pipe12_io_pipe_phv_out_data_133; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_134 = pipe12_io_pipe_phv_out_data_134; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_135 = pipe12_io_pipe_phv_out_data_135; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_136 = pipe12_io_pipe_phv_out_data_136; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_137 = pipe12_io_pipe_phv_out_data_137; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_138 = pipe12_io_pipe_phv_out_data_138; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_139 = pipe12_io_pipe_phv_out_data_139; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_140 = pipe12_io_pipe_phv_out_data_140; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_141 = pipe12_io_pipe_phv_out_data_141; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_142 = pipe12_io_pipe_phv_out_data_142; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_143 = pipe12_io_pipe_phv_out_data_143; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_144 = pipe12_io_pipe_phv_out_data_144; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_145 = pipe12_io_pipe_phv_out_data_145; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_146 = pipe12_io_pipe_phv_out_data_146; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_147 = pipe12_io_pipe_phv_out_data_147; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_148 = pipe12_io_pipe_phv_out_data_148; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_149 = pipe12_io_pipe_phv_out_data_149; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_150 = pipe12_io_pipe_phv_out_data_150; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_151 = pipe12_io_pipe_phv_out_data_151; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_152 = pipe12_io_pipe_phv_out_data_152; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_153 = pipe12_io_pipe_phv_out_data_153; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_154 = pipe12_io_pipe_phv_out_data_154; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_155 = pipe12_io_pipe_phv_out_data_155; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_156 = pipe12_io_pipe_phv_out_data_156; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_157 = pipe12_io_pipe_phv_out_data_157; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_158 = pipe12_io_pipe_phv_out_data_158; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_159 = pipe12_io_pipe_phv_out_data_159; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_160 = pipe12_io_pipe_phv_out_data_160; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_161 = pipe12_io_pipe_phv_out_data_161; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_162 = pipe12_io_pipe_phv_out_data_162; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_163 = pipe12_io_pipe_phv_out_data_163; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_164 = pipe12_io_pipe_phv_out_data_164; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_165 = pipe12_io_pipe_phv_out_data_165; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_166 = pipe12_io_pipe_phv_out_data_166; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_167 = pipe12_io_pipe_phv_out_data_167; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_168 = pipe12_io_pipe_phv_out_data_168; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_169 = pipe12_io_pipe_phv_out_data_169; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_170 = pipe12_io_pipe_phv_out_data_170; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_171 = pipe12_io_pipe_phv_out_data_171; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_172 = pipe12_io_pipe_phv_out_data_172; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_173 = pipe12_io_pipe_phv_out_data_173; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_174 = pipe12_io_pipe_phv_out_data_174; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_175 = pipe12_io_pipe_phv_out_data_175; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_176 = pipe12_io_pipe_phv_out_data_176; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_177 = pipe12_io_pipe_phv_out_data_177; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_178 = pipe12_io_pipe_phv_out_data_178; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_179 = pipe12_io_pipe_phv_out_data_179; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_180 = pipe12_io_pipe_phv_out_data_180; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_181 = pipe12_io_pipe_phv_out_data_181; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_182 = pipe12_io_pipe_phv_out_data_182; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_183 = pipe12_io_pipe_phv_out_data_183; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_184 = pipe12_io_pipe_phv_out_data_184; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_185 = pipe12_io_pipe_phv_out_data_185; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_186 = pipe12_io_pipe_phv_out_data_186; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_187 = pipe12_io_pipe_phv_out_data_187; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_188 = pipe12_io_pipe_phv_out_data_188; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_189 = pipe12_io_pipe_phv_out_data_189; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_190 = pipe12_io_pipe_phv_out_data_190; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_191 = pipe12_io_pipe_phv_out_data_191; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_192 = pipe12_io_pipe_phv_out_data_192; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_193 = pipe12_io_pipe_phv_out_data_193; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_194 = pipe12_io_pipe_phv_out_data_194; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_195 = pipe12_io_pipe_phv_out_data_195; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_196 = pipe12_io_pipe_phv_out_data_196; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_197 = pipe12_io_pipe_phv_out_data_197; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_198 = pipe12_io_pipe_phv_out_data_198; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_199 = pipe12_io_pipe_phv_out_data_199; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_200 = pipe12_io_pipe_phv_out_data_200; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_201 = pipe12_io_pipe_phv_out_data_201; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_202 = pipe12_io_pipe_phv_out_data_202; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_203 = pipe12_io_pipe_phv_out_data_203; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_204 = pipe12_io_pipe_phv_out_data_204; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_205 = pipe12_io_pipe_phv_out_data_205; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_206 = pipe12_io_pipe_phv_out_data_206; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_207 = pipe12_io_pipe_phv_out_data_207; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_208 = pipe12_io_pipe_phv_out_data_208; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_209 = pipe12_io_pipe_phv_out_data_209; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_210 = pipe12_io_pipe_phv_out_data_210; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_211 = pipe12_io_pipe_phv_out_data_211; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_212 = pipe12_io_pipe_phv_out_data_212; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_213 = pipe12_io_pipe_phv_out_data_213; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_214 = pipe12_io_pipe_phv_out_data_214; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_215 = pipe12_io_pipe_phv_out_data_215; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_216 = pipe12_io_pipe_phv_out_data_216; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_217 = pipe12_io_pipe_phv_out_data_217; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_218 = pipe12_io_pipe_phv_out_data_218; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_219 = pipe12_io_pipe_phv_out_data_219; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_220 = pipe12_io_pipe_phv_out_data_220; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_221 = pipe12_io_pipe_phv_out_data_221; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_222 = pipe12_io_pipe_phv_out_data_222; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_223 = pipe12_io_pipe_phv_out_data_223; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_224 = pipe12_io_pipe_phv_out_data_224; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_225 = pipe12_io_pipe_phv_out_data_225; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_226 = pipe12_io_pipe_phv_out_data_226; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_227 = pipe12_io_pipe_phv_out_data_227; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_228 = pipe12_io_pipe_phv_out_data_228; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_229 = pipe12_io_pipe_phv_out_data_229; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_230 = pipe12_io_pipe_phv_out_data_230; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_231 = pipe12_io_pipe_phv_out_data_231; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_232 = pipe12_io_pipe_phv_out_data_232; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_233 = pipe12_io_pipe_phv_out_data_233; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_234 = pipe12_io_pipe_phv_out_data_234; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_235 = pipe12_io_pipe_phv_out_data_235; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_236 = pipe12_io_pipe_phv_out_data_236; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_237 = pipe12_io_pipe_phv_out_data_237; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_238 = pipe12_io_pipe_phv_out_data_238; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_239 = pipe12_io_pipe_phv_out_data_239; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_240 = pipe12_io_pipe_phv_out_data_240; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_241 = pipe12_io_pipe_phv_out_data_241; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_242 = pipe12_io_pipe_phv_out_data_242; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_243 = pipe12_io_pipe_phv_out_data_243; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_244 = pipe12_io_pipe_phv_out_data_244; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_245 = pipe12_io_pipe_phv_out_data_245; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_246 = pipe12_io_pipe_phv_out_data_246; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_247 = pipe12_io_pipe_phv_out_data_247; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_248 = pipe12_io_pipe_phv_out_data_248; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_249 = pipe12_io_pipe_phv_out_data_249; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_250 = pipe12_io_pipe_phv_out_data_250; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_251 = pipe12_io_pipe_phv_out_data_251; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_252 = pipe12_io_pipe_phv_out_data_252; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_253 = pipe12_io_pipe_phv_out_data_253; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_254 = pipe12_io_pipe_phv_out_data_254; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_255 = pipe12_io_pipe_phv_out_data_255; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_256 = pipe12_io_pipe_phv_out_data_256; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_257 = pipe12_io_pipe_phv_out_data_257; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_258 = pipe12_io_pipe_phv_out_data_258; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_259 = pipe12_io_pipe_phv_out_data_259; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_260 = pipe12_io_pipe_phv_out_data_260; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_261 = pipe12_io_pipe_phv_out_data_261; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_262 = pipe12_io_pipe_phv_out_data_262; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_263 = pipe12_io_pipe_phv_out_data_263; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_264 = pipe12_io_pipe_phv_out_data_264; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_265 = pipe12_io_pipe_phv_out_data_265; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_266 = pipe12_io_pipe_phv_out_data_266; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_267 = pipe12_io_pipe_phv_out_data_267; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_268 = pipe12_io_pipe_phv_out_data_268; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_269 = pipe12_io_pipe_phv_out_data_269; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_270 = pipe12_io_pipe_phv_out_data_270; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_271 = pipe12_io_pipe_phv_out_data_271; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_272 = pipe12_io_pipe_phv_out_data_272; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_273 = pipe12_io_pipe_phv_out_data_273; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_274 = pipe12_io_pipe_phv_out_data_274; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_275 = pipe12_io_pipe_phv_out_data_275; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_276 = pipe12_io_pipe_phv_out_data_276; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_277 = pipe12_io_pipe_phv_out_data_277; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_278 = pipe12_io_pipe_phv_out_data_278; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_279 = pipe12_io_pipe_phv_out_data_279; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_280 = pipe12_io_pipe_phv_out_data_280; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_281 = pipe12_io_pipe_phv_out_data_281; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_282 = pipe12_io_pipe_phv_out_data_282; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_283 = pipe12_io_pipe_phv_out_data_283; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_284 = pipe12_io_pipe_phv_out_data_284; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_285 = pipe12_io_pipe_phv_out_data_285; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_286 = pipe12_io_pipe_phv_out_data_286; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_287 = pipe12_io_pipe_phv_out_data_287; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_288 = pipe12_io_pipe_phv_out_data_288; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_289 = pipe12_io_pipe_phv_out_data_289; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_290 = pipe12_io_pipe_phv_out_data_290; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_291 = pipe12_io_pipe_phv_out_data_291; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_292 = pipe12_io_pipe_phv_out_data_292; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_293 = pipe12_io_pipe_phv_out_data_293; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_294 = pipe12_io_pipe_phv_out_data_294; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_295 = pipe12_io_pipe_phv_out_data_295; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_296 = pipe12_io_pipe_phv_out_data_296; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_297 = pipe12_io_pipe_phv_out_data_297; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_298 = pipe12_io_pipe_phv_out_data_298; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_299 = pipe12_io_pipe_phv_out_data_299; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_300 = pipe12_io_pipe_phv_out_data_300; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_301 = pipe12_io_pipe_phv_out_data_301; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_302 = pipe12_io_pipe_phv_out_data_302; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_303 = pipe12_io_pipe_phv_out_data_303; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_304 = pipe12_io_pipe_phv_out_data_304; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_305 = pipe12_io_pipe_phv_out_data_305; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_306 = pipe12_io_pipe_phv_out_data_306; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_307 = pipe12_io_pipe_phv_out_data_307; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_308 = pipe12_io_pipe_phv_out_data_308; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_309 = pipe12_io_pipe_phv_out_data_309; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_310 = pipe12_io_pipe_phv_out_data_310; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_311 = pipe12_io_pipe_phv_out_data_311; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_312 = pipe12_io_pipe_phv_out_data_312; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_313 = pipe12_io_pipe_phv_out_data_313; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_314 = pipe12_io_pipe_phv_out_data_314; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_315 = pipe12_io_pipe_phv_out_data_315; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_316 = pipe12_io_pipe_phv_out_data_316; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_317 = pipe12_io_pipe_phv_out_data_317; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_318 = pipe12_io_pipe_phv_out_data_318; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_319 = pipe12_io_pipe_phv_out_data_319; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_320 = pipe12_io_pipe_phv_out_data_320; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_321 = pipe12_io_pipe_phv_out_data_321; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_322 = pipe12_io_pipe_phv_out_data_322; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_323 = pipe12_io_pipe_phv_out_data_323; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_324 = pipe12_io_pipe_phv_out_data_324; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_325 = pipe12_io_pipe_phv_out_data_325; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_326 = pipe12_io_pipe_phv_out_data_326; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_327 = pipe12_io_pipe_phv_out_data_327; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_328 = pipe12_io_pipe_phv_out_data_328; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_329 = pipe12_io_pipe_phv_out_data_329; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_330 = pipe12_io_pipe_phv_out_data_330; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_331 = pipe12_io_pipe_phv_out_data_331; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_332 = pipe12_io_pipe_phv_out_data_332; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_333 = pipe12_io_pipe_phv_out_data_333; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_334 = pipe12_io_pipe_phv_out_data_334; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_335 = pipe12_io_pipe_phv_out_data_335; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_336 = pipe12_io_pipe_phv_out_data_336; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_337 = pipe12_io_pipe_phv_out_data_337; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_338 = pipe12_io_pipe_phv_out_data_338; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_339 = pipe12_io_pipe_phv_out_data_339; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_340 = pipe12_io_pipe_phv_out_data_340; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_341 = pipe12_io_pipe_phv_out_data_341; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_342 = pipe12_io_pipe_phv_out_data_342; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_343 = pipe12_io_pipe_phv_out_data_343; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_344 = pipe12_io_pipe_phv_out_data_344; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_345 = pipe12_io_pipe_phv_out_data_345; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_346 = pipe12_io_pipe_phv_out_data_346; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_347 = pipe12_io_pipe_phv_out_data_347; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_348 = pipe12_io_pipe_phv_out_data_348; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_349 = pipe12_io_pipe_phv_out_data_349; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_350 = pipe12_io_pipe_phv_out_data_350; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_351 = pipe12_io_pipe_phv_out_data_351; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_352 = pipe12_io_pipe_phv_out_data_352; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_353 = pipe12_io_pipe_phv_out_data_353; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_354 = pipe12_io_pipe_phv_out_data_354; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_355 = pipe12_io_pipe_phv_out_data_355; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_356 = pipe12_io_pipe_phv_out_data_356; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_357 = pipe12_io_pipe_phv_out_data_357; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_358 = pipe12_io_pipe_phv_out_data_358; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_359 = pipe12_io_pipe_phv_out_data_359; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_360 = pipe12_io_pipe_phv_out_data_360; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_361 = pipe12_io_pipe_phv_out_data_361; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_362 = pipe12_io_pipe_phv_out_data_362; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_363 = pipe12_io_pipe_phv_out_data_363; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_364 = pipe12_io_pipe_phv_out_data_364; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_365 = pipe12_io_pipe_phv_out_data_365; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_366 = pipe12_io_pipe_phv_out_data_366; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_367 = pipe12_io_pipe_phv_out_data_367; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_368 = pipe12_io_pipe_phv_out_data_368; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_369 = pipe12_io_pipe_phv_out_data_369; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_370 = pipe12_io_pipe_phv_out_data_370; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_371 = pipe12_io_pipe_phv_out_data_371; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_372 = pipe12_io_pipe_phv_out_data_372; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_373 = pipe12_io_pipe_phv_out_data_373; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_374 = pipe12_io_pipe_phv_out_data_374; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_375 = pipe12_io_pipe_phv_out_data_375; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_376 = pipe12_io_pipe_phv_out_data_376; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_377 = pipe12_io_pipe_phv_out_data_377; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_378 = pipe12_io_pipe_phv_out_data_378; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_379 = pipe12_io_pipe_phv_out_data_379; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_380 = pipe12_io_pipe_phv_out_data_380; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_381 = pipe12_io_pipe_phv_out_data_381; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_382 = pipe12_io_pipe_phv_out_data_382; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_383 = pipe12_io_pipe_phv_out_data_383; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_384 = pipe12_io_pipe_phv_out_data_384; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_385 = pipe12_io_pipe_phv_out_data_385; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_386 = pipe12_io_pipe_phv_out_data_386; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_387 = pipe12_io_pipe_phv_out_data_387; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_388 = pipe12_io_pipe_phv_out_data_388; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_389 = pipe12_io_pipe_phv_out_data_389; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_390 = pipe12_io_pipe_phv_out_data_390; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_391 = pipe12_io_pipe_phv_out_data_391; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_392 = pipe12_io_pipe_phv_out_data_392; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_393 = pipe12_io_pipe_phv_out_data_393; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_394 = pipe12_io_pipe_phv_out_data_394; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_395 = pipe12_io_pipe_phv_out_data_395; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_396 = pipe12_io_pipe_phv_out_data_396; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_397 = pipe12_io_pipe_phv_out_data_397; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_398 = pipe12_io_pipe_phv_out_data_398; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_399 = pipe12_io_pipe_phv_out_data_399; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_400 = pipe12_io_pipe_phv_out_data_400; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_401 = pipe12_io_pipe_phv_out_data_401; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_402 = pipe12_io_pipe_phv_out_data_402; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_403 = pipe12_io_pipe_phv_out_data_403; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_404 = pipe12_io_pipe_phv_out_data_404; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_405 = pipe12_io_pipe_phv_out_data_405; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_406 = pipe12_io_pipe_phv_out_data_406; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_407 = pipe12_io_pipe_phv_out_data_407; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_408 = pipe12_io_pipe_phv_out_data_408; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_409 = pipe12_io_pipe_phv_out_data_409; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_410 = pipe12_io_pipe_phv_out_data_410; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_411 = pipe12_io_pipe_phv_out_data_411; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_412 = pipe12_io_pipe_phv_out_data_412; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_413 = pipe12_io_pipe_phv_out_data_413; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_414 = pipe12_io_pipe_phv_out_data_414; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_415 = pipe12_io_pipe_phv_out_data_415; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_416 = pipe12_io_pipe_phv_out_data_416; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_417 = pipe12_io_pipe_phv_out_data_417; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_418 = pipe12_io_pipe_phv_out_data_418; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_419 = pipe12_io_pipe_phv_out_data_419; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_420 = pipe12_io_pipe_phv_out_data_420; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_421 = pipe12_io_pipe_phv_out_data_421; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_422 = pipe12_io_pipe_phv_out_data_422; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_423 = pipe12_io_pipe_phv_out_data_423; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_424 = pipe12_io_pipe_phv_out_data_424; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_425 = pipe12_io_pipe_phv_out_data_425; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_426 = pipe12_io_pipe_phv_out_data_426; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_427 = pipe12_io_pipe_phv_out_data_427; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_428 = pipe12_io_pipe_phv_out_data_428; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_429 = pipe12_io_pipe_phv_out_data_429; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_430 = pipe12_io_pipe_phv_out_data_430; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_431 = pipe12_io_pipe_phv_out_data_431; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_432 = pipe12_io_pipe_phv_out_data_432; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_433 = pipe12_io_pipe_phv_out_data_433; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_434 = pipe12_io_pipe_phv_out_data_434; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_435 = pipe12_io_pipe_phv_out_data_435; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_436 = pipe12_io_pipe_phv_out_data_436; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_437 = pipe12_io_pipe_phv_out_data_437; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_438 = pipe12_io_pipe_phv_out_data_438; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_439 = pipe12_io_pipe_phv_out_data_439; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_440 = pipe12_io_pipe_phv_out_data_440; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_441 = pipe12_io_pipe_phv_out_data_441; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_442 = pipe12_io_pipe_phv_out_data_442; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_443 = pipe12_io_pipe_phv_out_data_443; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_444 = pipe12_io_pipe_phv_out_data_444; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_445 = pipe12_io_pipe_phv_out_data_445; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_446 = pipe12_io_pipe_phv_out_data_446; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_447 = pipe12_io_pipe_phv_out_data_447; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_448 = pipe12_io_pipe_phv_out_data_448; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_449 = pipe12_io_pipe_phv_out_data_449; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_450 = pipe12_io_pipe_phv_out_data_450; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_451 = pipe12_io_pipe_phv_out_data_451; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_452 = pipe12_io_pipe_phv_out_data_452; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_453 = pipe12_io_pipe_phv_out_data_453; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_454 = pipe12_io_pipe_phv_out_data_454; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_455 = pipe12_io_pipe_phv_out_data_455; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_456 = pipe12_io_pipe_phv_out_data_456; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_457 = pipe12_io_pipe_phv_out_data_457; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_458 = pipe12_io_pipe_phv_out_data_458; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_459 = pipe12_io_pipe_phv_out_data_459; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_460 = pipe12_io_pipe_phv_out_data_460; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_461 = pipe12_io_pipe_phv_out_data_461; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_462 = pipe12_io_pipe_phv_out_data_462; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_463 = pipe12_io_pipe_phv_out_data_463; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_464 = pipe12_io_pipe_phv_out_data_464; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_465 = pipe12_io_pipe_phv_out_data_465; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_466 = pipe12_io_pipe_phv_out_data_466; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_467 = pipe12_io_pipe_phv_out_data_467; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_468 = pipe12_io_pipe_phv_out_data_468; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_469 = pipe12_io_pipe_phv_out_data_469; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_470 = pipe12_io_pipe_phv_out_data_470; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_471 = pipe12_io_pipe_phv_out_data_471; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_472 = pipe12_io_pipe_phv_out_data_472; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_473 = pipe12_io_pipe_phv_out_data_473; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_474 = pipe12_io_pipe_phv_out_data_474; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_475 = pipe12_io_pipe_phv_out_data_475; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_476 = pipe12_io_pipe_phv_out_data_476; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_477 = pipe12_io_pipe_phv_out_data_477; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_478 = pipe12_io_pipe_phv_out_data_478; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_479 = pipe12_io_pipe_phv_out_data_479; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_480 = pipe12_io_pipe_phv_out_data_480; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_481 = pipe12_io_pipe_phv_out_data_481; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_482 = pipe12_io_pipe_phv_out_data_482; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_483 = pipe12_io_pipe_phv_out_data_483; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_484 = pipe12_io_pipe_phv_out_data_484; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_485 = pipe12_io_pipe_phv_out_data_485; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_486 = pipe12_io_pipe_phv_out_data_486; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_487 = pipe12_io_pipe_phv_out_data_487; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_488 = pipe12_io_pipe_phv_out_data_488; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_489 = pipe12_io_pipe_phv_out_data_489; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_490 = pipe12_io_pipe_phv_out_data_490; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_491 = pipe12_io_pipe_phv_out_data_491; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_492 = pipe12_io_pipe_phv_out_data_492; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_493 = pipe12_io_pipe_phv_out_data_493; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_494 = pipe12_io_pipe_phv_out_data_494; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_495 = pipe12_io_pipe_phv_out_data_495; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_496 = pipe12_io_pipe_phv_out_data_496; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_497 = pipe12_io_pipe_phv_out_data_497; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_498 = pipe12_io_pipe_phv_out_data_498; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_499 = pipe12_io_pipe_phv_out_data_499; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_500 = pipe12_io_pipe_phv_out_data_500; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_501 = pipe12_io_pipe_phv_out_data_501; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_502 = pipe12_io_pipe_phv_out_data_502; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_503 = pipe12_io_pipe_phv_out_data_503; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_504 = pipe12_io_pipe_phv_out_data_504; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_505 = pipe12_io_pipe_phv_out_data_505; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_506 = pipe12_io_pipe_phv_out_data_506; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_507 = pipe12_io_pipe_phv_out_data_507; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_508 = pipe12_io_pipe_phv_out_data_508; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_509 = pipe12_io_pipe_phv_out_data_509; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_510 = pipe12_io_pipe_phv_out_data_510; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_511 = pipe12_io_pipe_phv_out_data_511; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_0 = pipe12_io_pipe_phv_out_header_0; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_1 = pipe12_io_pipe_phv_out_header_1; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_2 = pipe12_io_pipe_phv_out_header_2; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_3 = pipe12_io_pipe_phv_out_header_3; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_4 = pipe12_io_pipe_phv_out_header_4; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_5 = pipe12_io_pipe_phv_out_header_5; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_6 = pipe12_io_pipe_phv_out_header_6; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_7 = pipe12_io_pipe_phv_out_header_7; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_8 = pipe12_io_pipe_phv_out_header_8; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_9 = pipe12_io_pipe_phv_out_header_9; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_10 = pipe12_io_pipe_phv_out_header_10; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_11 = pipe12_io_pipe_phv_out_header_11; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_12 = pipe12_io_pipe_phv_out_header_12; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_13 = pipe12_io_pipe_phv_out_header_13; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_14 = pipe12_io_pipe_phv_out_header_14; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_15 = pipe12_io_pipe_phv_out_header_15; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_parse_current_state = pipe12_io_pipe_phv_out_parse_current_state; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_parse_current_offset = pipe12_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_parse_transition_field = pipe12_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_next_processor_id = pipe12_io_pipe_phv_out_next_processor_id; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_next_config_id = pipe12_io_pipe_phv_out_next_config_id; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_is_valid_processor = pipe12_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 388:27]
  assign io_hit = pipe12_io_hit; // @[matcher.scala 389:27]
  assign io_match_value = pipe12_io_match_value; // @[matcher.scala 390:27]
  assign io_mem_cluster_0_en = pipe10_io_mem_cluster_0_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_0_addr = pipe10_io_mem_cluster_0_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_1_en = pipe10_io_mem_cluster_1_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_1_addr = pipe10_io_mem_cluster_1_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_2_en = pipe10_io_mem_cluster_2_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_2_addr = pipe10_io_mem_cluster_2_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_3_en = pipe10_io_mem_cluster_3_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_3_addr = pipe10_io_mem_cluster_3_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_4_en = pipe10_io_mem_cluster_4_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_4_addr = pipe10_io_mem_cluster_4_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_5_en = pipe10_io_mem_cluster_5_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_5_addr = pipe10_io_mem_cluster_5_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_6_en = pipe10_io_mem_cluster_6_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_6_addr = pipe10_io_mem_cluster_6_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_7_en = pipe10_io_mem_cluster_7_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_7_addr = pipe10_io_mem_cluster_7_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_8_en = pipe10_io_mem_cluster_8_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_8_addr = pipe10_io_mem_cluster_8_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_9_en = pipe10_io_mem_cluster_9_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_9_addr = pipe10_io_mem_cluster_9_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_10_en = pipe10_io_mem_cluster_10_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_10_addr = pipe10_io_mem_cluster_10_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_11_en = pipe10_io_mem_cluster_11_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_11_addr = pipe10_io_mem_cluster_11_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_12_en = pipe10_io_mem_cluster_12_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_12_addr = pipe10_io_mem_cluster_12_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_13_en = pipe10_io_mem_cluster_13_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_13_addr = pipe10_io_mem_cluster_13_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_14_en = pipe10_io_mem_cluster_14_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_14_addr = pipe10_io_mem_cluster_14_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_15_en = pipe10_io_mem_cluster_15_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_15_addr = pipe10_io_mem_cluster_15_addr; // @[matcher.scala 375:27]
  assign pipe1_clock = clock;
  assign pipe1_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_160 = io_pipe_phv_in_data_160; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_161 = io_pipe_phv_in_data_161; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_162 = io_pipe_phv_in_data_162; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_163 = io_pipe_phv_in_data_163; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_164 = io_pipe_phv_in_data_164; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_165 = io_pipe_phv_in_data_165; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_166 = io_pipe_phv_in_data_166; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_167 = io_pipe_phv_in_data_167; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_168 = io_pipe_phv_in_data_168; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_169 = io_pipe_phv_in_data_169; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_170 = io_pipe_phv_in_data_170; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_171 = io_pipe_phv_in_data_171; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_172 = io_pipe_phv_in_data_172; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_173 = io_pipe_phv_in_data_173; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_174 = io_pipe_phv_in_data_174; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_175 = io_pipe_phv_in_data_175; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_176 = io_pipe_phv_in_data_176; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_177 = io_pipe_phv_in_data_177; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_178 = io_pipe_phv_in_data_178; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_179 = io_pipe_phv_in_data_179; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_180 = io_pipe_phv_in_data_180; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_181 = io_pipe_phv_in_data_181; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_182 = io_pipe_phv_in_data_182; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_183 = io_pipe_phv_in_data_183; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_184 = io_pipe_phv_in_data_184; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_185 = io_pipe_phv_in_data_185; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_186 = io_pipe_phv_in_data_186; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_187 = io_pipe_phv_in_data_187; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_188 = io_pipe_phv_in_data_188; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_189 = io_pipe_phv_in_data_189; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_190 = io_pipe_phv_in_data_190; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_191 = io_pipe_phv_in_data_191; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_192 = io_pipe_phv_in_data_192; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_193 = io_pipe_phv_in_data_193; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_194 = io_pipe_phv_in_data_194; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_195 = io_pipe_phv_in_data_195; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_196 = io_pipe_phv_in_data_196; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_197 = io_pipe_phv_in_data_197; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_198 = io_pipe_phv_in_data_198; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_199 = io_pipe_phv_in_data_199; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_200 = io_pipe_phv_in_data_200; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_201 = io_pipe_phv_in_data_201; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_202 = io_pipe_phv_in_data_202; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_203 = io_pipe_phv_in_data_203; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_204 = io_pipe_phv_in_data_204; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_205 = io_pipe_phv_in_data_205; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_206 = io_pipe_phv_in_data_206; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_207 = io_pipe_phv_in_data_207; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_208 = io_pipe_phv_in_data_208; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_209 = io_pipe_phv_in_data_209; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_210 = io_pipe_phv_in_data_210; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_211 = io_pipe_phv_in_data_211; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_212 = io_pipe_phv_in_data_212; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_213 = io_pipe_phv_in_data_213; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_214 = io_pipe_phv_in_data_214; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_215 = io_pipe_phv_in_data_215; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_216 = io_pipe_phv_in_data_216; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_217 = io_pipe_phv_in_data_217; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_218 = io_pipe_phv_in_data_218; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_219 = io_pipe_phv_in_data_219; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_220 = io_pipe_phv_in_data_220; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_221 = io_pipe_phv_in_data_221; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_222 = io_pipe_phv_in_data_222; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_223 = io_pipe_phv_in_data_223; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_224 = io_pipe_phv_in_data_224; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_225 = io_pipe_phv_in_data_225; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_226 = io_pipe_phv_in_data_226; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_227 = io_pipe_phv_in_data_227; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_228 = io_pipe_phv_in_data_228; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_229 = io_pipe_phv_in_data_229; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_230 = io_pipe_phv_in_data_230; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_231 = io_pipe_phv_in_data_231; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_232 = io_pipe_phv_in_data_232; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_233 = io_pipe_phv_in_data_233; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_234 = io_pipe_phv_in_data_234; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_235 = io_pipe_phv_in_data_235; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_236 = io_pipe_phv_in_data_236; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_237 = io_pipe_phv_in_data_237; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_238 = io_pipe_phv_in_data_238; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_239 = io_pipe_phv_in_data_239; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_240 = io_pipe_phv_in_data_240; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_241 = io_pipe_phv_in_data_241; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_242 = io_pipe_phv_in_data_242; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_243 = io_pipe_phv_in_data_243; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_244 = io_pipe_phv_in_data_244; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_245 = io_pipe_phv_in_data_245; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_246 = io_pipe_phv_in_data_246; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_247 = io_pipe_phv_in_data_247; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_248 = io_pipe_phv_in_data_248; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_249 = io_pipe_phv_in_data_249; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_250 = io_pipe_phv_in_data_250; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_251 = io_pipe_phv_in_data_251; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_252 = io_pipe_phv_in_data_252; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_253 = io_pipe_phv_in_data_253; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_254 = io_pipe_phv_in_data_254; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_255 = io_pipe_phv_in_data_255; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_256 = io_pipe_phv_in_data_256; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_257 = io_pipe_phv_in_data_257; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_258 = io_pipe_phv_in_data_258; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_259 = io_pipe_phv_in_data_259; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_260 = io_pipe_phv_in_data_260; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_261 = io_pipe_phv_in_data_261; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_262 = io_pipe_phv_in_data_262; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_263 = io_pipe_phv_in_data_263; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_264 = io_pipe_phv_in_data_264; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_265 = io_pipe_phv_in_data_265; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_266 = io_pipe_phv_in_data_266; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_267 = io_pipe_phv_in_data_267; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_268 = io_pipe_phv_in_data_268; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_269 = io_pipe_phv_in_data_269; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_270 = io_pipe_phv_in_data_270; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_271 = io_pipe_phv_in_data_271; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_272 = io_pipe_phv_in_data_272; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_273 = io_pipe_phv_in_data_273; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_274 = io_pipe_phv_in_data_274; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_275 = io_pipe_phv_in_data_275; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_276 = io_pipe_phv_in_data_276; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_277 = io_pipe_phv_in_data_277; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_278 = io_pipe_phv_in_data_278; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_279 = io_pipe_phv_in_data_279; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_280 = io_pipe_phv_in_data_280; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_281 = io_pipe_phv_in_data_281; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_282 = io_pipe_phv_in_data_282; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_283 = io_pipe_phv_in_data_283; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_284 = io_pipe_phv_in_data_284; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_285 = io_pipe_phv_in_data_285; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_286 = io_pipe_phv_in_data_286; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_287 = io_pipe_phv_in_data_287; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_288 = io_pipe_phv_in_data_288; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_289 = io_pipe_phv_in_data_289; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_290 = io_pipe_phv_in_data_290; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_291 = io_pipe_phv_in_data_291; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_292 = io_pipe_phv_in_data_292; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_293 = io_pipe_phv_in_data_293; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_294 = io_pipe_phv_in_data_294; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_295 = io_pipe_phv_in_data_295; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_296 = io_pipe_phv_in_data_296; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_297 = io_pipe_phv_in_data_297; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_298 = io_pipe_phv_in_data_298; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_299 = io_pipe_phv_in_data_299; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_300 = io_pipe_phv_in_data_300; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_301 = io_pipe_phv_in_data_301; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_302 = io_pipe_phv_in_data_302; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_303 = io_pipe_phv_in_data_303; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_304 = io_pipe_phv_in_data_304; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_305 = io_pipe_phv_in_data_305; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_306 = io_pipe_phv_in_data_306; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_307 = io_pipe_phv_in_data_307; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_308 = io_pipe_phv_in_data_308; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_309 = io_pipe_phv_in_data_309; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_310 = io_pipe_phv_in_data_310; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_311 = io_pipe_phv_in_data_311; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_312 = io_pipe_phv_in_data_312; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_313 = io_pipe_phv_in_data_313; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_314 = io_pipe_phv_in_data_314; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_315 = io_pipe_phv_in_data_315; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_316 = io_pipe_phv_in_data_316; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_317 = io_pipe_phv_in_data_317; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_318 = io_pipe_phv_in_data_318; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_319 = io_pipe_phv_in_data_319; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_320 = io_pipe_phv_in_data_320; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_321 = io_pipe_phv_in_data_321; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_322 = io_pipe_phv_in_data_322; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_323 = io_pipe_phv_in_data_323; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_324 = io_pipe_phv_in_data_324; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_325 = io_pipe_phv_in_data_325; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_326 = io_pipe_phv_in_data_326; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_327 = io_pipe_phv_in_data_327; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_328 = io_pipe_phv_in_data_328; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_329 = io_pipe_phv_in_data_329; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_330 = io_pipe_phv_in_data_330; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_331 = io_pipe_phv_in_data_331; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_332 = io_pipe_phv_in_data_332; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_333 = io_pipe_phv_in_data_333; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_334 = io_pipe_phv_in_data_334; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_335 = io_pipe_phv_in_data_335; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_336 = io_pipe_phv_in_data_336; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_337 = io_pipe_phv_in_data_337; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_338 = io_pipe_phv_in_data_338; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_339 = io_pipe_phv_in_data_339; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_340 = io_pipe_phv_in_data_340; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_341 = io_pipe_phv_in_data_341; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_342 = io_pipe_phv_in_data_342; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_343 = io_pipe_phv_in_data_343; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_344 = io_pipe_phv_in_data_344; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_345 = io_pipe_phv_in_data_345; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_346 = io_pipe_phv_in_data_346; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_347 = io_pipe_phv_in_data_347; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_348 = io_pipe_phv_in_data_348; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_349 = io_pipe_phv_in_data_349; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_350 = io_pipe_phv_in_data_350; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_351 = io_pipe_phv_in_data_351; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_352 = io_pipe_phv_in_data_352; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_353 = io_pipe_phv_in_data_353; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_354 = io_pipe_phv_in_data_354; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_355 = io_pipe_phv_in_data_355; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_356 = io_pipe_phv_in_data_356; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_357 = io_pipe_phv_in_data_357; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_358 = io_pipe_phv_in_data_358; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_359 = io_pipe_phv_in_data_359; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_360 = io_pipe_phv_in_data_360; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_361 = io_pipe_phv_in_data_361; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_362 = io_pipe_phv_in_data_362; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_363 = io_pipe_phv_in_data_363; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_364 = io_pipe_phv_in_data_364; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_365 = io_pipe_phv_in_data_365; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_366 = io_pipe_phv_in_data_366; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_367 = io_pipe_phv_in_data_367; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_368 = io_pipe_phv_in_data_368; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_369 = io_pipe_phv_in_data_369; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_370 = io_pipe_phv_in_data_370; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_371 = io_pipe_phv_in_data_371; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_372 = io_pipe_phv_in_data_372; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_373 = io_pipe_phv_in_data_373; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_374 = io_pipe_phv_in_data_374; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_375 = io_pipe_phv_in_data_375; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_376 = io_pipe_phv_in_data_376; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_377 = io_pipe_phv_in_data_377; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_378 = io_pipe_phv_in_data_378; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_379 = io_pipe_phv_in_data_379; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_380 = io_pipe_phv_in_data_380; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_381 = io_pipe_phv_in_data_381; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_382 = io_pipe_phv_in_data_382; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_383 = io_pipe_phv_in_data_383; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_384 = io_pipe_phv_in_data_384; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_385 = io_pipe_phv_in_data_385; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_386 = io_pipe_phv_in_data_386; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_387 = io_pipe_phv_in_data_387; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_388 = io_pipe_phv_in_data_388; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_389 = io_pipe_phv_in_data_389; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_390 = io_pipe_phv_in_data_390; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_391 = io_pipe_phv_in_data_391; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_392 = io_pipe_phv_in_data_392; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_393 = io_pipe_phv_in_data_393; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_394 = io_pipe_phv_in_data_394; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_395 = io_pipe_phv_in_data_395; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_396 = io_pipe_phv_in_data_396; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_397 = io_pipe_phv_in_data_397; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_398 = io_pipe_phv_in_data_398; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_399 = io_pipe_phv_in_data_399; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_400 = io_pipe_phv_in_data_400; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_401 = io_pipe_phv_in_data_401; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_402 = io_pipe_phv_in_data_402; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_403 = io_pipe_phv_in_data_403; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_404 = io_pipe_phv_in_data_404; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_405 = io_pipe_phv_in_data_405; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_406 = io_pipe_phv_in_data_406; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_407 = io_pipe_phv_in_data_407; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_408 = io_pipe_phv_in_data_408; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_409 = io_pipe_phv_in_data_409; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_410 = io_pipe_phv_in_data_410; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_411 = io_pipe_phv_in_data_411; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_412 = io_pipe_phv_in_data_412; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_413 = io_pipe_phv_in_data_413; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_414 = io_pipe_phv_in_data_414; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_415 = io_pipe_phv_in_data_415; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_416 = io_pipe_phv_in_data_416; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_417 = io_pipe_phv_in_data_417; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_418 = io_pipe_phv_in_data_418; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_419 = io_pipe_phv_in_data_419; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_420 = io_pipe_phv_in_data_420; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_421 = io_pipe_phv_in_data_421; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_422 = io_pipe_phv_in_data_422; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_423 = io_pipe_phv_in_data_423; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_424 = io_pipe_phv_in_data_424; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_425 = io_pipe_phv_in_data_425; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_426 = io_pipe_phv_in_data_426; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_427 = io_pipe_phv_in_data_427; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_428 = io_pipe_phv_in_data_428; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_429 = io_pipe_phv_in_data_429; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_430 = io_pipe_phv_in_data_430; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_431 = io_pipe_phv_in_data_431; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_432 = io_pipe_phv_in_data_432; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_433 = io_pipe_phv_in_data_433; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_434 = io_pipe_phv_in_data_434; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_435 = io_pipe_phv_in_data_435; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_436 = io_pipe_phv_in_data_436; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_437 = io_pipe_phv_in_data_437; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_438 = io_pipe_phv_in_data_438; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_439 = io_pipe_phv_in_data_439; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_440 = io_pipe_phv_in_data_440; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_441 = io_pipe_phv_in_data_441; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_442 = io_pipe_phv_in_data_442; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_443 = io_pipe_phv_in_data_443; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_444 = io_pipe_phv_in_data_444; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_445 = io_pipe_phv_in_data_445; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_446 = io_pipe_phv_in_data_446; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_447 = io_pipe_phv_in_data_447; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_448 = io_pipe_phv_in_data_448; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_449 = io_pipe_phv_in_data_449; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_450 = io_pipe_phv_in_data_450; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_451 = io_pipe_phv_in_data_451; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_452 = io_pipe_phv_in_data_452; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_453 = io_pipe_phv_in_data_453; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_454 = io_pipe_phv_in_data_454; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_455 = io_pipe_phv_in_data_455; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_456 = io_pipe_phv_in_data_456; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_457 = io_pipe_phv_in_data_457; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_458 = io_pipe_phv_in_data_458; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_459 = io_pipe_phv_in_data_459; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_460 = io_pipe_phv_in_data_460; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_461 = io_pipe_phv_in_data_461; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_462 = io_pipe_phv_in_data_462; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_463 = io_pipe_phv_in_data_463; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_464 = io_pipe_phv_in_data_464; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_465 = io_pipe_phv_in_data_465; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_466 = io_pipe_phv_in_data_466; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_467 = io_pipe_phv_in_data_467; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_468 = io_pipe_phv_in_data_468; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_469 = io_pipe_phv_in_data_469; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_470 = io_pipe_phv_in_data_470; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_471 = io_pipe_phv_in_data_471; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_472 = io_pipe_phv_in_data_472; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_473 = io_pipe_phv_in_data_473; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_474 = io_pipe_phv_in_data_474; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_475 = io_pipe_phv_in_data_475; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_476 = io_pipe_phv_in_data_476; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_477 = io_pipe_phv_in_data_477; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_478 = io_pipe_phv_in_data_478; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_479 = io_pipe_phv_in_data_479; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_480 = io_pipe_phv_in_data_480; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_481 = io_pipe_phv_in_data_481; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_482 = io_pipe_phv_in_data_482; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_483 = io_pipe_phv_in_data_483; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_484 = io_pipe_phv_in_data_484; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_485 = io_pipe_phv_in_data_485; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_486 = io_pipe_phv_in_data_486; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_487 = io_pipe_phv_in_data_487; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_488 = io_pipe_phv_in_data_488; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_489 = io_pipe_phv_in_data_489; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_490 = io_pipe_phv_in_data_490; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_491 = io_pipe_phv_in_data_491; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_492 = io_pipe_phv_in_data_492; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_493 = io_pipe_phv_in_data_493; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_494 = io_pipe_phv_in_data_494; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_495 = io_pipe_phv_in_data_495; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_496 = io_pipe_phv_in_data_496; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_497 = io_pipe_phv_in_data_497; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_498 = io_pipe_phv_in_data_498; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_499 = io_pipe_phv_in_data_499; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_500 = io_pipe_phv_in_data_500; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_501 = io_pipe_phv_in_data_501; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_502 = io_pipe_phv_in_data_502; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_503 = io_pipe_phv_in_data_503; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_504 = io_pipe_phv_in_data_504; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_505 = io_pipe_phv_in_data_505; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_506 = io_pipe_phv_in_data_506; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_507 = io_pipe_phv_in_data_507; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_508 = io_pipe_phv_in_data_508; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_509 = io_pipe_phv_in_data_509; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_510 = io_pipe_phv_in_data_510; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_511 = io_pipe_phv_in_data_511; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[matcher.scala 351:26]
  assign pipe1_io_key_config_0_header_id = key_config_0_header_id; // @[matcher.scala 352:26]
  assign pipe1_io_key_config_0_internal_offset = key_config_0_internal_offset; // @[matcher.scala 352:26]
  assign pipe1_io_key_config_1_header_id = key_config_1_header_id; // @[matcher.scala 352:26]
  assign pipe1_io_key_config_1_internal_offset = key_config_1_internal_offset; // @[matcher.scala 352:26]
  assign pipe2_clock = clock;
  assign pipe2_io_pipe_phv_in_data_0 = pipe1_io_pipe_phv_out_data_0; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_1 = pipe1_io_pipe_phv_out_data_1; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_2 = pipe1_io_pipe_phv_out_data_2; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_3 = pipe1_io_pipe_phv_out_data_3; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_4 = pipe1_io_pipe_phv_out_data_4; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_5 = pipe1_io_pipe_phv_out_data_5; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_6 = pipe1_io_pipe_phv_out_data_6; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_7 = pipe1_io_pipe_phv_out_data_7; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_8 = pipe1_io_pipe_phv_out_data_8; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_9 = pipe1_io_pipe_phv_out_data_9; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_10 = pipe1_io_pipe_phv_out_data_10; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_11 = pipe1_io_pipe_phv_out_data_11; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_12 = pipe1_io_pipe_phv_out_data_12; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_13 = pipe1_io_pipe_phv_out_data_13; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_14 = pipe1_io_pipe_phv_out_data_14; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_15 = pipe1_io_pipe_phv_out_data_15; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_16 = pipe1_io_pipe_phv_out_data_16; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_17 = pipe1_io_pipe_phv_out_data_17; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_18 = pipe1_io_pipe_phv_out_data_18; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_19 = pipe1_io_pipe_phv_out_data_19; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_20 = pipe1_io_pipe_phv_out_data_20; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_21 = pipe1_io_pipe_phv_out_data_21; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_22 = pipe1_io_pipe_phv_out_data_22; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_23 = pipe1_io_pipe_phv_out_data_23; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_24 = pipe1_io_pipe_phv_out_data_24; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_25 = pipe1_io_pipe_phv_out_data_25; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_26 = pipe1_io_pipe_phv_out_data_26; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_27 = pipe1_io_pipe_phv_out_data_27; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_28 = pipe1_io_pipe_phv_out_data_28; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_29 = pipe1_io_pipe_phv_out_data_29; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_30 = pipe1_io_pipe_phv_out_data_30; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_31 = pipe1_io_pipe_phv_out_data_31; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_32 = pipe1_io_pipe_phv_out_data_32; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_33 = pipe1_io_pipe_phv_out_data_33; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_34 = pipe1_io_pipe_phv_out_data_34; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_35 = pipe1_io_pipe_phv_out_data_35; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_36 = pipe1_io_pipe_phv_out_data_36; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_37 = pipe1_io_pipe_phv_out_data_37; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_38 = pipe1_io_pipe_phv_out_data_38; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_39 = pipe1_io_pipe_phv_out_data_39; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_40 = pipe1_io_pipe_phv_out_data_40; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_41 = pipe1_io_pipe_phv_out_data_41; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_42 = pipe1_io_pipe_phv_out_data_42; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_43 = pipe1_io_pipe_phv_out_data_43; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_44 = pipe1_io_pipe_phv_out_data_44; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_45 = pipe1_io_pipe_phv_out_data_45; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_46 = pipe1_io_pipe_phv_out_data_46; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_47 = pipe1_io_pipe_phv_out_data_47; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_48 = pipe1_io_pipe_phv_out_data_48; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_49 = pipe1_io_pipe_phv_out_data_49; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_50 = pipe1_io_pipe_phv_out_data_50; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_51 = pipe1_io_pipe_phv_out_data_51; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_52 = pipe1_io_pipe_phv_out_data_52; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_53 = pipe1_io_pipe_phv_out_data_53; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_54 = pipe1_io_pipe_phv_out_data_54; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_55 = pipe1_io_pipe_phv_out_data_55; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_56 = pipe1_io_pipe_phv_out_data_56; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_57 = pipe1_io_pipe_phv_out_data_57; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_58 = pipe1_io_pipe_phv_out_data_58; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_59 = pipe1_io_pipe_phv_out_data_59; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_60 = pipe1_io_pipe_phv_out_data_60; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_61 = pipe1_io_pipe_phv_out_data_61; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_62 = pipe1_io_pipe_phv_out_data_62; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_63 = pipe1_io_pipe_phv_out_data_63; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_64 = pipe1_io_pipe_phv_out_data_64; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_65 = pipe1_io_pipe_phv_out_data_65; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_66 = pipe1_io_pipe_phv_out_data_66; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_67 = pipe1_io_pipe_phv_out_data_67; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_68 = pipe1_io_pipe_phv_out_data_68; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_69 = pipe1_io_pipe_phv_out_data_69; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_70 = pipe1_io_pipe_phv_out_data_70; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_71 = pipe1_io_pipe_phv_out_data_71; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_72 = pipe1_io_pipe_phv_out_data_72; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_73 = pipe1_io_pipe_phv_out_data_73; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_74 = pipe1_io_pipe_phv_out_data_74; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_75 = pipe1_io_pipe_phv_out_data_75; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_76 = pipe1_io_pipe_phv_out_data_76; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_77 = pipe1_io_pipe_phv_out_data_77; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_78 = pipe1_io_pipe_phv_out_data_78; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_79 = pipe1_io_pipe_phv_out_data_79; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_80 = pipe1_io_pipe_phv_out_data_80; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_81 = pipe1_io_pipe_phv_out_data_81; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_82 = pipe1_io_pipe_phv_out_data_82; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_83 = pipe1_io_pipe_phv_out_data_83; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_84 = pipe1_io_pipe_phv_out_data_84; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_85 = pipe1_io_pipe_phv_out_data_85; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_86 = pipe1_io_pipe_phv_out_data_86; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_87 = pipe1_io_pipe_phv_out_data_87; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_88 = pipe1_io_pipe_phv_out_data_88; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_89 = pipe1_io_pipe_phv_out_data_89; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_90 = pipe1_io_pipe_phv_out_data_90; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_91 = pipe1_io_pipe_phv_out_data_91; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_92 = pipe1_io_pipe_phv_out_data_92; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_93 = pipe1_io_pipe_phv_out_data_93; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_94 = pipe1_io_pipe_phv_out_data_94; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_95 = pipe1_io_pipe_phv_out_data_95; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_96 = pipe1_io_pipe_phv_out_data_96; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_97 = pipe1_io_pipe_phv_out_data_97; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_98 = pipe1_io_pipe_phv_out_data_98; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_99 = pipe1_io_pipe_phv_out_data_99; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_100 = pipe1_io_pipe_phv_out_data_100; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_101 = pipe1_io_pipe_phv_out_data_101; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_102 = pipe1_io_pipe_phv_out_data_102; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_103 = pipe1_io_pipe_phv_out_data_103; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_104 = pipe1_io_pipe_phv_out_data_104; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_105 = pipe1_io_pipe_phv_out_data_105; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_106 = pipe1_io_pipe_phv_out_data_106; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_107 = pipe1_io_pipe_phv_out_data_107; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_108 = pipe1_io_pipe_phv_out_data_108; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_109 = pipe1_io_pipe_phv_out_data_109; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_110 = pipe1_io_pipe_phv_out_data_110; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_111 = pipe1_io_pipe_phv_out_data_111; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_112 = pipe1_io_pipe_phv_out_data_112; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_113 = pipe1_io_pipe_phv_out_data_113; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_114 = pipe1_io_pipe_phv_out_data_114; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_115 = pipe1_io_pipe_phv_out_data_115; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_116 = pipe1_io_pipe_phv_out_data_116; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_117 = pipe1_io_pipe_phv_out_data_117; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_118 = pipe1_io_pipe_phv_out_data_118; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_119 = pipe1_io_pipe_phv_out_data_119; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_120 = pipe1_io_pipe_phv_out_data_120; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_121 = pipe1_io_pipe_phv_out_data_121; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_122 = pipe1_io_pipe_phv_out_data_122; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_123 = pipe1_io_pipe_phv_out_data_123; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_124 = pipe1_io_pipe_phv_out_data_124; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_125 = pipe1_io_pipe_phv_out_data_125; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_126 = pipe1_io_pipe_phv_out_data_126; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_127 = pipe1_io_pipe_phv_out_data_127; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_128 = pipe1_io_pipe_phv_out_data_128; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_129 = pipe1_io_pipe_phv_out_data_129; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_130 = pipe1_io_pipe_phv_out_data_130; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_131 = pipe1_io_pipe_phv_out_data_131; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_132 = pipe1_io_pipe_phv_out_data_132; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_133 = pipe1_io_pipe_phv_out_data_133; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_134 = pipe1_io_pipe_phv_out_data_134; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_135 = pipe1_io_pipe_phv_out_data_135; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_136 = pipe1_io_pipe_phv_out_data_136; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_137 = pipe1_io_pipe_phv_out_data_137; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_138 = pipe1_io_pipe_phv_out_data_138; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_139 = pipe1_io_pipe_phv_out_data_139; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_140 = pipe1_io_pipe_phv_out_data_140; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_141 = pipe1_io_pipe_phv_out_data_141; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_142 = pipe1_io_pipe_phv_out_data_142; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_143 = pipe1_io_pipe_phv_out_data_143; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_144 = pipe1_io_pipe_phv_out_data_144; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_145 = pipe1_io_pipe_phv_out_data_145; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_146 = pipe1_io_pipe_phv_out_data_146; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_147 = pipe1_io_pipe_phv_out_data_147; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_148 = pipe1_io_pipe_phv_out_data_148; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_149 = pipe1_io_pipe_phv_out_data_149; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_150 = pipe1_io_pipe_phv_out_data_150; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_151 = pipe1_io_pipe_phv_out_data_151; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_152 = pipe1_io_pipe_phv_out_data_152; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_153 = pipe1_io_pipe_phv_out_data_153; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_154 = pipe1_io_pipe_phv_out_data_154; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_155 = pipe1_io_pipe_phv_out_data_155; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_156 = pipe1_io_pipe_phv_out_data_156; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_157 = pipe1_io_pipe_phv_out_data_157; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_158 = pipe1_io_pipe_phv_out_data_158; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_159 = pipe1_io_pipe_phv_out_data_159; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_160 = pipe1_io_pipe_phv_out_data_160; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_161 = pipe1_io_pipe_phv_out_data_161; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_162 = pipe1_io_pipe_phv_out_data_162; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_163 = pipe1_io_pipe_phv_out_data_163; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_164 = pipe1_io_pipe_phv_out_data_164; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_165 = pipe1_io_pipe_phv_out_data_165; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_166 = pipe1_io_pipe_phv_out_data_166; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_167 = pipe1_io_pipe_phv_out_data_167; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_168 = pipe1_io_pipe_phv_out_data_168; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_169 = pipe1_io_pipe_phv_out_data_169; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_170 = pipe1_io_pipe_phv_out_data_170; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_171 = pipe1_io_pipe_phv_out_data_171; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_172 = pipe1_io_pipe_phv_out_data_172; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_173 = pipe1_io_pipe_phv_out_data_173; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_174 = pipe1_io_pipe_phv_out_data_174; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_175 = pipe1_io_pipe_phv_out_data_175; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_176 = pipe1_io_pipe_phv_out_data_176; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_177 = pipe1_io_pipe_phv_out_data_177; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_178 = pipe1_io_pipe_phv_out_data_178; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_179 = pipe1_io_pipe_phv_out_data_179; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_180 = pipe1_io_pipe_phv_out_data_180; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_181 = pipe1_io_pipe_phv_out_data_181; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_182 = pipe1_io_pipe_phv_out_data_182; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_183 = pipe1_io_pipe_phv_out_data_183; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_184 = pipe1_io_pipe_phv_out_data_184; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_185 = pipe1_io_pipe_phv_out_data_185; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_186 = pipe1_io_pipe_phv_out_data_186; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_187 = pipe1_io_pipe_phv_out_data_187; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_188 = pipe1_io_pipe_phv_out_data_188; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_189 = pipe1_io_pipe_phv_out_data_189; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_190 = pipe1_io_pipe_phv_out_data_190; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_191 = pipe1_io_pipe_phv_out_data_191; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_192 = pipe1_io_pipe_phv_out_data_192; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_193 = pipe1_io_pipe_phv_out_data_193; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_194 = pipe1_io_pipe_phv_out_data_194; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_195 = pipe1_io_pipe_phv_out_data_195; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_196 = pipe1_io_pipe_phv_out_data_196; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_197 = pipe1_io_pipe_phv_out_data_197; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_198 = pipe1_io_pipe_phv_out_data_198; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_199 = pipe1_io_pipe_phv_out_data_199; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_200 = pipe1_io_pipe_phv_out_data_200; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_201 = pipe1_io_pipe_phv_out_data_201; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_202 = pipe1_io_pipe_phv_out_data_202; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_203 = pipe1_io_pipe_phv_out_data_203; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_204 = pipe1_io_pipe_phv_out_data_204; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_205 = pipe1_io_pipe_phv_out_data_205; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_206 = pipe1_io_pipe_phv_out_data_206; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_207 = pipe1_io_pipe_phv_out_data_207; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_208 = pipe1_io_pipe_phv_out_data_208; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_209 = pipe1_io_pipe_phv_out_data_209; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_210 = pipe1_io_pipe_phv_out_data_210; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_211 = pipe1_io_pipe_phv_out_data_211; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_212 = pipe1_io_pipe_phv_out_data_212; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_213 = pipe1_io_pipe_phv_out_data_213; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_214 = pipe1_io_pipe_phv_out_data_214; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_215 = pipe1_io_pipe_phv_out_data_215; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_216 = pipe1_io_pipe_phv_out_data_216; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_217 = pipe1_io_pipe_phv_out_data_217; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_218 = pipe1_io_pipe_phv_out_data_218; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_219 = pipe1_io_pipe_phv_out_data_219; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_220 = pipe1_io_pipe_phv_out_data_220; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_221 = pipe1_io_pipe_phv_out_data_221; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_222 = pipe1_io_pipe_phv_out_data_222; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_223 = pipe1_io_pipe_phv_out_data_223; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_224 = pipe1_io_pipe_phv_out_data_224; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_225 = pipe1_io_pipe_phv_out_data_225; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_226 = pipe1_io_pipe_phv_out_data_226; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_227 = pipe1_io_pipe_phv_out_data_227; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_228 = pipe1_io_pipe_phv_out_data_228; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_229 = pipe1_io_pipe_phv_out_data_229; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_230 = pipe1_io_pipe_phv_out_data_230; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_231 = pipe1_io_pipe_phv_out_data_231; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_232 = pipe1_io_pipe_phv_out_data_232; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_233 = pipe1_io_pipe_phv_out_data_233; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_234 = pipe1_io_pipe_phv_out_data_234; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_235 = pipe1_io_pipe_phv_out_data_235; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_236 = pipe1_io_pipe_phv_out_data_236; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_237 = pipe1_io_pipe_phv_out_data_237; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_238 = pipe1_io_pipe_phv_out_data_238; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_239 = pipe1_io_pipe_phv_out_data_239; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_240 = pipe1_io_pipe_phv_out_data_240; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_241 = pipe1_io_pipe_phv_out_data_241; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_242 = pipe1_io_pipe_phv_out_data_242; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_243 = pipe1_io_pipe_phv_out_data_243; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_244 = pipe1_io_pipe_phv_out_data_244; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_245 = pipe1_io_pipe_phv_out_data_245; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_246 = pipe1_io_pipe_phv_out_data_246; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_247 = pipe1_io_pipe_phv_out_data_247; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_248 = pipe1_io_pipe_phv_out_data_248; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_249 = pipe1_io_pipe_phv_out_data_249; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_250 = pipe1_io_pipe_phv_out_data_250; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_251 = pipe1_io_pipe_phv_out_data_251; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_252 = pipe1_io_pipe_phv_out_data_252; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_253 = pipe1_io_pipe_phv_out_data_253; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_254 = pipe1_io_pipe_phv_out_data_254; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_255 = pipe1_io_pipe_phv_out_data_255; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_256 = pipe1_io_pipe_phv_out_data_256; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_257 = pipe1_io_pipe_phv_out_data_257; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_258 = pipe1_io_pipe_phv_out_data_258; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_259 = pipe1_io_pipe_phv_out_data_259; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_260 = pipe1_io_pipe_phv_out_data_260; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_261 = pipe1_io_pipe_phv_out_data_261; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_262 = pipe1_io_pipe_phv_out_data_262; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_263 = pipe1_io_pipe_phv_out_data_263; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_264 = pipe1_io_pipe_phv_out_data_264; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_265 = pipe1_io_pipe_phv_out_data_265; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_266 = pipe1_io_pipe_phv_out_data_266; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_267 = pipe1_io_pipe_phv_out_data_267; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_268 = pipe1_io_pipe_phv_out_data_268; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_269 = pipe1_io_pipe_phv_out_data_269; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_270 = pipe1_io_pipe_phv_out_data_270; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_271 = pipe1_io_pipe_phv_out_data_271; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_272 = pipe1_io_pipe_phv_out_data_272; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_273 = pipe1_io_pipe_phv_out_data_273; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_274 = pipe1_io_pipe_phv_out_data_274; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_275 = pipe1_io_pipe_phv_out_data_275; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_276 = pipe1_io_pipe_phv_out_data_276; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_277 = pipe1_io_pipe_phv_out_data_277; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_278 = pipe1_io_pipe_phv_out_data_278; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_279 = pipe1_io_pipe_phv_out_data_279; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_280 = pipe1_io_pipe_phv_out_data_280; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_281 = pipe1_io_pipe_phv_out_data_281; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_282 = pipe1_io_pipe_phv_out_data_282; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_283 = pipe1_io_pipe_phv_out_data_283; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_284 = pipe1_io_pipe_phv_out_data_284; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_285 = pipe1_io_pipe_phv_out_data_285; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_286 = pipe1_io_pipe_phv_out_data_286; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_287 = pipe1_io_pipe_phv_out_data_287; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_288 = pipe1_io_pipe_phv_out_data_288; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_289 = pipe1_io_pipe_phv_out_data_289; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_290 = pipe1_io_pipe_phv_out_data_290; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_291 = pipe1_io_pipe_phv_out_data_291; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_292 = pipe1_io_pipe_phv_out_data_292; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_293 = pipe1_io_pipe_phv_out_data_293; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_294 = pipe1_io_pipe_phv_out_data_294; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_295 = pipe1_io_pipe_phv_out_data_295; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_296 = pipe1_io_pipe_phv_out_data_296; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_297 = pipe1_io_pipe_phv_out_data_297; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_298 = pipe1_io_pipe_phv_out_data_298; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_299 = pipe1_io_pipe_phv_out_data_299; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_300 = pipe1_io_pipe_phv_out_data_300; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_301 = pipe1_io_pipe_phv_out_data_301; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_302 = pipe1_io_pipe_phv_out_data_302; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_303 = pipe1_io_pipe_phv_out_data_303; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_304 = pipe1_io_pipe_phv_out_data_304; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_305 = pipe1_io_pipe_phv_out_data_305; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_306 = pipe1_io_pipe_phv_out_data_306; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_307 = pipe1_io_pipe_phv_out_data_307; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_308 = pipe1_io_pipe_phv_out_data_308; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_309 = pipe1_io_pipe_phv_out_data_309; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_310 = pipe1_io_pipe_phv_out_data_310; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_311 = pipe1_io_pipe_phv_out_data_311; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_312 = pipe1_io_pipe_phv_out_data_312; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_313 = pipe1_io_pipe_phv_out_data_313; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_314 = pipe1_io_pipe_phv_out_data_314; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_315 = pipe1_io_pipe_phv_out_data_315; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_316 = pipe1_io_pipe_phv_out_data_316; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_317 = pipe1_io_pipe_phv_out_data_317; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_318 = pipe1_io_pipe_phv_out_data_318; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_319 = pipe1_io_pipe_phv_out_data_319; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_320 = pipe1_io_pipe_phv_out_data_320; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_321 = pipe1_io_pipe_phv_out_data_321; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_322 = pipe1_io_pipe_phv_out_data_322; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_323 = pipe1_io_pipe_phv_out_data_323; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_324 = pipe1_io_pipe_phv_out_data_324; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_325 = pipe1_io_pipe_phv_out_data_325; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_326 = pipe1_io_pipe_phv_out_data_326; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_327 = pipe1_io_pipe_phv_out_data_327; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_328 = pipe1_io_pipe_phv_out_data_328; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_329 = pipe1_io_pipe_phv_out_data_329; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_330 = pipe1_io_pipe_phv_out_data_330; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_331 = pipe1_io_pipe_phv_out_data_331; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_332 = pipe1_io_pipe_phv_out_data_332; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_333 = pipe1_io_pipe_phv_out_data_333; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_334 = pipe1_io_pipe_phv_out_data_334; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_335 = pipe1_io_pipe_phv_out_data_335; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_336 = pipe1_io_pipe_phv_out_data_336; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_337 = pipe1_io_pipe_phv_out_data_337; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_338 = pipe1_io_pipe_phv_out_data_338; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_339 = pipe1_io_pipe_phv_out_data_339; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_340 = pipe1_io_pipe_phv_out_data_340; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_341 = pipe1_io_pipe_phv_out_data_341; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_342 = pipe1_io_pipe_phv_out_data_342; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_343 = pipe1_io_pipe_phv_out_data_343; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_344 = pipe1_io_pipe_phv_out_data_344; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_345 = pipe1_io_pipe_phv_out_data_345; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_346 = pipe1_io_pipe_phv_out_data_346; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_347 = pipe1_io_pipe_phv_out_data_347; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_348 = pipe1_io_pipe_phv_out_data_348; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_349 = pipe1_io_pipe_phv_out_data_349; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_350 = pipe1_io_pipe_phv_out_data_350; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_351 = pipe1_io_pipe_phv_out_data_351; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_352 = pipe1_io_pipe_phv_out_data_352; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_353 = pipe1_io_pipe_phv_out_data_353; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_354 = pipe1_io_pipe_phv_out_data_354; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_355 = pipe1_io_pipe_phv_out_data_355; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_356 = pipe1_io_pipe_phv_out_data_356; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_357 = pipe1_io_pipe_phv_out_data_357; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_358 = pipe1_io_pipe_phv_out_data_358; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_359 = pipe1_io_pipe_phv_out_data_359; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_360 = pipe1_io_pipe_phv_out_data_360; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_361 = pipe1_io_pipe_phv_out_data_361; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_362 = pipe1_io_pipe_phv_out_data_362; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_363 = pipe1_io_pipe_phv_out_data_363; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_364 = pipe1_io_pipe_phv_out_data_364; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_365 = pipe1_io_pipe_phv_out_data_365; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_366 = pipe1_io_pipe_phv_out_data_366; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_367 = pipe1_io_pipe_phv_out_data_367; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_368 = pipe1_io_pipe_phv_out_data_368; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_369 = pipe1_io_pipe_phv_out_data_369; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_370 = pipe1_io_pipe_phv_out_data_370; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_371 = pipe1_io_pipe_phv_out_data_371; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_372 = pipe1_io_pipe_phv_out_data_372; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_373 = pipe1_io_pipe_phv_out_data_373; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_374 = pipe1_io_pipe_phv_out_data_374; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_375 = pipe1_io_pipe_phv_out_data_375; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_376 = pipe1_io_pipe_phv_out_data_376; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_377 = pipe1_io_pipe_phv_out_data_377; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_378 = pipe1_io_pipe_phv_out_data_378; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_379 = pipe1_io_pipe_phv_out_data_379; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_380 = pipe1_io_pipe_phv_out_data_380; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_381 = pipe1_io_pipe_phv_out_data_381; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_382 = pipe1_io_pipe_phv_out_data_382; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_383 = pipe1_io_pipe_phv_out_data_383; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_384 = pipe1_io_pipe_phv_out_data_384; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_385 = pipe1_io_pipe_phv_out_data_385; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_386 = pipe1_io_pipe_phv_out_data_386; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_387 = pipe1_io_pipe_phv_out_data_387; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_388 = pipe1_io_pipe_phv_out_data_388; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_389 = pipe1_io_pipe_phv_out_data_389; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_390 = pipe1_io_pipe_phv_out_data_390; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_391 = pipe1_io_pipe_phv_out_data_391; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_392 = pipe1_io_pipe_phv_out_data_392; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_393 = pipe1_io_pipe_phv_out_data_393; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_394 = pipe1_io_pipe_phv_out_data_394; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_395 = pipe1_io_pipe_phv_out_data_395; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_396 = pipe1_io_pipe_phv_out_data_396; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_397 = pipe1_io_pipe_phv_out_data_397; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_398 = pipe1_io_pipe_phv_out_data_398; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_399 = pipe1_io_pipe_phv_out_data_399; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_400 = pipe1_io_pipe_phv_out_data_400; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_401 = pipe1_io_pipe_phv_out_data_401; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_402 = pipe1_io_pipe_phv_out_data_402; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_403 = pipe1_io_pipe_phv_out_data_403; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_404 = pipe1_io_pipe_phv_out_data_404; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_405 = pipe1_io_pipe_phv_out_data_405; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_406 = pipe1_io_pipe_phv_out_data_406; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_407 = pipe1_io_pipe_phv_out_data_407; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_408 = pipe1_io_pipe_phv_out_data_408; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_409 = pipe1_io_pipe_phv_out_data_409; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_410 = pipe1_io_pipe_phv_out_data_410; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_411 = pipe1_io_pipe_phv_out_data_411; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_412 = pipe1_io_pipe_phv_out_data_412; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_413 = pipe1_io_pipe_phv_out_data_413; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_414 = pipe1_io_pipe_phv_out_data_414; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_415 = pipe1_io_pipe_phv_out_data_415; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_416 = pipe1_io_pipe_phv_out_data_416; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_417 = pipe1_io_pipe_phv_out_data_417; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_418 = pipe1_io_pipe_phv_out_data_418; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_419 = pipe1_io_pipe_phv_out_data_419; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_420 = pipe1_io_pipe_phv_out_data_420; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_421 = pipe1_io_pipe_phv_out_data_421; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_422 = pipe1_io_pipe_phv_out_data_422; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_423 = pipe1_io_pipe_phv_out_data_423; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_424 = pipe1_io_pipe_phv_out_data_424; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_425 = pipe1_io_pipe_phv_out_data_425; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_426 = pipe1_io_pipe_phv_out_data_426; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_427 = pipe1_io_pipe_phv_out_data_427; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_428 = pipe1_io_pipe_phv_out_data_428; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_429 = pipe1_io_pipe_phv_out_data_429; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_430 = pipe1_io_pipe_phv_out_data_430; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_431 = pipe1_io_pipe_phv_out_data_431; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_432 = pipe1_io_pipe_phv_out_data_432; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_433 = pipe1_io_pipe_phv_out_data_433; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_434 = pipe1_io_pipe_phv_out_data_434; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_435 = pipe1_io_pipe_phv_out_data_435; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_436 = pipe1_io_pipe_phv_out_data_436; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_437 = pipe1_io_pipe_phv_out_data_437; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_438 = pipe1_io_pipe_phv_out_data_438; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_439 = pipe1_io_pipe_phv_out_data_439; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_440 = pipe1_io_pipe_phv_out_data_440; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_441 = pipe1_io_pipe_phv_out_data_441; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_442 = pipe1_io_pipe_phv_out_data_442; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_443 = pipe1_io_pipe_phv_out_data_443; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_444 = pipe1_io_pipe_phv_out_data_444; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_445 = pipe1_io_pipe_phv_out_data_445; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_446 = pipe1_io_pipe_phv_out_data_446; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_447 = pipe1_io_pipe_phv_out_data_447; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_448 = pipe1_io_pipe_phv_out_data_448; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_449 = pipe1_io_pipe_phv_out_data_449; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_450 = pipe1_io_pipe_phv_out_data_450; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_451 = pipe1_io_pipe_phv_out_data_451; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_452 = pipe1_io_pipe_phv_out_data_452; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_453 = pipe1_io_pipe_phv_out_data_453; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_454 = pipe1_io_pipe_phv_out_data_454; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_455 = pipe1_io_pipe_phv_out_data_455; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_456 = pipe1_io_pipe_phv_out_data_456; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_457 = pipe1_io_pipe_phv_out_data_457; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_458 = pipe1_io_pipe_phv_out_data_458; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_459 = pipe1_io_pipe_phv_out_data_459; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_460 = pipe1_io_pipe_phv_out_data_460; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_461 = pipe1_io_pipe_phv_out_data_461; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_462 = pipe1_io_pipe_phv_out_data_462; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_463 = pipe1_io_pipe_phv_out_data_463; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_464 = pipe1_io_pipe_phv_out_data_464; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_465 = pipe1_io_pipe_phv_out_data_465; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_466 = pipe1_io_pipe_phv_out_data_466; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_467 = pipe1_io_pipe_phv_out_data_467; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_468 = pipe1_io_pipe_phv_out_data_468; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_469 = pipe1_io_pipe_phv_out_data_469; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_470 = pipe1_io_pipe_phv_out_data_470; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_471 = pipe1_io_pipe_phv_out_data_471; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_472 = pipe1_io_pipe_phv_out_data_472; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_473 = pipe1_io_pipe_phv_out_data_473; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_474 = pipe1_io_pipe_phv_out_data_474; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_475 = pipe1_io_pipe_phv_out_data_475; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_476 = pipe1_io_pipe_phv_out_data_476; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_477 = pipe1_io_pipe_phv_out_data_477; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_478 = pipe1_io_pipe_phv_out_data_478; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_479 = pipe1_io_pipe_phv_out_data_479; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_480 = pipe1_io_pipe_phv_out_data_480; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_481 = pipe1_io_pipe_phv_out_data_481; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_482 = pipe1_io_pipe_phv_out_data_482; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_483 = pipe1_io_pipe_phv_out_data_483; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_484 = pipe1_io_pipe_phv_out_data_484; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_485 = pipe1_io_pipe_phv_out_data_485; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_486 = pipe1_io_pipe_phv_out_data_486; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_487 = pipe1_io_pipe_phv_out_data_487; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_488 = pipe1_io_pipe_phv_out_data_488; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_489 = pipe1_io_pipe_phv_out_data_489; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_490 = pipe1_io_pipe_phv_out_data_490; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_491 = pipe1_io_pipe_phv_out_data_491; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_492 = pipe1_io_pipe_phv_out_data_492; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_493 = pipe1_io_pipe_phv_out_data_493; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_494 = pipe1_io_pipe_phv_out_data_494; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_495 = pipe1_io_pipe_phv_out_data_495; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_496 = pipe1_io_pipe_phv_out_data_496; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_497 = pipe1_io_pipe_phv_out_data_497; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_498 = pipe1_io_pipe_phv_out_data_498; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_499 = pipe1_io_pipe_phv_out_data_499; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_500 = pipe1_io_pipe_phv_out_data_500; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_501 = pipe1_io_pipe_phv_out_data_501; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_502 = pipe1_io_pipe_phv_out_data_502; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_503 = pipe1_io_pipe_phv_out_data_503; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_504 = pipe1_io_pipe_phv_out_data_504; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_505 = pipe1_io_pipe_phv_out_data_505; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_506 = pipe1_io_pipe_phv_out_data_506; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_507 = pipe1_io_pipe_phv_out_data_507; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_508 = pipe1_io_pipe_phv_out_data_508; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_509 = pipe1_io_pipe_phv_out_data_509; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_510 = pipe1_io_pipe_phv_out_data_510; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_511 = pipe1_io_pipe_phv_out_data_511; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_0 = pipe1_io_pipe_phv_out_header_0; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_1 = pipe1_io_pipe_phv_out_header_1; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_2 = pipe1_io_pipe_phv_out_header_2; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_3 = pipe1_io_pipe_phv_out_header_3; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_4 = pipe1_io_pipe_phv_out_header_4; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_5 = pipe1_io_pipe_phv_out_header_5; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_6 = pipe1_io_pipe_phv_out_header_6; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_7 = pipe1_io_pipe_phv_out_header_7; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_8 = pipe1_io_pipe_phv_out_header_8; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_9 = pipe1_io_pipe_phv_out_header_9; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_10 = pipe1_io_pipe_phv_out_header_10; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_11 = pipe1_io_pipe_phv_out_header_11; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_12 = pipe1_io_pipe_phv_out_header_12; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_13 = pipe1_io_pipe_phv_out_header_13; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_14 = pipe1_io_pipe_phv_out_header_14; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_15 = pipe1_io_pipe_phv_out_header_15; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_parse_current_state = pipe1_io_pipe_phv_out_parse_current_state; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_parse_current_offset = pipe1_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_parse_transition_field = pipe1_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_next_processor_id = pipe1_io_pipe_phv_out_next_processor_id; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_next_config_id = pipe1_io_pipe_phv_out_next_config_id; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_is_valid_processor = pipe1_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 354:26]
  assign pipe2_io_key_config_0_key_length = key_config_0_key_length; // @[matcher.scala 356:26]
  assign pipe2_io_key_config_1_key_length = key_config_1_key_length; // @[matcher.scala 356:26]
  assign pipe2_io_key_offset = pipe1_io_key_offset; // @[matcher.scala 355:26]
  assign pipe3to8_clock = clock;
  assign pipe3to8_io_pipe_phv_in_data_0 = pipe2_io_pipe_phv_out_data_0; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_1 = pipe2_io_pipe_phv_out_data_1; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_2 = pipe2_io_pipe_phv_out_data_2; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_3 = pipe2_io_pipe_phv_out_data_3; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_4 = pipe2_io_pipe_phv_out_data_4; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_5 = pipe2_io_pipe_phv_out_data_5; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_6 = pipe2_io_pipe_phv_out_data_6; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_7 = pipe2_io_pipe_phv_out_data_7; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_8 = pipe2_io_pipe_phv_out_data_8; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_9 = pipe2_io_pipe_phv_out_data_9; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_10 = pipe2_io_pipe_phv_out_data_10; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_11 = pipe2_io_pipe_phv_out_data_11; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_12 = pipe2_io_pipe_phv_out_data_12; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_13 = pipe2_io_pipe_phv_out_data_13; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_14 = pipe2_io_pipe_phv_out_data_14; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_15 = pipe2_io_pipe_phv_out_data_15; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_16 = pipe2_io_pipe_phv_out_data_16; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_17 = pipe2_io_pipe_phv_out_data_17; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_18 = pipe2_io_pipe_phv_out_data_18; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_19 = pipe2_io_pipe_phv_out_data_19; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_20 = pipe2_io_pipe_phv_out_data_20; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_21 = pipe2_io_pipe_phv_out_data_21; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_22 = pipe2_io_pipe_phv_out_data_22; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_23 = pipe2_io_pipe_phv_out_data_23; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_24 = pipe2_io_pipe_phv_out_data_24; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_25 = pipe2_io_pipe_phv_out_data_25; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_26 = pipe2_io_pipe_phv_out_data_26; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_27 = pipe2_io_pipe_phv_out_data_27; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_28 = pipe2_io_pipe_phv_out_data_28; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_29 = pipe2_io_pipe_phv_out_data_29; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_30 = pipe2_io_pipe_phv_out_data_30; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_31 = pipe2_io_pipe_phv_out_data_31; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_32 = pipe2_io_pipe_phv_out_data_32; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_33 = pipe2_io_pipe_phv_out_data_33; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_34 = pipe2_io_pipe_phv_out_data_34; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_35 = pipe2_io_pipe_phv_out_data_35; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_36 = pipe2_io_pipe_phv_out_data_36; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_37 = pipe2_io_pipe_phv_out_data_37; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_38 = pipe2_io_pipe_phv_out_data_38; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_39 = pipe2_io_pipe_phv_out_data_39; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_40 = pipe2_io_pipe_phv_out_data_40; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_41 = pipe2_io_pipe_phv_out_data_41; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_42 = pipe2_io_pipe_phv_out_data_42; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_43 = pipe2_io_pipe_phv_out_data_43; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_44 = pipe2_io_pipe_phv_out_data_44; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_45 = pipe2_io_pipe_phv_out_data_45; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_46 = pipe2_io_pipe_phv_out_data_46; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_47 = pipe2_io_pipe_phv_out_data_47; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_48 = pipe2_io_pipe_phv_out_data_48; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_49 = pipe2_io_pipe_phv_out_data_49; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_50 = pipe2_io_pipe_phv_out_data_50; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_51 = pipe2_io_pipe_phv_out_data_51; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_52 = pipe2_io_pipe_phv_out_data_52; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_53 = pipe2_io_pipe_phv_out_data_53; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_54 = pipe2_io_pipe_phv_out_data_54; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_55 = pipe2_io_pipe_phv_out_data_55; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_56 = pipe2_io_pipe_phv_out_data_56; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_57 = pipe2_io_pipe_phv_out_data_57; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_58 = pipe2_io_pipe_phv_out_data_58; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_59 = pipe2_io_pipe_phv_out_data_59; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_60 = pipe2_io_pipe_phv_out_data_60; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_61 = pipe2_io_pipe_phv_out_data_61; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_62 = pipe2_io_pipe_phv_out_data_62; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_63 = pipe2_io_pipe_phv_out_data_63; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_64 = pipe2_io_pipe_phv_out_data_64; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_65 = pipe2_io_pipe_phv_out_data_65; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_66 = pipe2_io_pipe_phv_out_data_66; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_67 = pipe2_io_pipe_phv_out_data_67; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_68 = pipe2_io_pipe_phv_out_data_68; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_69 = pipe2_io_pipe_phv_out_data_69; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_70 = pipe2_io_pipe_phv_out_data_70; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_71 = pipe2_io_pipe_phv_out_data_71; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_72 = pipe2_io_pipe_phv_out_data_72; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_73 = pipe2_io_pipe_phv_out_data_73; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_74 = pipe2_io_pipe_phv_out_data_74; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_75 = pipe2_io_pipe_phv_out_data_75; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_76 = pipe2_io_pipe_phv_out_data_76; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_77 = pipe2_io_pipe_phv_out_data_77; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_78 = pipe2_io_pipe_phv_out_data_78; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_79 = pipe2_io_pipe_phv_out_data_79; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_80 = pipe2_io_pipe_phv_out_data_80; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_81 = pipe2_io_pipe_phv_out_data_81; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_82 = pipe2_io_pipe_phv_out_data_82; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_83 = pipe2_io_pipe_phv_out_data_83; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_84 = pipe2_io_pipe_phv_out_data_84; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_85 = pipe2_io_pipe_phv_out_data_85; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_86 = pipe2_io_pipe_phv_out_data_86; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_87 = pipe2_io_pipe_phv_out_data_87; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_88 = pipe2_io_pipe_phv_out_data_88; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_89 = pipe2_io_pipe_phv_out_data_89; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_90 = pipe2_io_pipe_phv_out_data_90; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_91 = pipe2_io_pipe_phv_out_data_91; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_92 = pipe2_io_pipe_phv_out_data_92; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_93 = pipe2_io_pipe_phv_out_data_93; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_94 = pipe2_io_pipe_phv_out_data_94; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_95 = pipe2_io_pipe_phv_out_data_95; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_96 = pipe2_io_pipe_phv_out_data_96; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_97 = pipe2_io_pipe_phv_out_data_97; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_98 = pipe2_io_pipe_phv_out_data_98; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_99 = pipe2_io_pipe_phv_out_data_99; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_100 = pipe2_io_pipe_phv_out_data_100; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_101 = pipe2_io_pipe_phv_out_data_101; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_102 = pipe2_io_pipe_phv_out_data_102; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_103 = pipe2_io_pipe_phv_out_data_103; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_104 = pipe2_io_pipe_phv_out_data_104; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_105 = pipe2_io_pipe_phv_out_data_105; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_106 = pipe2_io_pipe_phv_out_data_106; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_107 = pipe2_io_pipe_phv_out_data_107; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_108 = pipe2_io_pipe_phv_out_data_108; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_109 = pipe2_io_pipe_phv_out_data_109; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_110 = pipe2_io_pipe_phv_out_data_110; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_111 = pipe2_io_pipe_phv_out_data_111; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_112 = pipe2_io_pipe_phv_out_data_112; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_113 = pipe2_io_pipe_phv_out_data_113; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_114 = pipe2_io_pipe_phv_out_data_114; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_115 = pipe2_io_pipe_phv_out_data_115; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_116 = pipe2_io_pipe_phv_out_data_116; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_117 = pipe2_io_pipe_phv_out_data_117; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_118 = pipe2_io_pipe_phv_out_data_118; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_119 = pipe2_io_pipe_phv_out_data_119; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_120 = pipe2_io_pipe_phv_out_data_120; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_121 = pipe2_io_pipe_phv_out_data_121; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_122 = pipe2_io_pipe_phv_out_data_122; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_123 = pipe2_io_pipe_phv_out_data_123; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_124 = pipe2_io_pipe_phv_out_data_124; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_125 = pipe2_io_pipe_phv_out_data_125; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_126 = pipe2_io_pipe_phv_out_data_126; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_127 = pipe2_io_pipe_phv_out_data_127; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_128 = pipe2_io_pipe_phv_out_data_128; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_129 = pipe2_io_pipe_phv_out_data_129; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_130 = pipe2_io_pipe_phv_out_data_130; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_131 = pipe2_io_pipe_phv_out_data_131; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_132 = pipe2_io_pipe_phv_out_data_132; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_133 = pipe2_io_pipe_phv_out_data_133; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_134 = pipe2_io_pipe_phv_out_data_134; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_135 = pipe2_io_pipe_phv_out_data_135; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_136 = pipe2_io_pipe_phv_out_data_136; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_137 = pipe2_io_pipe_phv_out_data_137; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_138 = pipe2_io_pipe_phv_out_data_138; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_139 = pipe2_io_pipe_phv_out_data_139; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_140 = pipe2_io_pipe_phv_out_data_140; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_141 = pipe2_io_pipe_phv_out_data_141; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_142 = pipe2_io_pipe_phv_out_data_142; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_143 = pipe2_io_pipe_phv_out_data_143; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_144 = pipe2_io_pipe_phv_out_data_144; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_145 = pipe2_io_pipe_phv_out_data_145; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_146 = pipe2_io_pipe_phv_out_data_146; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_147 = pipe2_io_pipe_phv_out_data_147; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_148 = pipe2_io_pipe_phv_out_data_148; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_149 = pipe2_io_pipe_phv_out_data_149; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_150 = pipe2_io_pipe_phv_out_data_150; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_151 = pipe2_io_pipe_phv_out_data_151; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_152 = pipe2_io_pipe_phv_out_data_152; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_153 = pipe2_io_pipe_phv_out_data_153; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_154 = pipe2_io_pipe_phv_out_data_154; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_155 = pipe2_io_pipe_phv_out_data_155; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_156 = pipe2_io_pipe_phv_out_data_156; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_157 = pipe2_io_pipe_phv_out_data_157; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_158 = pipe2_io_pipe_phv_out_data_158; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_159 = pipe2_io_pipe_phv_out_data_159; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_160 = pipe2_io_pipe_phv_out_data_160; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_161 = pipe2_io_pipe_phv_out_data_161; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_162 = pipe2_io_pipe_phv_out_data_162; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_163 = pipe2_io_pipe_phv_out_data_163; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_164 = pipe2_io_pipe_phv_out_data_164; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_165 = pipe2_io_pipe_phv_out_data_165; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_166 = pipe2_io_pipe_phv_out_data_166; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_167 = pipe2_io_pipe_phv_out_data_167; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_168 = pipe2_io_pipe_phv_out_data_168; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_169 = pipe2_io_pipe_phv_out_data_169; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_170 = pipe2_io_pipe_phv_out_data_170; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_171 = pipe2_io_pipe_phv_out_data_171; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_172 = pipe2_io_pipe_phv_out_data_172; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_173 = pipe2_io_pipe_phv_out_data_173; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_174 = pipe2_io_pipe_phv_out_data_174; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_175 = pipe2_io_pipe_phv_out_data_175; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_176 = pipe2_io_pipe_phv_out_data_176; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_177 = pipe2_io_pipe_phv_out_data_177; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_178 = pipe2_io_pipe_phv_out_data_178; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_179 = pipe2_io_pipe_phv_out_data_179; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_180 = pipe2_io_pipe_phv_out_data_180; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_181 = pipe2_io_pipe_phv_out_data_181; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_182 = pipe2_io_pipe_phv_out_data_182; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_183 = pipe2_io_pipe_phv_out_data_183; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_184 = pipe2_io_pipe_phv_out_data_184; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_185 = pipe2_io_pipe_phv_out_data_185; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_186 = pipe2_io_pipe_phv_out_data_186; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_187 = pipe2_io_pipe_phv_out_data_187; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_188 = pipe2_io_pipe_phv_out_data_188; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_189 = pipe2_io_pipe_phv_out_data_189; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_190 = pipe2_io_pipe_phv_out_data_190; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_191 = pipe2_io_pipe_phv_out_data_191; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_192 = pipe2_io_pipe_phv_out_data_192; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_193 = pipe2_io_pipe_phv_out_data_193; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_194 = pipe2_io_pipe_phv_out_data_194; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_195 = pipe2_io_pipe_phv_out_data_195; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_196 = pipe2_io_pipe_phv_out_data_196; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_197 = pipe2_io_pipe_phv_out_data_197; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_198 = pipe2_io_pipe_phv_out_data_198; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_199 = pipe2_io_pipe_phv_out_data_199; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_200 = pipe2_io_pipe_phv_out_data_200; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_201 = pipe2_io_pipe_phv_out_data_201; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_202 = pipe2_io_pipe_phv_out_data_202; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_203 = pipe2_io_pipe_phv_out_data_203; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_204 = pipe2_io_pipe_phv_out_data_204; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_205 = pipe2_io_pipe_phv_out_data_205; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_206 = pipe2_io_pipe_phv_out_data_206; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_207 = pipe2_io_pipe_phv_out_data_207; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_208 = pipe2_io_pipe_phv_out_data_208; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_209 = pipe2_io_pipe_phv_out_data_209; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_210 = pipe2_io_pipe_phv_out_data_210; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_211 = pipe2_io_pipe_phv_out_data_211; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_212 = pipe2_io_pipe_phv_out_data_212; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_213 = pipe2_io_pipe_phv_out_data_213; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_214 = pipe2_io_pipe_phv_out_data_214; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_215 = pipe2_io_pipe_phv_out_data_215; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_216 = pipe2_io_pipe_phv_out_data_216; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_217 = pipe2_io_pipe_phv_out_data_217; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_218 = pipe2_io_pipe_phv_out_data_218; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_219 = pipe2_io_pipe_phv_out_data_219; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_220 = pipe2_io_pipe_phv_out_data_220; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_221 = pipe2_io_pipe_phv_out_data_221; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_222 = pipe2_io_pipe_phv_out_data_222; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_223 = pipe2_io_pipe_phv_out_data_223; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_224 = pipe2_io_pipe_phv_out_data_224; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_225 = pipe2_io_pipe_phv_out_data_225; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_226 = pipe2_io_pipe_phv_out_data_226; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_227 = pipe2_io_pipe_phv_out_data_227; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_228 = pipe2_io_pipe_phv_out_data_228; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_229 = pipe2_io_pipe_phv_out_data_229; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_230 = pipe2_io_pipe_phv_out_data_230; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_231 = pipe2_io_pipe_phv_out_data_231; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_232 = pipe2_io_pipe_phv_out_data_232; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_233 = pipe2_io_pipe_phv_out_data_233; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_234 = pipe2_io_pipe_phv_out_data_234; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_235 = pipe2_io_pipe_phv_out_data_235; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_236 = pipe2_io_pipe_phv_out_data_236; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_237 = pipe2_io_pipe_phv_out_data_237; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_238 = pipe2_io_pipe_phv_out_data_238; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_239 = pipe2_io_pipe_phv_out_data_239; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_240 = pipe2_io_pipe_phv_out_data_240; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_241 = pipe2_io_pipe_phv_out_data_241; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_242 = pipe2_io_pipe_phv_out_data_242; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_243 = pipe2_io_pipe_phv_out_data_243; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_244 = pipe2_io_pipe_phv_out_data_244; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_245 = pipe2_io_pipe_phv_out_data_245; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_246 = pipe2_io_pipe_phv_out_data_246; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_247 = pipe2_io_pipe_phv_out_data_247; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_248 = pipe2_io_pipe_phv_out_data_248; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_249 = pipe2_io_pipe_phv_out_data_249; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_250 = pipe2_io_pipe_phv_out_data_250; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_251 = pipe2_io_pipe_phv_out_data_251; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_252 = pipe2_io_pipe_phv_out_data_252; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_253 = pipe2_io_pipe_phv_out_data_253; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_254 = pipe2_io_pipe_phv_out_data_254; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_255 = pipe2_io_pipe_phv_out_data_255; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_256 = pipe2_io_pipe_phv_out_data_256; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_257 = pipe2_io_pipe_phv_out_data_257; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_258 = pipe2_io_pipe_phv_out_data_258; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_259 = pipe2_io_pipe_phv_out_data_259; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_260 = pipe2_io_pipe_phv_out_data_260; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_261 = pipe2_io_pipe_phv_out_data_261; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_262 = pipe2_io_pipe_phv_out_data_262; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_263 = pipe2_io_pipe_phv_out_data_263; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_264 = pipe2_io_pipe_phv_out_data_264; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_265 = pipe2_io_pipe_phv_out_data_265; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_266 = pipe2_io_pipe_phv_out_data_266; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_267 = pipe2_io_pipe_phv_out_data_267; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_268 = pipe2_io_pipe_phv_out_data_268; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_269 = pipe2_io_pipe_phv_out_data_269; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_270 = pipe2_io_pipe_phv_out_data_270; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_271 = pipe2_io_pipe_phv_out_data_271; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_272 = pipe2_io_pipe_phv_out_data_272; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_273 = pipe2_io_pipe_phv_out_data_273; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_274 = pipe2_io_pipe_phv_out_data_274; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_275 = pipe2_io_pipe_phv_out_data_275; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_276 = pipe2_io_pipe_phv_out_data_276; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_277 = pipe2_io_pipe_phv_out_data_277; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_278 = pipe2_io_pipe_phv_out_data_278; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_279 = pipe2_io_pipe_phv_out_data_279; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_280 = pipe2_io_pipe_phv_out_data_280; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_281 = pipe2_io_pipe_phv_out_data_281; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_282 = pipe2_io_pipe_phv_out_data_282; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_283 = pipe2_io_pipe_phv_out_data_283; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_284 = pipe2_io_pipe_phv_out_data_284; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_285 = pipe2_io_pipe_phv_out_data_285; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_286 = pipe2_io_pipe_phv_out_data_286; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_287 = pipe2_io_pipe_phv_out_data_287; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_288 = pipe2_io_pipe_phv_out_data_288; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_289 = pipe2_io_pipe_phv_out_data_289; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_290 = pipe2_io_pipe_phv_out_data_290; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_291 = pipe2_io_pipe_phv_out_data_291; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_292 = pipe2_io_pipe_phv_out_data_292; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_293 = pipe2_io_pipe_phv_out_data_293; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_294 = pipe2_io_pipe_phv_out_data_294; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_295 = pipe2_io_pipe_phv_out_data_295; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_296 = pipe2_io_pipe_phv_out_data_296; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_297 = pipe2_io_pipe_phv_out_data_297; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_298 = pipe2_io_pipe_phv_out_data_298; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_299 = pipe2_io_pipe_phv_out_data_299; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_300 = pipe2_io_pipe_phv_out_data_300; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_301 = pipe2_io_pipe_phv_out_data_301; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_302 = pipe2_io_pipe_phv_out_data_302; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_303 = pipe2_io_pipe_phv_out_data_303; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_304 = pipe2_io_pipe_phv_out_data_304; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_305 = pipe2_io_pipe_phv_out_data_305; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_306 = pipe2_io_pipe_phv_out_data_306; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_307 = pipe2_io_pipe_phv_out_data_307; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_308 = pipe2_io_pipe_phv_out_data_308; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_309 = pipe2_io_pipe_phv_out_data_309; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_310 = pipe2_io_pipe_phv_out_data_310; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_311 = pipe2_io_pipe_phv_out_data_311; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_312 = pipe2_io_pipe_phv_out_data_312; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_313 = pipe2_io_pipe_phv_out_data_313; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_314 = pipe2_io_pipe_phv_out_data_314; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_315 = pipe2_io_pipe_phv_out_data_315; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_316 = pipe2_io_pipe_phv_out_data_316; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_317 = pipe2_io_pipe_phv_out_data_317; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_318 = pipe2_io_pipe_phv_out_data_318; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_319 = pipe2_io_pipe_phv_out_data_319; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_320 = pipe2_io_pipe_phv_out_data_320; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_321 = pipe2_io_pipe_phv_out_data_321; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_322 = pipe2_io_pipe_phv_out_data_322; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_323 = pipe2_io_pipe_phv_out_data_323; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_324 = pipe2_io_pipe_phv_out_data_324; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_325 = pipe2_io_pipe_phv_out_data_325; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_326 = pipe2_io_pipe_phv_out_data_326; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_327 = pipe2_io_pipe_phv_out_data_327; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_328 = pipe2_io_pipe_phv_out_data_328; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_329 = pipe2_io_pipe_phv_out_data_329; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_330 = pipe2_io_pipe_phv_out_data_330; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_331 = pipe2_io_pipe_phv_out_data_331; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_332 = pipe2_io_pipe_phv_out_data_332; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_333 = pipe2_io_pipe_phv_out_data_333; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_334 = pipe2_io_pipe_phv_out_data_334; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_335 = pipe2_io_pipe_phv_out_data_335; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_336 = pipe2_io_pipe_phv_out_data_336; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_337 = pipe2_io_pipe_phv_out_data_337; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_338 = pipe2_io_pipe_phv_out_data_338; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_339 = pipe2_io_pipe_phv_out_data_339; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_340 = pipe2_io_pipe_phv_out_data_340; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_341 = pipe2_io_pipe_phv_out_data_341; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_342 = pipe2_io_pipe_phv_out_data_342; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_343 = pipe2_io_pipe_phv_out_data_343; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_344 = pipe2_io_pipe_phv_out_data_344; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_345 = pipe2_io_pipe_phv_out_data_345; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_346 = pipe2_io_pipe_phv_out_data_346; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_347 = pipe2_io_pipe_phv_out_data_347; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_348 = pipe2_io_pipe_phv_out_data_348; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_349 = pipe2_io_pipe_phv_out_data_349; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_350 = pipe2_io_pipe_phv_out_data_350; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_351 = pipe2_io_pipe_phv_out_data_351; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_352 = pipe2_io_pipe_phv_out_data_352; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_353 = pipe2_io_pipe_phv_out_data_353; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_354 = pipe2_io_pipe_phv_out_data_354; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_355 = pipe2_io_pipe_phv_out_data_355; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_356 = pipe2_io_pipe_phv_out_data_356; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_357 = pipe2_io_pipe_phv_out_data_357; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_358 = pipe2_io_pipe_phv_out_data_358; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_359 = pipe2_io_pipe_phv_out_data_359; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_360 = pipe2_io_pipe_phv_out_data_360; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_361 = pipe2_io_pipe_phv_out_data_361; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_362 = pipe2_io_pipe_phv_out_data_362; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_363 = pipe2_io_pipe_phv_out_data_363; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_364 = pipe2_io_pipe_phv_out_data_364; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_365 = pipe2_io_pipe_phv_out_data_365; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_366 = pipe2_io_pipe_phv_out_data_366; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_367 = pipe2_io_pipe_phv_out_data_367; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_368 = pipe2_io_pipe_phv_out_data_368; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_369 = pipe2_io_pipe_phv_out_data_369; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_370 = pipe2_io_pipe_phv_out_data_370; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_371 = pipe2_io_pipe_phv_out_data_371; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_372 = pipe2_io_pipe_phv_out_data_372; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_373 = pipe2_io_pipe_phv_out_data_373; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_374 = pipe2_io_pipe_phv_out_data_374; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_375 = pipe2_io_pipe_phv_out_data_375; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_376 = pipe2_io_pipe_phv_out_data_376; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_377 = pipe2_io_pipe_phv_out_data_377; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_378 = pipe2_io_pipe_phv_out_data_378; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_379 = pipe2_io_pipe_phv_out_data_379; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_380 = pipe2_io_pipe_phv_out_data_380; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_381 = pipe2_io_pipe_phv_out_data_381; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_382 = pipe2_io_pipe_phv_out_data_382; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_383 = pipe2_io_pipe_phv_out_data_383; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_384 = pipe2_io_pipe_phv_out_data_384; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_385 = pipe2_io_pipe_phv_out_data_385; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_386 = pipe2_io_pipe_phv_out_data_386; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_387 = pipe2_io_pipe_phv_out_data_387; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_388 = pipe2_io_pipe_phv_out_data_388; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_389 = pipe2_io_pipe_phv_out_data_389; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_390 = pipe2_io_pipe_phv_out_data_390; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_391 = pipe2_io_pipe_phv_out_data_391; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_392 = pipe2_io_pipe_phv_out_data_392; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_393 = pipe2_io_pipe_phv_out_data_393; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_394 = pipe2_io_pipe_phv_out_data_394; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_395 = pipe2_io_pipe_phv_out_data_395; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_396 = pipe2_io_pipe_phv_out_data_396; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_397 = pipe2_io_pipe_phv_out_data_397; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_398 = pipe2_io_pipe_phv_out_data_398; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_399 = pipe2_io_pipe_phv_out_data_399; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_400 = pipe2_io_pipe_phv_out_data_400; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_401 = pipe2_io_pipe_phv_out_data_401; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_402 = pipe2_io_pipe_phv_out_data_402; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_403 = pipe2_io_pipe_phv_out_data_403; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_404 = pipe2_io_pipe_phv_out_data_404; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_405 = pipe2_io_pipe_phv_out_data_405; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_406 = pipe2_io_pipe_phv_out_data_406; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_407 = pipe2_io_pipe_phv_out_data_407; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_408 = pipe2_io_pipe_phv_out_data_408; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_409 = pipe2_io_pipe_phv_out_data_409; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_410 = pipe2_io_pipe_phv_out_data_410; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_411 = pipe2_io_pipe_phv_out_data_411; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_412 = pipe2_io_pipe_phv_out_data_412; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_413 = pipe2_io_pipe_phv_out_data_413; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_414 = pipe2_io_pipe_phv_out_data_414; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_415 = pipe2_io_pipe_phv_out_data_415; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_416 = pipe2_io_pipe_phv_out_data_416; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_417 = pipe2_io_pipe_phv_out_data_417; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_418 = pipe2_io_pipe_phv_out_data_418; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_419 = pipe2_io_pipe_phv_out_data_419; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_420 = pipe2_io_pipe_phv_out_data_420; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_421 = pipe2_io_pipe_phv_out_data_421; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_422 = pipe2_io_pipe_phv_out_data_422; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_423 = pipe2_io_pipe_phv_out_data_423; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_424 = pipe2_io_pipe_phv_out_data_424; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_425 = pipe2_io_pipe_phv_out_data_425; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_426 = pipe2_io_pipe_phv_out_data_426; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_427 = pipe2_io_pipe_phv_out_data_427; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_428 = pipe2_io_pipe_phv_out_data_428; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_429 = pipe2_io_pipe_phv_out_data_429; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_430 = pipe2_io_pipe_phv_out_data_430; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_431 = pipe2_io_pipe_phv_out_data_431; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_432 = pipe2_io_pipe_phv_out_data_432; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_433 = pipe2_io_pipe_phv_out_data_433; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_434 = pipe2_io_pipe_phv_out_data_434; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_435 = pipe2_io_pipe_phv_out_data_435; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_436 = pipe2_io_pipe_phv_out_data_436; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_437 = pipe2_io_pipe_phv_out_data_437; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_438 = pipe2_io_pipe_phv_out_data_438; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_439 = pipe2_io_pipe_phv_out_data_439; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_440 = pipe2_io_pipe_phv_out_data_440; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_441 = pipe2_io_pipe_phv_out_data_441; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_442 = pipe2_io_pipe_phv_out_data_442; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_443 = pipe2_io_pipe_phv_out_data_443; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_444 = pipe2_io_pipe_phv_out_data_444; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_445 = pipe2_io_pipe_phv_out_data_445; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_446 = pipe2_io_pipe_phv_out_data_446; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_447 = pipe2_io_pipe_phv_out_data_447; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_448 = pipe2_io_pipe_phv_out_data_448; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_449 = pipe2_io_pipe_phv_out_data_449; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_450 = pipe2_io_pipe_phv_out_data_450; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_451 = pipe2_io_pipe_phv_out_data_451; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_452 = pipe2_io_pipe_phv_out_data_452; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_453 = pipe2_io_pipe_phv_out_data_453; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_454 = pipe2_io_pipe_phv_out_data_454; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_455 = pipe2_io_pipe_phv_out_data_455; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_456 = pipe2_io_pipe_phv_out_data_456; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_457 = pipe2_io_pipe_phv_out_data_457; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_458 = pipe2_io_pipe_phv_out_data_458; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_459 = pipe2_io_pipe_phv_out_data_459; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_460 = pipe2_io_pipe_phv_out_data_460; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_461 = pipe2_io_pipe_phv_out_data_461; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_462 = pipe2_io_pipe_phv_out_data_462; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_463 = pipe2_io_pipe_phv_out_data_463; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_464 = pipe2_io_pipe_phv_out_data_464; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_465 = pipe2_io_pipe_phv_out_data_465; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_466 = pipe2_io_pipe_phv_out_data_466; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_467 = pipe2_io_pipe_phv_out_data_467; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_468 = pipe2_io_pipe_phv_out_data_468; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_469 = pipe2_io_pipe_phv_out_data_469; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_470 = pipe2_io_pipe_phv_out_data_470; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_471 = pipe2_io_pipe_phv_out_data_471; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_472 = pipe2_io_pipe_phv_out_data_472; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_473 = pipe2_io_pipe_phv_out_data_473; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_474 = pipe2_io_pipe_phv_out_data_474; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_475 = pipe2_io_pipe_phv_out_data_475; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_476 = pipe2_io_pipe_phv_out_data_476; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_477 = pipe2_io_pipe_phv_out_data_477; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_478 = pipe2_io_pipe_phv_out_data_478; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_479 = pipe2_io_pipe_phv_out_data_479; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_480 = pipe2_io_pipe_phv_out_data_480; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_481 = pipe2_io_pipe_phv_out_data_481; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_482 = pipe2_io_pipe_phv_out_data_482; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_483 = pipe2_io_pipe_phv_out_data_483; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_484 = pipe2_io_pipe_phv_out_data_484; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_485 = pipe2_io_pipe_phv_out_data_485; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_486 = pipe2_io_pipe_phv_out_data_486; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_487 = pipe2_io_pipe_phv_out_data_487; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_488 = pipe2_io_pipe_phv_out_data_488; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_489 = pipe2_io_pipe_phv_out_data_489; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_490 = pipe2_io_pipe_phv_out_data_490; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_491 = pipe2_io_pipe_phv_out_data_491; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_492 = pipe2_io_pipe_phv_out_data_492; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_493 = pipe2_io_pipe_phv_out_data_493; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_494 = pipe2_io_pipe_phv_out_data_494; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_495 = pipe2_io_pipe_phv_out_data_495; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_496 = pipe2_io_pipe_phv_out_data_496; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_497 = pipe2_io_pipe_phv_out_data_497; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_498 = pipe2_io_pipe_phv_out_data_498; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_499 = pipe2_io_pipe_phv_out_data_499; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_500 = pipe2_io_pipe_phv_out_data_500; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_501 = pipe2_io_pipe_phv_out_data_501; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_502 = pipe2_io_pipe_phv_out_data_502; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_503 = pipe2_io_pipe_phv_out_data_503; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_504 = pipe2_io_pipe_phv_out_data_504; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_505 = pipe2_io_pipe_phv_out_data_505; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_506 = pipe2_io_pipe_phv_out_data_506; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_507 = pipe2_io_pipe_phv_out_data_507; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_508 = pipe2_io_pipe_phv_out_data_508; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_509 = pipe2_io_pipe_phv_out_data_509; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_510 = pipe2_io_pipe_phv_out_data_510; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_511 = pipe2_io_pipe_phv_out_data_511; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_0 = pipe2_io_pipe_phv_out_header_0; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_1 = pipe2_io_pipe_phv_out_header_1; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_2 = pipe2_io_pipe_phv_out_header_2; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_3 = pipe2_io_pipe_phv_out_header_3; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_4 = pipe2_io_pipe_phv_out_header_4; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_5 = pipe2_io_pipe_phv_out_header_5; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_6 = pipe2_io_pipe_phv_out_header_6; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_7 = pipe2_io_pipe_phv_out_header_7; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_8 = pipe2_io_pipe_phv_out_header_8; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_9 = pipe2_io_pipe_phv_out_header_9; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_10 = pipe2_io_pipe_phv_out_header_10; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_11 = pipe2_io_pipe_phv_out_header_11; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_12 = pipe2_io_pipe_phv_out_header_12; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_13 = pipe2_io_pipe_phv_out_header_13; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_14 = pipe2_io_pipe_phv_out_header_14; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_15 = pipe2_io_pipe_phv_out_header_15; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_parse_current_state = pipe2_io_pipe_phv_out_parse_current_state; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_parse_current_offset = pipe2_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_parse_transition_field = pipe2_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_next_processor_id = pipe2_io_pipe_phv_out_next_processor_id; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_next_config_id = pipe2_io_pipe_phv_out_next_config_id; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_is_valid_processor = pipe2_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 358:29]
  assign pipe3to8_io_mod_hash_depth_mod = io_mod_en; // @[matcher.scala 359:36]
  assign pipe3to8_io_mod_config_id = io_mod_config_id; // @[matcher.scala 360:36]
  assign pipe3to8_io_mod_hash_depth = io_mod_table_mod_table_depth[3:0]; // @[matcher.scala 361:36]
  assign pipe3to8_io_key_in = pipe2_io_match_key; // @[matcher.scala 362:26]
  assign pipe9_clock = clock;
  assign pipe9_io_pipe_phv_in_data_0 = pipe3to8_io_pipe_phv_out_data_0; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_1 = pipe3to8_io_pipe_phv_out_data_1; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_2 = pipe3to8_io_pipe_phv_out_data_2; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_3 = pipe3to8_io_pipe_phv_out_data_3; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_4 = pipe3to8_io_pipe_phv_out_data_4; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_5 = pipe3to8_io_pipe_phv_out_data_5; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_6 = pipe3to8_io_pipe_phv_out_data_6; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_7 = pipe3to8_io_pipe_phv_out_data_7; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_8 = pipe3to8_io_pipe_phv_out_data_8; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_9 = pipe3to8_io_pipe_phv_out_data_9; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_10 = pipe3to8_io_pipe_phv_out_data_10; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_11 = pipe3to8_io_pipe_phv_out_data_11; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_12 = pipe3to8_io_pipe_phv_out_data_12; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_13 = pipe3to8_io_pipe_phv_out_data_13; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_14 = pipe3to8_io_pipe_phv_out_data_14; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_15 = pipe3to8_io_pipe_phv_out_data_15; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_16 = pipe3to8_io_pipe_phv_out_data_16; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_17 = pipe3to8_io_pipe_phv_out_data_17; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_18 = pipe3to8_io_pipe_phv_out_data_18; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_19 = pipe3to8_io_pipe_phv_out_data_19; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_20 = pipe3to8_io_pipe_phv_out_data_20; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_21 = pipe3to8_io_pipe_phv_out_data_21; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_22 = pipe3to8_io_pipe_phv_out_data_22; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_23 = pipe3to8_io_pipe_phv_out_data_23; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_24 = pipe3to8_io_pipe_phv_out_data_24; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_25 = pipe3to8_io_pipe_phv_out_data_25; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_26 = pipe3to8_io_pipe_phv_out_data_26; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_27 = pipe3to8_io_pipe_phv_out_data_27; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_28 = pipe3to8_io_pipe_phv_out_data_28; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_29 = pipe3to8_io_pipe_phv_out_data_29; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_30 = pipe3to8_io_pipe_phv_out_data_30; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_31 = pipe3to8_io_pipe_phv_out_data_31; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_32 = pipe3to8_io_pipe_phv_out_data_32; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_33 = pipe3to8_io_pipe_phv_out_data_33; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_34 = pipe3to8_io_pipe_phv_out_data_34; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_35 = pipe3to8_io_pipe_phv_out_data_35; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_36 = pipe3to8_io_pipe_phv_out_data_36; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_37 = pipe3to8_io_pipe_phv_out_data_37; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_38 = pipe3to8_io_pipe_phv_out_data_38; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_39 = pipe3to8_io_pipe_phv_out_data_39; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_40 = pipe3to8_io_pipe_phv_out_data_40; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_41 = pipe3to8_io_pipe_phv_out_data_41; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_42 = pipe3to8_io_pipe_phv_out_data_42; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_43 = pipe3to8_io_pipe_phv_out_data_43; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_44 = pipe3to8_io_pipe_phv_out_data_44; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_45 = pipe3to8_io_pipe_phv_out_data_45; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_46 = pipe3to8_io_pipe_phv_out_data_46; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_47 = pipe3to8_io_pipe_phv_out_data_47; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_48 = pipe3to8_io_pipe_phv_out_data_48; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_49 = pipe3to8_io_pipe_phv_out_data_49; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_50 = pipe3to8_io_pipe_phv_out_data_50; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_51 = pipe3to8_io_pipe_phv_out_data_51; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_52 = pipe3to8_io_pipe_phv_out_data_52; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_53 = pipe3to8_io_pipe_phv_out_data_53; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_54 = pipe3to8_io_pipe_phv_out_data_54; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_55 = pipe3to8_io_pipe_phv_out_data_55; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_56 = pipe3to8_io_pipe_phv_out_data_56; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_57 = pipe3to8_io_pipe_phv_out_data_57; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_58 = pipe3to8_io_pipe_phv_out_data_58; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_59 = pipe3to8_io_pipe_phv_out_data_59; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_60 = pipe3to8_io_pipe_phv_out_data_60; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_61 = pipe3to8_io_pipe_phv_out_data_61; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_62 = pipe3to8_io_pipe_phv_out_data_62; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_63 = pipe3to8_io_pipe_phv_out_data_63; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_64 = pipe3to8_io_pipe_phv_out_data_64; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_65 = pipe3to8_io_pipe_phv_out_data_65; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_66 = pipe3to8_io_pipe_phv_out_data_66; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_67 = pipe3to8_io_pipe_phv_out_data_67; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_68 = pipe3to8_io_pipe_phv_out_data_68; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_69 = pipe3to8_io_pipe_phv_out_data_69; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_70 = pipe3to8_io_pipe_phv_out_data_70; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_71 = pipe3to8_io_pipe_phv_out_data_71; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_72 = pipe3to8_io_pipe_phv_out_data_72; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_73 = pipe3to8_io_pipe_phv_out_data_73; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_74 = pipe3to8_io_pipe_phv_out_data_74; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_75 = pipe3to8_io_pipe_phv_out_data_75; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_76 = pipe3to8_io_pipe_phv_out_data_76; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_77 = pipe3to8_io_pipe_phv_out_data_77; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_78 = pipe3to8_io_pipe_phv_out_data_78; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_79 = pipe3to8_io_pipe_phv_out_data_79; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_80 = pipe3to8_io_pipe_phv_out_data_80; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_81 = pipe3to8_io_pipe_phv_out_data_81; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_82 = pipe3to8_io_pipe_phv_out_data_82; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_83 = pipe3to8_io_pipe_phv_out_data_83; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_84 = pipe3to8_io_pipe_phv_out_data_84; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_85 = pipe3to8_io_pipe_phv_out_data_85; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_86 = pipe3to8_io_pipe_phv_out_data_86; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_87 = pipe3to8_io_pipe_phv_out_data_87; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_88 = pipe3to8_io_pipe_phv_out_data_88; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_89 = pipe3to8_io_pipe_phv_out_data_89; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_90 = pipe3to8_io_pipe_phv_out_data_90; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_91 = pipe3to8_io_pipe_phv_out_data_91; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_92 = pipe3to8_io_pipe_phv_out_data_92; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_93 = pipe3to8_io_pipe_phv_out_data_93; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_94 = pipe3to8_io_pipe_phv_out_data_94; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_95 = pipe3to8_io_pipe_phv_out_data_95; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_96 = pipe3to8_io_pipe_phv_out_data_96; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_97 = pipe3to8_io_pipe_phv_out_data_97; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_98 = pipe3to8_io_pipe_phv_out_data_98; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_99 = pipe3to8_io_pipe_phv_out_data_99; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_100 = pipe3to8_io_pipe_phv_out_data_100; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_101 = pipe3to8_io_pipe_phv_out_data_101; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_102 = pipe3to8_io_pipe_phv_out_data_102; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_103 = pipe3to8_io_pipe_phv_out_data_103; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_104 = pipe3to8_io_pipe_phv_out_data_104; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_105 = pipe3to8_io_pipe_phv_out_data_105; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_106 = pipe3to8_io_pipe_phv_out_data_106; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_107 = pipe3to8_io_pipe_phv_out_data_107; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_108 = pipe3to8_io_pipe_phv_out_data_108; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_109 = pipe3to8_io_pipe_phv_out_data_109; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_110 = pipe3to8_io_pipe_phv_out_data_110; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_111 = pipe3to8_io_pipe_phv_out_data_111; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_112 = pipe3to8_io_pipe_phv_out_data_112; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_113 = pipe3to8_io_pipe_phv_out_data_113; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_114 = pipe3to8_io_pipe_phv_out_data_114; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_115 = pipe3to8_io_pipe_phv_out_data_115; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_116 = pipe3to8_io_pipe_phv_out_data_116; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_117 = pipe3to8_io_pipe_phv_out_data_117; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_118 = pipe3to8_io_pipe_phv_out_data_118; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_119 = pipe3to8_io_pipe_phv_out_data_119; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_120 = pipe3to8_io_pipe_phv_out_data_120; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_121 = pipe3to8_io_pipe_phv_out_data_121; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_122 = pipe3to8_io_pipe_phv_out_data_122; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_123 = pipe3to8_io_pipe_phv_out_data_123; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_124 = pipe3to8_io_pipe_phv_out_data_124; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_125 = pipe3to8_io_pipe_phv_out_data_125; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_126 = pipe3to8_io_pipe_phv_out_data_126; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_127 = pipe3to8_io_pipe_phv_out_data_127; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_128 = pipe3to8_io_pipe_phv_out_data_128; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_129 = pipe3to8_io_pipe_phv_out_data_129; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_130 = pipe3to8_io_pipe_phv_out_data_130; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_131 = pipe3to8_io_pipe_phv_out_data_131; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_132 = pipe3to8_io_pipe_phv_out_data_132; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_133 = pipe3to8_io_pipe_phv_out_data_133; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_134 = pipe3to8_io_pipe_phv_out_data_134; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_135 = pipe3to8_io_pipe_phv_out_data_135; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_136 = pipe3to8_io_pipe_phv_out_data_136; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_137 = pipe3to8_io_pipe_phv_out_data_137; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_138 = pipe3to8_io_pipe_phv_out_data_138; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_139 = pipe3to8_io_pipe_phv_out_data_139; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_140 = pipe3to8_io_pipe_phv_out_data_140; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_141 = pipe3to8_io_pipe_phv_out_data_141; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_142 = pipe3to8_io_pipe_phv_out_data_142; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_143 = pipe3to8_io_pipe_phv_out_data_143; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_144 = pipe3to8_io_pipe_phv_out_data_144; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_145 = pipe3to8_io_pipe_phv_out_data_145; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_146 = pipe3to8_io_pipe_phv_out_data_146; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_147 = pipe3to8_io_pipe_phv_out_data_147; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_148 = pipe3to8_io_pipe_phv_out_data_148; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_149 = pipe3to8_io_pipe_phv_out_data_149; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_150 = pipe3to8_io_pipe_phv_out_data_150; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_151 = pipe3to8_io_pipe_phv_out_data_151; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_152 = pipe3to8_io_pipe_phv_out_data_152; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_153 = pipe3to8_io_pipe_phv_out_data_153; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_154 = pipe3to8_io_pipe_phv_out_data_154; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_155 = pipe3to8_io_pipe_phv_out_data_155; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_156 = pipe3to8_io_pipe_phv_out_data_156; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_157 = pipe3to8_io_pipe_phv_out_data_157; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_158 = pipe3to8_io_pipe_phv_out_data_158; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_159 = pipe3to8_io_pipe_phv_out_data_159; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_160 = pipe3to8_io_pipe_phv_out_data_160; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_161 = pipe3to8_io_pipe_phv_out_data_161; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_162 = pipe3to8_io_pipe_phv_out_data_162; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_163 = pipe3to8_io_pipe_phv_out_data_163; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_164 = pipe3to8_io_pipe_phv_out_data_164; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_165 = pipe3to8_io_pipe_phv_out_data_165; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_166 = pipe3to8_io_pipe_phv_out_data_166; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_167 = pipe3to8_io_pipe_phv_out_data_167; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_168 = pipe3to8_io_pipe_phv_out_data_168; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_169 = pipe3to8_io_pipe_phv_out_data_169; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_170 = pipe3to8_io_pipe_phv_out_data_170; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_171 = pipe3to8_io_pipe_phv_out_data_171; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_172 = pipe3to8_io_pipe_phv_out_data_172; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_173 = pipe3to8_io_pipe_phv_out_data_173; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_174 = pipe3to8_io_pipe_phv_out_data_174; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_175 = pipe3to8_io_pipe_phv_out_data_175; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_176 = pipe3to8_io_pipe_phv_out_data_176; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_177 = pipe3to8_io_pipe_phv_out_data_177; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_178 = pipe3to8_io_pipe_phv_out_data_178; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_179 = pipe3to8_io_pipe_phv_out_data_179; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_180 = pipe3to8_io_pipe_phv_out_data_180; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_181 = pipe3to8_io_pipe_phv_out_data_181; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_182 = pipe3to8_io_pipe_phv_out_data_182; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_183 = pipe3to8_io_pipe_phv_out_data_183; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_184 = pipe3to8_io_pipe_phv_out_data_184; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_185 = pipe3to8_io_pipe_phv_out_data_185; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_186 = pipe3to8_io_pipe_phv_out_data_186; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_187 = pipe3to8_io_pipe_phv_out_data_187; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_188 = pipe3to8_io_pipe_phv_out_data_188; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_189 = pipe3to8_io_pipe_phv_out_data_189; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_190 = pipe3to8_io_pipe_phv_out_data_190; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_191 = pipe3to8_io_pipe_phv_out_data_191; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_192 = pipe3to8_io_pipe_phv_out_data_192; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_193 = pipe3to8_io_pipe_phv_out_data_193; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_194 = pipe3to8_io_pipe_phv_out_data_194; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_195 = pipe3to8_io_pipe_phv_out_data_195; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_196 = pipe3to8_io_pipe_phv_out_data_196; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_197 = pipe3to8_io_pipe_phv_out_data_197; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_198 = pipe3to8_io_pipe_phv_out_data_198; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_199 = pipe3to8_io_pipe_phv_out_data_199; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_200 = pipe3to8_io_pipe_phv_out_data_200; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_201 = pipe3to8_io_pipe_phv_out_data_201; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_202 = pipe3to8_io_pipe_phv_out_data_202; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_203 = pipe3to8_io_pipe_phv_out_data_203; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_204 = pipe3to8_io_pipe_phv_out_data_204; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_205 = pipe3to8_io_pipe_phv_out_data_205; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_206 = pipe3to8_io_pipe_phv_out_data_206; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_207 = pipe3to8_io_pipe_phv_out_data_207; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_208 = pipe3to8_io_pipe_phv_out_data_208; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_209 = pipe3to8_io_pipe_phv_out_data_209; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_210 = pipe3to8_io_pipe_phv_out_data_210; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_211 = pipe3to8_io_pipe_phv_out_data_211; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_212 = pipe3to8_io_pipe_phv_out_data_212; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_213 = pipe3to8_io_pipe_phv_out_data_213; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_214 = pipe3to8_io_pipe_phv_out_data_214; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_215 = pipe3to8_io_pipe_phv_out_data_215; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_216 = pipe3to8_io_pipe_phv_out_data_216; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_217 = pipe3to8_io_pipe_phv_out_data_217; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_218 = pipe3to8_io_pipe_phv_out_data_218; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_219 = pipe3to8_io_pipe_phv_out_data_219; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_220 = pipe3to8_io_pipe_phv_out_data_220; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_221 = pipe3to8_io_pipe_phv_out_data_221; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_222 = pipe3to8_io_pipe_phv_out_data_222; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_223 = pipe3to8_io_pipe_phv_out_data_223; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_224 = pipe3to8_io_pipe_phv_out_data_224; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_225 = pipe3to8_io_pipe_phv_out_data_225; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_226 = pipe3to8_io_pipe_phv_out_data_226; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_227 = pipe3to8_io_pipe_phv_out_data_227; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_228 = pipe3to8_io_pipe_phv_out_data_228; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_229 = pipe3to8_io_pipe_phv_out_data_229; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_230 = pipe3to8_io_pipe_phv_out_data_230; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_231 = pipe3to8_io_pipe_phv_out_data_231; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_232 = pipe3to8_io_pipe_phv_out_data_232; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_233 = pipe3to8_io_pipe_phv_out_data_233; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_234 = pipe3to8_io_pipe_phv_out_data_234; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_235 = pipe3to8_io_pipe_phv_out_data_235; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_236 = pipe3to8_io_pipe_phv_out_data_236; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_237 = pipe3to8_io_pipe_phv_out_data_237; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_238 = pipe3to8_io_pipe_phv_out_data_238; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_239 = pipe3to8_io_pipe_phv_out_data_239; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_240 = pipe3to8_io_pipe_phv_out_data_240; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_241 = pipe3to8_io_pipe_phv_out_data_241; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_242 = pipe3to8_io_pipe_phv_out_data_242; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_243 = pipe3to8_io_pipe_phv_out_data_243; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_244 = pipe3to8_io_pipe_phv_out_data_244; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_245 = pipe3to8_io_pipe_phv_out_data_245; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_246 = pipe3to8_io_pipe_phv_out_data_246; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_247 = pipe3to8_io_pipe_phv_out_data_247; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_248 = pipe3to8_io_pipe_phv_out_data_248; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_249 = pipe3to8_io_pipe_phv_out_data_249; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_250 = pipe3to8_io_pipe_phv_out_data_250; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_251 = pipe3to8_io_pipe_phv_out_data_251; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_252 = pipe3to8_io_pipe_phv_out_data_252; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_253 = pipe3to8_io_pipe_phv_out_data_253; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_254 = pipe3to8_io_pipe_phv_out_data_254; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_255 = pipe3to8_io_pipe_phv_out_data_255; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_256 = pipe3to8_io_pipe_phv_out_data_256; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_257 = pipe3to8_io_pipe_phv_out_data_257; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_258 = pipe3to8_io_pipe_phv_out_data_258; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_259 = pipe3to8_io_pipe_phv_out_data_259; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_260 = pipe3to8_io_pipe_phv_out_data_260; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_261 = pipe3to8_io_pipe_phv_out_data_261; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_262 = pipe3to8_io_pipe_phv_out_data_262; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_263 = pipe3to8_io_pipe_phv_out_data_263; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_264 = pipe3to8_io_pipe_phv_out_data_264; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_265 = pipe3to8_io_pipe_phv_out_data_265; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_266 = pipe3to8_io_pipe_phv_out_data_266; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_267 = pipe3to8_io_pipe_phv_out_data_267; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_268 = pipe3to8_io_pipe_phv_out_data_268; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_269 = pipe3to8_io_pipe_phv_out_data_269; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_270 = pipe3to8_io_pipe_phv_out_data_270; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_271 = pipe3to8_io_pipe_phv_out_data_271; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_272 = pipe3to8_io_pipe_phv_out_data_272; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_273 = pipe3to8_io_pipe_phv_out_data_273; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_274 = pipe3to8_io_pipe_phv_out_data_274; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_275 = pipe3to8_io_pipe_phv_out_data_275; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_276 = pipe3to8_io_pipe_phv_out_data_276; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_277 = pipe3to8_io_pipe_phv_out_data_277; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_278 = pipe3to8_io_pipe_phv_out_data_278; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_279 = pipe3to8_io_pipe_phv_out_data_279; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_280 = pipe3to8_io_pipe_phv_out_data_280; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_281 = pipe3to8_io_pipe_phv_out_data_281; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_282 = pipe3to8_io_pipe_phv_out_data_282; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_283 = pipe3to8_io_pipe_phv_out_data_283; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_284 = pipe3to8_io_pipe_phv_out_data_284; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_285 = pipe3to8_io_pipe_phv_out_data_285; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_286 = pipe3to8_io_pipe_phv_out_data_286; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_287 = pipe3to8_io_pipe_phv_out_data_287; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_288 = pipe3to8_io_pipe_phv_out_data_288; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_289 = pipe3to8_io_pipe_phv_out_data_289; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_290 = pipe3to8_io_pipe_phv_out_data_290; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_291 = pipe3to8_io_pipe_phv_out_data_291; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_292 = pipe3to8_io_pipe_phv_out_data_292; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_293 = pipe3to8_io_pipe_phv_out_data_293; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_294 = pipe3to8_io_pipe_phv_out_data_294; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_295 = pipe3to8_io_pipe_phv_out_data_295; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_296 = pipe3to8_io_pipe_phv_out_data_296; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_297 = pipe3to8_io_pipe_phv_out_data_297; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_298 = pipe3to8_io_pipe_phv_out_data_298; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_299 = pipe3to8_io_pipe_phv_out_data_299; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_300 = pipe3to8_io_pipe_phv_out_data_300; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_301 = pipe3to8_io_pipe_phv_out_data_301; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_302 = pipe3to8_io_pipe_phv_out_data_302; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_303 = pipe3to8_io_pipe_phv_out_data_303; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_304 = pipe3to8_io_pipe_phv_out_data_304; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_305 = pipe3to8_io_pipe_phv_out_data_305; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_306 = pipe3to8_io_pipe_phv_out_data_306; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_307 = pipe3to8_io_pipe_phv_out_data_307; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_308 = pipe3to8_io_pipe_phv_out_data_308; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_309 = pipe3to8_io_pipe_phv_out_data_309; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_310 = pipe3to8_io_pipe_phv_out_data_310; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_311 = pipe3to8_io_pipe_phv_out_data_311; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_312 = pipe3to8_io_pipe_phv_out_data_312; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_313 = pipe3to8_io_pipe_phv_out_data_313; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_314 = pipe3to8_io_pipe_phv_out_data_314; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_315 = pipe3to8_io_pipe_phv_out_data_315; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_316 = pipe3to8_io_pipe_phv_out_data_316; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_317 = pipe3to8_io_pipe_phv_out_data_317; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_318 = pipe3to8_io_pipe_phv_out_data_318; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_319 = pipe3to8_io_pipe_phv_out_data_319; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_320 = pipe3to8_io_pipe_phv_out_data_320; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_321 = pipe3to8_io_pipe_phv_out_data_321; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_322 = pipe3to8_io_pipe_phv_out_data_322; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_323 = pipe3to8_io_pipe_phv_out_data_323; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_324 = pipe3to8_io_pipe_phv_out_data_324; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_325 = pipe3to8_io_pipe_phv_out_data_325; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_326 = pipe3to8_io_pipe_phv_out_data_326; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_327 = pipe3to8_io_pipe_phv_out_data_327; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_328 = pipe3to8_io_pipe_phv_out_data_328; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_329 = pipe3to8_io_pipe_phv_out_data_329; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_330 = pipe3to8_io_pipe_phv_out_data_330; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_331 = pipe3to8_io_pipe_phv_out_data_331; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_332 = pipe3to8_io_pipe_phv_out_data_332; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_333 = pipe3to8_io_pipe_phv_out_data_333; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_334 = pipe3to8_io_pipe_phv_out_data_334; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_335 = pipe3to8_io_pipe_phv_out_data_335; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_336 = pipe3to8_io_pipe_phv_out_data_336; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_337 = pipe3to8_io_pipe_phv_out_data_337; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_338 = pipe3to8_io_pipe_phv_out_data_338; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_339 = pipe3to8_io_pipe_phv_out_data_339; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_340 = pipe3to8_io_pipe_phv_out_data_340; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_341 = pipe3to8_io_pipe_phv_out_data_341; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_342 = pipe3to8_io_pipe_phv_out_data_342; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_343 = pipe3to8_io_pipe_phv_out_data_343; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_344 = pipe3to8_io_pipe_phv_out_data_344; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_345 = pipe3to8_io_pipe_phv_out_data_345; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_346 = pipe3to8_io_pipe_phv_out_data_346; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_347 = pipe3to8_io_pipe_phv_out_data_347; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_348 = pipe3to8_io_pipe_phv_out_data_348; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_349 = pipe3to8_io_pipe_phv_out_data_349; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_350 = pipe3to8_io_pipe_phv_out_data_350; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_351 = pipe3to8_io_pipe_phv_out_data_351; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_352 = pipe3to8_io_pipe_phv_out_data_352; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_353 = pipe3to8_io_pipe_phv_out_data_353; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_354 = pipe3to8_io_pipe_phv_out_data_354; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_355 = pipe3to8_io_pipe_phv_out_data_355; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_356 = pipe3to8_io_pipe_phv_out_data_356; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_357 = pipe3to8_io_pipe_phv_out_data_357; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_358 = pipe3to8_io_pipe_phv_out_data_358; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_359 = pipe3to8_io_pipe_phv_out_data_359; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_360 = pipe3to8_io_pipe_phv_out_data_360; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_361 = pipe3to8_io_pipe_phv_out_data_361; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_362 = pipe3to8_io_pipe_phv_out_data_362; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_363 = pipe3to8_io_pipe_phv_out_data_363; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_364 = pipe3to8_io_pipe_phv_out_data_364; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_365 = pipe3to8_io_pipe_phv_out_data_365; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_366 = pipe3to8_io_pipe_phv_out_data_366; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_367 = pipe3to8_io_pipe_phv_out_data_367; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_368 = pipe3to8_io_pipe_phv_out_data_368; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_369 = pipe3to8_io_pipe_phv_out_data_369; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_370 = pipe3to8_io_pipe_phv_out_data_370; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_371 = pipe3to8_io_pipe_phv_out_data_371; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_372 = pipe3to8_io_pipe_phv_out_data_372; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_373 = pipe3to8_io_pipe_phv_out_data_373; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_374 = pipe3to8_io_pipe_phv_out_data_374; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_375 = pipe3to8_io_pipe_phv_out_data_375; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_376 = pipe3to8_io_pipe_phv_out_data_376; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_377 = pipe3to8_io_pipe_phv_out_data_377; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_378 = pipe3to8_io_pipe_phv_out_data_378; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_379 = pipe3to8_io_pipe_phv_out_data_379; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_380 = pipe3to8_io_pipe_phv_out_data_380; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_381 = pipe3to8_io_pipe_phv_out_data_381; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_382 = pipe3to8_io_pipe_phv_out_data_382; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_383 = pipe3to8_io_pipe_phv_out_data_383; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_384 = pipe3to8_io_pipe_phv_out_data_384; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_385 = pipe3to8_io_pipe_phv_out_data_385; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_386 = pipe3to8_io_pipe_phv_out_data_386; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_387 = pipe3to8_io_pipe_phv_out_data_387; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_388 = pipe3to8_io_pipe_phv_out_data_388; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_389 = pipe3to8_io_pipe_phv_out_data_389; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_390 = pipe3to8_io_pipe_phv_out_data_390; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_391 = pipe3to8_io_pipe_phv_out_data_391; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_392 = pipe3to8_io_pipe_phv_out_data_392; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_393 = pipe3to8_io_pipe_phv_out_data_393; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_394 = pipe3to8_io_pipe_phv_out_data_394; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_395 = pipe3to8_io_pipe_phv_out_data_395; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_396 = pipe3to8_io_pipe_phv_out_data_396; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_397 = pipe3to8_io_pipe_phv_out_data_397; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_398 = pipe3to8_io_pipe_phv_out_data_398; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_399 = pipe3to8_io_pipe_phv_out_data_399; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_400 = pipe3to8_io_pipe_phv_out_data_400; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_401 = pipe3to8_io_pipe_phv_out_data_401; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_402 = pipe3to8_io_pipe_phv_out_data_402; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_403 = pipe3to8_io_pipe_phv_out_data_403; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_404 = pipe3to8_io_pipe_phv_out_data_404; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_405 = pipe3to8_io_pipe_phv_out_data_405; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_406 = pipe3to8_io_pipe_phv_out_data_406; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_407 = pipe3to8_io_pipe_phv_out_data_407; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_408 = pipe3to8_io_pipe_phv_out_data_408; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_409 = pipe3to8_io_pipe_phv_out_data_409; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_410 = pipe3to8_io_pipe_phv_out_data_410; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_411 = pipe3to8_io_pipe_phv_out_data_411; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_412 = pipe3to8_io_pipe_phv_out_data_412; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_413 = pipe3to8_io_pipe_phv_out_data_413; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_414 = pipe3to8_io_pipe_phv_out_data_414; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_415 = pipe3to8_io_pipe_phv_out_data_415; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_416 = pipe3to8_io_pipe_phv_out_data_416; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_417 = pipe3to8_io_pipe_phv_out_data_417; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_418 = pipe3to8_io_pipe_phv_out_data_418; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_419 = pipe3to8_io_pipe_phv_out_data_419; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_420 = pipe3to8_io_pipe_phv_out_data_420; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_421 = pipe3to8_io_pipe_phv_out_data_421; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_422 = pipe3to8_io_pipe_phv_out_data_422; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_423 = pipe3to8_io_pipe_phv_out_data_423; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_424 = pipe3to8_io_pipe_phv_out_data_424; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_425 = pipe3to8_io_pipe_phv_out_data_425; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_426 = pipe3to8_io_pipe_phv_out_data_426; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_427 = pipe3to8_io_pipe_phv_out_data_427; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_428 = pipe3to8_io_pipe_phv_out_data_428; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_429 = pipe3to8_io_pipe_phv_out_data_429; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_430 = pipe3to8_io_pipe_phv_out_data_430; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_431 = pipe3to8_io_pipe_phv_out_data_431; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_432 = pipe3to8_io_pipe_phv_out_data_432; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_433 = pipe3to8_io_pipe_phv_out_data_433; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_434 = pipe3to8_io_pipe_phv_out_data_434; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_435 = pipe3to8_io_pipe_phv_out_data_435; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_436 = pipe3to8_io_pipe_phv_out_data_436; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_437 = pipe3to8_io_pipe_phv_out_data_437; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_438 = pipe3to8_io_pipe_phv_out_data_438; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_439 = pipe3to8_io_pipe_phv_out_data_439; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_440 = pipe3to8_io_pipe_phv_out_data_440; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_441 = pipe3to8_io_pipe_phv_out_data_441; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_442 = pipe3to8_io_pipe_phv_out_data_442; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_443 = pipe3to8_io_pipe_phv_out_data_443; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_444 = pipe3to8_io_pipe_phv_out_data_444; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_445 = pipe3to8_io_pipe_phv_out_data_445; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_446 = pipe3to8_io_pipe_phv_out_data_446; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_447 = pipe3to8_io_pipe_phv_out_data_447; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_448 = pipe3to8_io_pipe_phv_out_data_448; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_449 = pipe3to8_io_pipe_phv_out_data_449; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_450 = pipe3to8_io_pipe_phv_out_data_450; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_451 = pipe3to8_io_pipe_phv_out_data_451; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_452 = pipe3to8_io_pipe_phv_out_data_452; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_453 = pipe3to8_io_pipe_phv_out_data_453; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_454 = pipe3to8_io_pipe_phv_out_data_454; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_455 = pipe3to8_io_pipe_phv_out_data_455; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_456 = pipe3to8_io_pipe_phv_out_data_456; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_457 = pipe3to8_io_pipe_phv_out_data_457; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_458 = pipe3to8_io_pipe_phv_out_data_458; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_459 = pipe3to8_io_pipe_phv_out_data_459; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_460 = pipe3to8_io_pipe_phv_out_data_460; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_461 = pipe3to8_io_pipe_phv_out_data_461; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_462 = pipe3to8_io_pipe_phv_out_data_462; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_463 = pipe3to8_io_pipe_phv_out_data_463; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_464 = pipe3to8_io_pipe_phv_out_data_464; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_465 = pipe3to8_io_pipe_phv_out_data_465; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_466 = pipe3to8_io_pipe_phv_out_data_466; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_467 = pipe3to8_io_pipe_phv_out_data_467; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_468 = pipe3to8_io_pipe_phv_out_data_468; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_469 = pipe3to8_io_pipe_phv_out_data_469; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_470 = pipe3to8_io_pipe_phv_out_data_470; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_471 = pipe3to8_io_pipe_phv_out_data_471; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_472 = pipe3to8_io_pipe_phv_out_data_472; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_473 = pipe3to8_io_pipe_phv_out_data_473; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_474 = pipe3to8_io_pipe_phv_out_data_474; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_475 = pipe3to8_io_pipe_phv_out_data_475; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_476 = pipe3to8_io_pipe_phv_out_data_476; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_477 = pipe3to8_io_pipe_phv_out_data_477; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_478 = pipe3to8_io_pipe_phv_out_data_478; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_479 = pipe3to8_io_pipe_phv_out_data_479; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_480 = pipe3to8_io_pipe_phv_out_data_480; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_481 = pipe3to8_io_pipe_phv_out_data_481; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_482 = pipe3to8_io_pipe_phv_out_data_482; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_483 = pipe3to8_io_pipe_phv_out_data_483; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_484 = pipe3to8_io_pipe_phv_out_data_484; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_485 = pipe3to8_io_pipe_phv_out_data_485; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_486 = pipe3to8_io_pipe_phv_out_data_486; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_487 = pipe3to8_io_pipe_phv_out_data_487; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_488 = pipe3to8_io_pipe_phv_out_data_488; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_489 = pipe3to8_io_pipe_phv_out_data_489; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_490 = pipe3to8_io_pipe_phv_out_data_490; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_491 = pipe3to8_io_pipe_phv_out_data_491; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_492 = pipe3to8_io_pipe_phv_out_data_492; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_493 = pipe3to8_io_pipe_phv_out_data_493; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_494 = pipe3to8_io_pipe_phv_out_data_494; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_495 = pipe3to8_io_pipe_phv_out_data_495; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_496 = pipe3to8_io_pipe_phv_out_data_496; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_497 = pipe3to8_io_pipe_phv_out_data_497; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_498 = pipe3to8_io_pipe_phv_out_data_498; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_499 = pipe3to8_io_pipe_phv_out_data_499; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_500 = pipe3to8_io_pipe_phv_out_data_500; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_501 = pipe3to8_io_pipe_phv_out_data_501; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_502 = pipe3to8_io_pipe_phv_out_data_502; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_503 = pipe3to8_io_pipe_phv_out_data_503; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_504 = pipe3to8_io_pipe_phv_out_data_504; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_505 = pipe3to8_io_pipe_phv_out_data_505; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_506 = pipe3to8_io_pipe_phv_out_data_506; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_507 = pipe3to8_io_pipe_phv_out_data_507; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_508 = pipe3to8_io_pipe_phv_out_data_508; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_509 = pipe3to8_io_pipe_phv_out_data_509; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_510 = pipe3to8_io_pipe_phv_out_data_510; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_511 = pipe3to8_io_pipe_phv_out_data_511; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_0 = pipe3to8_io_pipe_phv_out_header_0; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_1 = pipe3to8_io_pipe_phv_out_header_1; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_2 = pipe3to8_io_pipe_phv_out_header_2; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_3 = pipe3to8_io_pipe_phv_out_header_3; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_4 = pipe3to8_io_pipe_phv_out_header_4; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_5 = pipe3to8_io_pipe_phv_out_header_5; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_6 = pipe3to8_io_pipe_phv_out_header_6; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_7 = pipe3to8_io_pipe_phv_out_header_7; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_8 = pipe3to8_io_pipe_phv_out_header_8; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_9 = pipe3to8_io_pipe_phv_out_header_9; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_10 = pipe3to8_io_pipe_phv_out_header_10; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_11 = pipe3to8_io_pipe_phv_out_header_11; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_12 = pipe3to8_io_pipe_phv_out_header_12; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_13 = pipe3to8_io_pipe_phv_out_header_13; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_14 = pipe3to8_io_pipe_phv_out_header_14; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_15 = pipe3to8_io_pipe_phv_out_header_15; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_parse_current_state = pipe3to8_io_pipe_phv_out_parse_current_state; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_parse_current_offset = pipe3to8_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_parse_transition_field = pipe3to8_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_next_processor_id = pipe3to8_io_pipe_phv_out_next_processor_id; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_next_config_id = pipe3to8_io_pipe_phv_out_next_config_id; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_is_valid_processor = pipe3to8_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 364:27]
  assign pipe9_io_table_config_0_table_width = table_config_0_table_width; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_table_depth = table_config_0_table_depth; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_table_width = table_config_1_table_width; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_table_depth = table_config_1_table_depth; // @[matcher.scala 368:27]
  assign pipe9_io_key_in = pipe3to8_io_key_out; // @[matcher.scala 365:27]
  assign pipe9_io_addr_in = pipe3to8_io_hash_val; // @[matcher.scala 366:27]
  assign pipe9_io_cs_in = pipe3to8_io_hash_val_cs; // @[matcher.scala 367:27]
  assign pipe10_clock = clock;
  assign pipe10_io_pipe_phv_in_data_0 = pipe9_io_pipe_phv_out_data_0; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_1 = pipe9_io_pipe_phv_out_data_1; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_2 = pipe9_io_pipe_phv_out_data_2; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_3 = pipe9_io_pipe_phv_out_data_3; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_4 = pipe9_io_pipe_phv_out_data_4; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_5 = pipe9_io_pipe_phv_out_data_5; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_6 = pipe9_io_pipe_phv_out_data_6; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_7 = pipe9_io_pipe_phv_out_data_7; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_8 = pipe9_io_pipe_phv_out_data_8; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_9 = pipe9_io_pipe_phv_out_data_9; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_10 = pipe9_io_pipe_phv_out_data_10; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_11 = pipe9_io_pipe_phv_out_data_11; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_12 = pipe9_io_pipe_phv_out_data_12; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_13 = pipe9_io_pipe_phv_out_data_13; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_14 = pipe9_io_pipe_phv_out_data_14; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_15 = pipe9_io_pipe_phv_out_data_15; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_16 = pipe9_io_pipe_phv_out_data_16; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_17 = pipe9_io_pipe_phv_out_data_17; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_18 = pipe9_io_pipe_phv_out_data_18; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_19 = pipe9_io_pipe_phv_out_data_19; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_20 = pipe9_io_pipe_phv_out_data_20; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_21 = pipe9_io_pipe_phv_out_data_21; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_22 = pipe9_io_pipe_phv_out_data_22; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_23 = pipe9_io_pipe_phv_out_data_23; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_24 = pipe9_io_pipe_phv_out_data_24; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_25 = pipe9_io_pipe_phv_out_data_25; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_26 = pipe9_io_pipe_phv_out_data_26; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_27 = pipe9_io_pipe_phv_out_data_27; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_28 = pipe9_io_pipe_phv_out_data_28; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_29 = pipe9_io_pipe_phv_out_data_29; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_30 = pipe9_io_pipe_phv_out_data_30; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_31 = pipe9_io_pipe_phv_out_data_31; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_32 = pipe9_io_pipe_phv_out_data_32; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_33 = pipe9_io_pipe_phv_out_data_33; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_34 = pipe9_io_pipe_phv_out_data_34; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_35 = pipe9_io_pipe_phv_out_data_35; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_36 = pipe9_io_pipe_phv_out_data_36; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_37 = pipe9_io_pipe_phv_out_data_37; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_38 = pipe9_io_pipe_phv_out_data_38; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_39 = pipe9_io_pipe_phv_out_data_39; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_40 = pipe9_io_pipe_phv_out_data_40; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_41 = pipe9_io_pipe_phv_out_data_41; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_42 = pipe9_io_pipe_phv_out_data_42; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_43 = pipe9_io_pipe_phv_out_data_43; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_44 = pipe9_io_pipe_phv_out_data_44; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_45 = pipe9_io_pipe_phv_out_data_45; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_46 = pipe9_io_pipe_phv_out_data_46; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_47 = pipe9_io_pipe_phv_out_data_47; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_48 = pipe9_io_pipe_phv_out_data_48; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_49 = pipe9_io_pipe_phv_out_data_49; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_50 = pipe9_io_pipe_phv_out_data_50; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_51 = pipe9_io_pipe_phv_out_data_51; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_52 = pipe9_io_pipe_phv_out_data_52; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_53 = pipe9_io_pipe_phv_out_data_53; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_54 = pipe9_io_pipe_phv_out_data_54; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_55 = pipe9_io_pipe_phv_out_data_55; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_56 = pipe9_io_pipe_phv_out_data_56; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_57 = pipe9_io_pipe_phv_out_data_57; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_58 = pipe9_io_pipe_phv_out_data_58; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_59 = pipe9_io_pipe_phv_out_data_59; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_60 = pipe9_io_pipe_phv_out_data_60; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_61 = pipe9_io_pipe_phv_out_data_61; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_62 = pipe9_io_pipe_phv_out_data_62; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_63 = pipe9_io_pipe_phv_out_data_63; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_64 = pipe9_io_pipe_phv_out_data_64; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_65 = pipe9_io_pipe_phv_out_data_65; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_66 = pipe9_io_pipe_phv_out_data_66; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_67 = pipe9_io_pipe_phv_out_data_67; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_68 = pipe9_io_pipe_phv_out_data_68; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_69 = pipe9_io_pipe_phv_out_data_69; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_70 = pipe9_io_pipe_phv_out_data_70; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_71 = pipe9_io_pipe_phv_out_data_71; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_72 = pipe9_io_pipe_phv_out_data_72; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_73 = pipe9_io_pipe_phv_out_data_73; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_74 = pipe9_io_pipe_phv_out_data_74; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_75 = pipe9_io_pipe_phv_out_data_75; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_76 = pipe9_io_pipe_phv_out_data_76; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_77 = pipe9_io_pipe_phv_out_data_77; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_78 = pipe9_io_pipe_phv_out_data_78; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_79 = pipe9_io_pipe_phv_out_data_79; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_80 = pipe9_io_pipe_phv_out_data_80; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_81 = pipe9_io_pipe_phv_out_data_81; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_82 = pipe9_io_pipe_phv_out_data_82; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_83 = pipe9_io_pipe_phv_out_data_83; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_84 = pipe9_io_pipe_phv_out_data_84; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_85 = pipe9_io_pipe_phv_out_data_85; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_86 = pipe9_io_pipe_phv_out_data_86; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_87 = pipe9_io_pipe_phv_out_data_87; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_88 = pipe9_io_pipe_phv_out_data_88; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_89 = pipe9_io_pipe_phv_out_data_89; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_90 = pipe9_io_pipe_phv_out_data_90; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_91 = pipe9_io_pipe_phv_out_data_91; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_92 = pipe9_io_pipe_phv_out_data_92; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_93 = pipe9_io_pipe_phv_out_data_93; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_94 = pipe9_io_pipe_phv_out_data_94; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_95 = pipe9_io_pipe_phv_out_data_95; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_96 = pipe9_io_pipe_phv_out_data_96; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_97 = pipe9_io_pipe_phv_out_data_97; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_98 = pipe9_io_pipe_phv_out_data_98; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_99 = pipe9_io_pipe_phv_out_data_99; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_100 = pipe9_io_pipe_phv_out_data_100; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_101 = pipe9_io_pipe_phv_out_data_101; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_102 = pipe9_io_pipe_phv_out_data_102; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_103 = pipe9_io_pipe_phv_out_data_103; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_104 = pipe9_io_pipe_phv_out_data_104; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_105 = pipe9_io_pipe_phv_out_data_105; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_106 = pipe9_io_pipe_phv_out_data_106; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_107 = pipe9_io_pipe_phv_out_data_107; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_108 = pipe9_io_pipe_phv_out_data_108; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_109 = pipe9_io_pipe_phv_out_data_109; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_110 = pipe9_io_pipe_phv_out_data_110; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_111 = pipe9_io_pipe_phv_out_data_111; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_112 = pipe9_io_pipe_phv_out_data_112; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_113 = pipe9_io_pipe_phv_out_data_113; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_114 = pipe9_io_pipe_phv_out_data_114; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_115 = pipe9_io_pipe_phv_out_data_115; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_116 = pipe9_io_pipe_phv_out_data_116; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_117 = pipe9_io_pipe_phv_out_data_117; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_118 = pipe9_io_pipe_phv_out_data_118; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_119 = pipe9_io_pipe_phv_out_data_119; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_120 = pipe9_io_pipe_phv_out_data_120; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_121 = pipe9_io_pipe_phv_out_data_121; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_122 = pipe9_io_pipe_phv_out_data_122; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_123 = pipe9_io_pipe_phv_out_data_123; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_124 = pipe9_io_pipe_phv_out_data_124; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_125 = pipe9_io_pipe_phv_out_data_125; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_126 = pipe9_io_pipe_phv_out_data_126; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_127 = pipe9_io_pipe_phv_out_data_127; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_128 = pipe9_io_pipe_phv_out_data_128; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_129 = pipe9_io_pipe_phv_out_data_129; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_130 = pipe9_io_pipe_phv_out_data_130; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_131 = pipe9_io_pipe_phv_out_data_131; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_132 = pipe9_io_pipe_phv_out_data_132; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_133 = pipe9_io_pipe_phv_out_data_133; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_134 = pipe9_io_pipe_phv_out_data_134; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_135 = pipe9_io_pipe_phv_out_data_135; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_136 = pipe9_io_pipe_phv_out_data_136; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_137 = pipe9_io_pipe_phv_out_data_137; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_138 = pipe9_io_pipe_phv_out_data_138; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_139 = pipe9_io_pipe_phv_out_data_139; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_140 = pipe9_io_pipe_phv_out_data_140; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_141 = pipe9_io_pipe_phv_out_data_141; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_142 = pipe9_io_pipe_phv_out_data_142; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_143 = pipe9_io_pipe_phv_out_data_143; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_144 = pipe9_io_pipe_phv_out_data_144; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_145 = pipe9_io_pipe_phv_out_data_145; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_146 = pipe9_io_pipe_phv_out_data_146; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_147 = pipe9_io_pipe_phv_out_data_147; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_148 = pipe9_io_pipe_phv_out_data_148; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_149 = pipe9_io_pipe_phv_out_data_149; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_150 = pipe9_io_pipe_phv_out_data_150; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_151 = pipe9_io_pipe_phv_out_data_151; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_152 = pipe9_io_pipe_phv_out_data_152; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_153 = pipe9_io_pipe_phv_out_data_153; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_154 = pipe9_io_pipe_phv_out_data_154; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_155 = pipe9_io_pipe_phv_out_data_155; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_156 = pipe9_io_pipe_phv_out_data_156; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_157 = pipe9_io_pipe_phv_out_data_157; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_158 = pipe9_io_pipe_phv_out_data_158; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_159 = pipe9_io_pipe_phv_out_data_159; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_160 = pipe9_io_pipe_phv_out_data_160; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_161 = pipe9_io_pipe_phv_out_data_161; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_162 = pipe9_io_pipe_phv_out_data_162; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_163 = pipe9_io_pipe_phv_out_data_163; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_164 = pipe9_io_pipe_phv_out_data_164; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_165 = pipe9_io_pipe_phv_out_data_165; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_166 = pipe9_io_pipe_phv_out_data_166; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_167 = pipe9_io_pipe_phv_out_data_167; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_168 = pipe9_io_pipe_phv_out_data_168; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_169 = pipe9_io_pipe_phv_out_data_169; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_170 = pipe9_io_pipe_phv_out_data_170; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_171 = pipe9_io_pipe_phv_out_data_171; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_172 = pipe9_io_pipe_phv_out_data_172; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_173 = pipe9_io_pipe_phv_out_data_173; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_174 = pipe9_io_pipe_phv_out_data_174; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_175 = pipe9_io_pipe_phv_out_data_175; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_176 = pipe9_io_pipe_phv_out_data_176; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_177 = pipe9_io_pipe_phv_out_data_177; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_178 = pipe9_io_pipe_phv_out_data_178; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_179 = pipe9_io_pipe_phv_out_data_179; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_180 = pipe9_io_pipe_phv_out_data_180; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_181 = pipe9_io_pipe_phv_out_data_181; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_182 = pipe9_io_pipe_phv_out_data_182; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_183 = pipe9_io_pipe_phv_out_data_183; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_184 = pipe9_io_pipe_phv_out_data_184; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_185 = pipe9_io_pipe_phv_out_data_185; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_186 = pipe9_io_pipe_phv_out_data_186; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_187 = pipe9_io_pipe_phv_out_data_187; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_188 = pipe9_io_pipe_phv_out_data_188; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_189 = pipe9_io_pipe_phv_out_data_189; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_190 = pipe9_io_pipe_phv_out_data_190; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_191 = pipe9_io_pipe_phv_out_data_191; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_192 = pipe9_io_pipe_phv_out_data_192; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_193 = pipe9_io_pipe_phv_out_data_193; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_194 = pipe9_io_pipe_phv_out_data_194; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_195 = pipe9_io_pipe_phv_out_data_195; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_196 = pipe9_io_pipe_phv_out_data_196; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_197 = pipe9_io_pipe_phv_out_data_197; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_198 = pipe9_io_pipe_phv_out_data_198; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_199 = pipe9_io_pipe_phv_out_data_199; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_200 = pipe9_io_pipe_phv_out_data_200; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_201 = pipe9_io_pipe_phv_out_data_201; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_202 = pipe9_io_pipe_phv_out_data_202; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_203 = pipe9_io_pipe_phv_out_data_203; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_204 = pipe9_io_pipe_phv_out_data_204; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_205 = pipe9_io_pipe_phv_out_data_205; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_206 = pipe9_io_pipe_phv_out_data_206; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_207 = pipe9_io_pipe_phv_out_data_207; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_208 = pipe9_io_pipe_phv_out_data_208; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_209 = pipe9_io_pipe_phv_out_data_209; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_210 = pipe9_io_pipe_phv_out_data_210; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_211 = pipe9_io_pipe_phv_out_data_211; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_212 = pipe9_io_pipe_phv_out_data_212; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_213 = pipe9_io_pipe_phv_out_data_213; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_214 = pipe9_io_pipe_phv_out_data_214; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_215 = pipe9_io_pipe_phv_out_data_215; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_216 = pipe9_io_pipe_phv_out_data_216; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_217 = pipe9_io_pipe_phv_out_data_217; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_218 = pipe9_io_pipe_phv_out_data_218; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_219 = pipe9_io_pipe_phv_out_data_219; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_220 = pipe9_io_pipe_phv_out_data_220; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_221 = pipe9_io_pipe_phv_out_data_221; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_222 = pipe9_io_pipe_phv_out_data_222; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_223 = pipe9_io_pipe_phv_out_data_223; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_224 = pipe9_io_pipe_phv_out_data_224; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_225 = pipe9_io_pipe_phv_out_data_225; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_226 = pipe9_io_pipe_phv_out_data_226; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_227 = pipe9_io_pipe_phv_out_data_227; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_228 = pipe9_io_pipe_phv_out_data_228; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_229 = pipe9_io_pipe_phv_out_data_229; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_230 = pipe9_io_pipe_phv_out_data_230; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_231 = pipe9_io_pipe_phv_out_data_231; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_232 = pipe9_io_pipe_phv_out_data_232; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_233 = pipe9_io_pipe_phv_out_data_233; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_234 = pipe9_io_pipe_phv_out_data_234; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_235 = pipe9_io_pipe_phv_out_data_235; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_236 = pipe9_io_pipe_phv_out_data_236; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_237 = pipe9_io_pipe_phv_out_data_237; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_238 = pipe9_io_pipe_phv_out_data_238; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_239 = pipe9_io_pipe_phv_out_data_239; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_240 = pipe9_io_pipe_phv_out_data_240; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_241 = pipe9_io_pipe_phv_out_data_241; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_242 = pipe9_io_pipe_phv_out_data_242; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_243 = pipe9_io_pipe_phv_out_data_243; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_244 = pipe9_io_pipe_phv_out_data_244; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_245 = pipe9_io_pipe_phv_out_data_245; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_246 = pipe9_io_pipe_phv_out_data_246; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_247 = pipe9_io_pipe_phv_out_data_247; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_248 = pipe9_io_pipe_phv_out_data_248; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_249 = pipe9_io_pipe_phv_out_data_249; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_250 = pipe9_io_pipe_phv_out_data_250; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_251 = pipe9_io_pipe_phv_out_data_251; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_252 = pipe9_io_pipe_phv_out_data_252; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_253 = pipe9_io_pipe_phv_out_data_253; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_254 = pipe9_io_pipe_phv_out_data_254; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_255 = pipe9_io_pipe_phv_out_data_255; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_256 = pipe9_io_pipe_phv_out_data_256; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_257 = pipe9_io_pipe_phv_out_data_257; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_258 = pipe9_io_pipe_phv_out_data_258; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_259 = pipe9_io_pipe_phv_out_data_259; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_260 = pipe9_io_pipe_phv_out_data_260; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_261 = pipe9_io_pipe_phv_out_data_261; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_262 = pipe9_io_pipe_phv_out_data_262; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_263 = pipe9_io_pipe_phv_out_data_263; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_264 = pipe9_io_pipe_phv_out_data_264; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_265 = pipe9_io_pipe_phv_out_data_265; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_266 = pipe9_io_pipe_phv_out_data_266; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_267 = pipe9_io_pipe_phv_out_data_267; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_268 = pipe9_io_pipe_phv_out_data_268; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_269 = pipe9_io_pipe_phv_out_data_269; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_270 = pipe9_io_pipe_phv_out_data_270; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_271 = pipe9_io_pipe_phv_out_data_271; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_272 = pipe9_io_pipe_phv_out_data_272; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_273 = pipe9_io_pipe_phv_out_data_273; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_274 = pipe9_io_pipe_phv_out_data_274; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_275 = pipe9_io_pipe_phv_out_data_275; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_276 = pipe9_io_pipe_phv_out_data_276; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_277 = pipe9_io_pipe_phv_out_data_277; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_278 = pipe9_io_pipe_phv_out_data_278; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_279 = pipe9_io_pipe_phv_out_data_279; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_280 = pipe9_io_pipe_phv_out_data_280; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_281 = pipe9_io_pipe_phv_out_data_281; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_282 = pipe9_io_pipe_phv_out_data_282; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_283 = pipe9_io_pipe_phv_out_data_283; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_284 = pipe9_io_pipe_phv_out_data_284; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_285 = pipe9_io_pipe_phv_out_data_285; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_286 = pipe9_io_pipe_phv_out_data_286; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_287 = pipe9_io_pipe_phv_out_data_287; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_288 = pipe9_io_pipe_phv_out_data_288; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_289 = pipe9_io_pipe_phv_out_data_289; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_290 = pipe9_io_pipe_phv_out_data_290; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_291 = pipe9_io_pipe_phv_out_data_291; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_292 = pipe9_io_pipe_phv_out_data_292; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_293 = pipe9_io_pipe_phv_out_data_293; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_294 = pipe9_io_pipe_phv_out_data_294; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_295 = pipe9_io_pipe_phv_out_data_295; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_296 = pipe9_io_pipe_phv_out_data_296; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_297 = pipe9_io_pipe_phv_out_data_297; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_298 = pipe9_io_pipe_phv_out_data_298; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_299 = pipe9_io_pipe_phv_out_data_299; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_300 = pipe9_io_pipe_phv_out_data_300; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_301 = pipe9_io_pipe_phv_out_data_301; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_302 = pipe9_io_pipe_phv_out_data_302; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_303 = pipe9_io_pipe_phv_out_data_303; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_304 = pipe9_io_pipe_phv_out_data_304; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_305 = pipe9_io_pipe_phv_out_data_305; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_306 = pipe9_io_pipe_phv_out_data_306; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_307 = pipe9_io_pipe_phv_out_data_307; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_308 = pipe9_io_pipe_phv_out_data_308; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_309 = pipe9_io_pipe_phv_out_data_309; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_310 = pipe9_io_pipe_phv_out_data_310; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_311 = pipe9_io_pipe_phv_out_data_311; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_312 = pipe9_io_pipe_phv_out_data_312; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_313 = pipe9_io_pipe_phv_out_data_313; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_314 = pipe9_io_pipe_phv_out_data_314; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_315 = pipe9_io_pipe_phv_out_data_315; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_316 = pipe9_io_pipe_phv_out_data_316; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_317 = pipe9_io_pipe_phv_out_data_317; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_318 = pipe9_io_pipe_phv_out_data_318; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_319 = pipe9_io_pipe_phv_out_data_319; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_320 = pipe9_io_pipe_phv_out_data_320; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_321 = pipe9_io_pipe_phv_out_data_321; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_322 = pipe9_io_pipe_phv_out_data_322; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_323 = pipe9_io_pipe_phv_out_data_323; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_324 = pipe9_io_pipe_phv_out_data_324; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_325 = pipe9_io_pipe_phv_out_data_325; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_326 = pipe9_io_pipe_phv_out_data_326; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_327 = pipe9_io_pipe_phv_out_data_327; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_328 = pipe9_io_pipe_phv_out_data_328; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_329 = pipe9_io_pipe_phv_out_data_329; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_330 = pipe9_io_pipe_phv_out_data_330; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_331 = pipe9_io_pipe_phv_out_data_331; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_332 = pipe9_io_pipe_phv_out_data_332; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_333 = pipe9_io_pipe_phv_out_data_333; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_334 = pipe9_io_pipe_phv_out_data_334; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_335 = pipe9_io_pipe_phv_out_data_335; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_336 = pipe9_io_pipe_phv_out_data_336; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_337 = pipe9_io_pipe_phv_out_data_337; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_338 = pipe9_io_pipe_phv_out_data_338; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_339 = pipe9_io_pipe_phv_out_data_339; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_340 = pipe9_io_pipe_phv_out_data_340; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_341 = pipe9_io_pipe_phv_out_data_341; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_342 = pipe9_io_pipe_phv_out_data_342; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_343 = pipe9_io_pipe_phv_out_data_343; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_344 = pipe9_io_pipe_phv_out_data_344; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_345 = pipe9_io_pipe_phv_out_data_345; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_346 = pipe9_io_pipe_phv_out_data_346; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_347 = pipe9_io_pipe_phv_out_data_347; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_348 = pipe9_io_pipe_phv_out_data_348; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_349 = pipe9_io_pipe_phv_out_data_349; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_350 = pipe9_io_pipe_phv_out_data_350; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_351 = pipe9_io_pipe_phv_out_data_351; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_352 = pipe9_io_pipe_phv_out_data_352; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_353 = pipe9_io_pipe_phv_out_data_353; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_354 = pipe9_io_pipe_phv_out_data_354; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_355 = pipe9_io_pipe_phv_out_data_355; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_356 = pipe9_io_pipe_phv_out_data_356; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_357 = pipe9_io_pipe_phv_out_data_357; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_358 = pipe9_io_pipe_phv_out_data_358; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_359 = pipe9_io_pipe_phv_out_data_359; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_360 = pipe9_io_pipe_phv_out_data_360; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_361 = pipe9_io_pipe_phv_out_data_361; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_362 = pipe9_io_pipe_phv_out_data_362; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_363 = pipe9_io_pipe_phv_out_data_363; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_364 = pipe9_io_pipe_phv_out_data_364; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_365 = pipe9_io_pipe_phv_out_data_365; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_366 = pipe9_io_pipe_phv_out_data_366; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_367 = pipe9_io_pipe_phv_out_data_367; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_368 = pipe9_io_pipe_phv_out_data_368; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_369 = pipe9_io_pipe_phv_out_data_369; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_370 = pipe9_io_pipe_phv_out_data_370; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_371 = pipe9_io_pipe_phv_out_data_371; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_372 = pipe9_io_pipe_phv_out_data_372; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_373 = pipe9_io_pipe_phv_out_data_373; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_374 = pipe9_io_pipe_phv_out_data_374; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_375 = pipe9_io_pipe_phv_out_data_375; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_376 = pipe9_io_pipe_phv_out_data_376; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_377 = pipe9_io_pipe_phv_out_data_377; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_378 = pipe9_io_pipe_phv_out_data_378; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_379 = pipe9_io_pipe_phv_out_data_379; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_380 = pipe9_io_pipe_phv_out_data_380; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_381 = pipe9_io_pipe_phv_out_data_381; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_382 = pipe9_io_pipe_phv_out_data_382; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_383 = pipe9_io_pipe_phv_out_data_383; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_384 = pipe9_io_pipe_phv_out_data_384; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_385 = pipe9_io_pipe_phv_out_data_385; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_386 = pipe9_io_pipe_phv_out_data_386; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_387 = pipe9_io_pipe_phv_out_data_387; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_388 = pipe9_io_pipe_phv_out_data_388; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_389 = pipe9_io_pipe_phv_out_data_389; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_390 = pipe9_io_pipe_phv_out_data_390; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_391 = pipe9_io_pipe_phv_out_data_391; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_392 = pipe9_io_pipe_phv_out_data_392; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_393 = pipe9_io_pipe_phv_out_data_393; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_394 = pipe9_io_pipe_phv_out_data_394; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_395 = pipe9_io_pipe_phv_out_data_395; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_396 = pipe9_io_pipe_phv_out_data_396; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_397 = pipe9_io_pipe_phv_out_data_397; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_398 = pipe9_io_pipe_phv_out_data_398; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_399 = pipe9_io_pipe_phv_out_data_399; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_400 = pipe9_io_pipe_phv_out_data_400; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_401 = pipe9_io_pipe_phv_out_data_401; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_402 = pipe9_io_pipe_phv_out_data_402; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_403 = pipe9_io_pipe_phv_out_data_403; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_404 = pipe9_io_pipe_phv_out_data_404; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_405 = pipe9_io_pipe_phv_out_data_405; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_406 = pipe9_io_pipe_phv_out_data_406; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_407 = pipe9_io_pipe_phv_out_data_407; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_408 = pipe9_io_pipe_phv_out_data_408; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_409 = pipe9_io_pipe_phv_out_data_409; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_410 = pipe9_io_pipe_phv_out_data_410; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_411 = pipe9_io_pipe_phv_out_data_411; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_412 = pipe9_io_pipe_phv_out_data_412; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_413 = pipe9_io_pipe_phv_out_data_413; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_414 = pipe9_io_pipe_phv_out_data_414; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_415 = pipe9_io_pipe_phv_out_data_415; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_416 = pipe9_io_pipe_phv_out_data_416; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_417 = pipe9_io_pipe_phv_out_data_417; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_418 = pipe9_io_pipe_phv_out_data_418; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_419 = pipe9_io_pipe_phv_out_data_419; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_420 = pipe9_io_pipe_phv_out_data_420; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_421 = pipe9_io_pipe_phv_out_data_421; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_422 = pipe9_io_pipe_phv_out_data_422; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_423 = pipe9_io_pipe_phv_out_data_423; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_424 = pipe9_io_pipe_phv_out_data_424; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_425 = pipe9_io_pipe_phv_out_data_425; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_426 = pipe9_io_pipe_phv_out_data_426; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_427 = pipe9_io_pipe_phv_out_data_427; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_428 = pipe9_io_pipe_phv_out_data_428; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_429 = pipe9_io_pipe_phv_out_data_429; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_430 = pipe9_io_pipe_phv_out_data_430; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_431 = pipe9_io_pipe_phv_out_data_431; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_432 = pipe9_io_pipe_phv_out_data_432; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_433 = pipe9_io_pipe_phv_out_data_433; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_434 = pipe9_io_pipe_phv_out_data_434; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_435 = pipe9_io_pipe_phv_out_data_435; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_436 = pipe9_io_pipe_phv_out_data_436; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_437 = pipe9_io_pipe_phv_out_data_437; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_438 = pipe9_io_pipe_phv_out_data_438; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_439 = pipe9_io_pipe_phv_out_data_439; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_440 = pipe9_io_pipe_phv_out_data_440; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_441 = pipe9_io_pipe_phv_out_data_441; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_442 = pipe9_io_pipe_phv_out_data_442; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_443 = pipe9_io_pipe_phv_out_data_443; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_444 = pipe9_io_pipe_phv_out_data_444; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_445 = pipe9_io_pipe_phv_out_data_445; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_446 = pipe9_io_pipe_phv_out_data_446; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_447 = pipe9_io_pipe_phv_out_data_447; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_448 = pipe9_io_pipe_phv_out_data_448; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_449 = pipe9_io_pipe_phv_out_data_449; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_450 = pipe9_io_pipe_phv_out_data_450; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_451 = pipe9_io_pipe_phv_out_data_451; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_452 = pipe9_io_pipe_phv_out_data_452; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_453 = pipe9_io_pipe_phv_out_data_453; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_454 = pipe9_io_pipe_phv_out_data_454; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_455 = pipe9_io_pipe_phv_out_data_455; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_456 = pipe9_io_pipe_phv_out_data_456; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_457 = pipe9_io_pipe_phv_out_data_457; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_458 = pipe9_io_pipe_phv_out_data_458; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_459 = pipe9_io_pipe_phv_out_data_459; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_460 = pipe9_io_pipe_phv_out_data_460; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_461 = pipe9_io_pipe_phv_out_data_461; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_462 = pipe9_io_pipe_phv_out_data_462; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_463 = pipe9_io_pipe_phv_out_data_463; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_464 = pipe9_io_pipe_phv_out_data_464; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_465 = pipe9_io_pipe_phv_out_data_465; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_466 = pipe9_io_pipe_phv_out_data_466; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_467 = pipe9_io_pipe_phv_out_data_467; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_468 = pipe9_io_pipe_phv_out_data_468; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_469 = pipe9_io_pipe_phv_out_data_469; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_470 = pipe9_io_pipe_phv_out_data_470; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_471 = pipe9_io_pipe_phv_out_data_471; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_472 = pipe9_io_pipe_phv_out_data_472; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_473 = pipe9_io_pipe_phv_out_data_473; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_474 = pipe9_io_pipe_phv_out_data_474; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_475 = pipe9_io_pipe_phv_out_data_475; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_476 = pipe9_io_pipe_phv_out_data_476; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_477 = pipe9_io_pipe_phv_out_data_477; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_478 = pipe9_io_pipe_phv_out_data_478; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_479 = pipe9_io_pipe_phv_out_data_479; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_480 = pipe9_io_pipe_phv_out_data_480; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_481 = pipe9_io_pipe_phv_out_data_481; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_482 = pipe9_io_pipe_phv_out_data_482; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_483 = pipe9_io_pipe_phv_out_data_483; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_484 = pipe9_io_pipe_phv_out_data_484; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_485 = pipe9_io_pipe_phv_out_data_485; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_486 = pipe9_io_pipe_phv_out_data_486; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_487 = pipe9_io_pipe_phv_out_data_487; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_488 = pipe9_io_pipe_phv_out_data_488; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_489 = pipe9_io_pipe_phv_out_data_489; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_490 = pipe9_io_pipe_phv_out_data_490; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_491 = pipe9_io_pipe_phv_out_data_491; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_492 = pipe9_io_pipe_phv_out_data_492; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_493 = pipe9_io_pipe_phv_out_data_493; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_494 = pipe9_io_pipe_phv_out_data_494; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_495 = pipe9_io_pipe_phv_out_data_495; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_496 = pipe9_io_pipe_phv_out_data_496; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_497 = pipe9_io_pipe_phv_out_data_497; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_498 = pipe9_io_pipe_phv_out_data_498; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_499 = pipe9_io_pipe_phv_out_data_499; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_500 = pipe9_io_pipe_phv_out_data_500; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_501 = pipe9_io_pipe_phv_out_data_501; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_502 = pipe9_io_pipe_phv_out_data_502; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_503 = pipe9_io_pipe_phv_out_data_503; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_504 = pipe9_io_pipe_phv_out_data_504; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_505 = pipe9_io_pipe_phv_out_data_505; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_506 = pipe9_io_pipe_phv_out_data_506; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_507 = pipe9_io_pipe_phv_out_data_507; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_508 = pipe9_io_pipe_phv_out_data_508; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_509 = pipe9_io_pipe_phv_out_data_509; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_510 = pipe9_io_pipe_phv_out_data_510; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_511 = pipe9_io_pipe_phv_out_data_511; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_0 = pipe9_io_pipe_phv_out_header_0; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_1 = pipe9_io_pipe_phv_out_header_1; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_2 = pipe9_io_pipe_phv_out_header_2; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_3 = pipe9_io_pipe_phv_out_header_3; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_4 = pipe9_io_pipe_phv_out_header_4; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_5 = pipe9_io_pipe_phv_out_header_5; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_6 = pipe9_io_pipe_phv_out_header_6; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_7 = pipe9_io_pipe_phv_out_header_7; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_8 = pipe9_io_pipe_phv_out_header_8; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_9 = pipe9_io_pipe_phv_out_header_9; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_10 = pipe9_io_pipe_phv_out_header_10; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_11 = pipe9_io_pipe_phv_out_header_11; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_12 = pipe9_io_pipe_phv_out_header_12; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_13 = pipe9_io_pipe_phv_out_header_13; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_14 = pipe9_io_pipe_phv_out_header_14; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_15 = pipe9_io_pipe_phv_out_header_15; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_parse_current_state = pipe9_io_pipe_phv_out_parse_current_state; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_parse_current_offset = pipe9_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_parse_transition_field = pipe9_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_next_processor_id = pipe9_io_pipe_phv_out_next_processor_id; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_next_config_id = pipe9_io_pipe_phv_out_next_config_id; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_is_valid_processor = pipe9_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 370:27]
  assign pipe10_io_key_in = pipe9_io_key_out; // @[matcher.scala 371:27]
  assign pipe10_io_cs_in = pipe9_io_cs_out; // @[matcher.scala 372:27]
  assign pipe10_io_addr_in = pipe9_io_addr_out; // @[matcher.scala 373:27]
  assign pipe10_io_cs_vec_in_0 = pipe9_io_cs_vec_out_0; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_1 = pipe9_io_cs_vec_out_1; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_2 = pipe9_io_cs_vec_out_2; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_3 = pipe9_io_cs_vec_out_3; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_4 = pipe9_io_cs_vec_out_4; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_5 = pipe9_io_cs_vec_out_5; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_6 = pipe9_io_cs_vec_out_6; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_7 = pipe9_io_cs_vec_out_7; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_8 = pipe9_io_cs_vec_out_8; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_9 = pipe9_io_cs_vec_out_9; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_10 = pipe9_io_cs_vec_out_10; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_11 = pipe9_io_cs_vec_out_11; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_12 = pipe9_io_cs_vec_out_12; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_13 = pipe9_io_cs_vec_out_13; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_14 = pipe9_io_cs_vec_out_14; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_15 = pipe9_io_cs_vec_out_15; // @[matcher.scala 374:27]
  assign pipe10_io_mem_cluster_0_data = io_mem_cluster_0_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_1_data = io_mem_cluster_1_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_2_data = io_mem_cluster_2_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_3_data = io_mem_cluster_3_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_4_data = io_mem_cluster_4_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_5_data = io_mem_cluster_5_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_6_data = io_mem_cluster_6_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_7_data = io_mem_cluster_7_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_8_data = io_mem_cluster_8_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_9_data = io_mem_cluster_9_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_10_data = io_mem_cluster_10_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_11_data = io_mem_cluster_11_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_12_data = io_mem_cluster_12_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_13_data = io_mem_cluster_13_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_14_data = io_mem_cluster_14_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_15_data = io_mem_cluster_15_data; // @[matcher.scala 375:27]
  assign pipe11_clock = clock;
  assign pipe11_io_pipe_phv_in_data_0 = pipe10_io_pipe_phv_out_data_0; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_1 = pipe10_io_pipe_phv_out_data_1; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_2 = pipe10_io_pipe_phv_out_data_2; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_3 = pipe10_io_pipe_phv_out_data_3; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_4 = pipe10_io_pipe_phv_out_data_4; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_5 = pipe10_io_pipe_phv_out_data_5; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_6 = pipe10_io_pipe_phv_out_data_6; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_7 = pipe10_io_pipe_phv_out_data_7; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_8 = pipe10_io_pipe_phv_out_data_8; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_9 = pipe10_io_pipe_phv_out_data_9; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_10 = pipe10_io_pipe_phv_out_data_10; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_11 = pipe10_io_pipe_phv_out_data_11; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_12 = pipe10_io_pipe_phv_out_data_12; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_13 = pipe10_io_pipe_phv_out_data_13; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_14 = pipe10_io_pipe_phv_out_data_14; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_15 = pipe10_io_pipe_phv_out_data_15; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_16 = pipe10_io_pipe_phv_out_data_16; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_17 = pipe10_io_pipe_phv_out_data_17; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_18 = pipe10_io_pipe_phv_out_data_18; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_19 = pipe10_io_pipe_phv_out_data_19; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_20 = pipe10_io_pipe_phv_out_data_20; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_21 = pipe10_io_pipe_phv_out_data_21; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_22 = pipe10_io_pipe_phv_out_data_22; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_23 = pipe10_io_pipe_phv_out_data_23; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_24 = pipe10_io_pipe_phv_out_data_24; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_25 = pipe10_io_pipe_phv_out_data_25; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_26 = pipe10_io_pipe_phv_out_data_26; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_27 = pipe10_io_pipe_phv_out_data_27; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_28 = pipe10_io_pipe_phv_out_data_28; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_29 = pipe10_io_pipe_phv_out_data_29; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_30 = pipe10_io_pipe_phv_out_data_30; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_31 = pipe10_io_pipe_phv_out_data_31; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_32 = pipe10_io_pipe_phv_out_data_32; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_33 = pipe10_io_pipe_phv_out_data_33; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_34 = pipe10_io_pipe_phv_out_data_34; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_35 = pipe10_io_pipe_phv_out_data_35; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_36 = pipe10_io_pipe_phv_out_data_36; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_37 = pipe10_io_pipe_phv_out_data_37; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_38 = pipe10_io_pipe_phv_out_data_38; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_39 = pipe10_io_pipe_phv_out_data_39; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_40 = pipe10_io_pipe_phv_out_data_40; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_41 = pipe10_io_pipe_phv_out_data_41; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_42 = pipe10_io_pipe_phv_out_data_42; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_43 = pipe10_io_pipe_phv_out_data_43; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_44 = pipe10_io_pipe_phv_out_data_44; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_45 = pipe10_io_pipe_phv_out_data_45; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_46 = pipe10_io_pipe_phv_out_data_46; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_47 = pipe10_io_pipe_phv_out_data_47; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_48 = pipe10_io_pipe_phv_out_data_48; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_49 = pipe10_io_pipe_phv_out_data_49; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_50 = pipe10_io_pipe_phv_out_data_50; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_51 = pipe10_io_pipe_phv_out_data_51; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_52 = pipe10_io_pipe_phv_out_data_52; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_53 = pipe10_io_pipe_phv_out_data_53; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_54 = pipe10_io_pipe_phv_out_data_54; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_55 = pipe10_io_pipe_phv_out_data_55; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_56 = pipe10_io_pipe_phv_out_data_56; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_57 = pipe10_io_pipe_phv_out_data_57; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_58 = pipe10_io_pipe_phv_out_data_58; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_59 = pipe10_io_pipe_phv_out_data_59; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_60 = pipe10_io_pipe_phv_out_data_60; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_61 = pipe10_io_pipe_phv_out_data_61; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_62 = pipe10_io_pipe_phv_out_data_62; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_63 = pipe10_io_pipe_phv_out_data_63; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_64 = pipe10_io_pipe_phv_out_data_64; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_65 = pipe10_io_pipe_phv_out_data_65; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_66 = pipe10_io_pipe_phv_out_data_66; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_67 = pipe10_io_pipe_phv_out_data_67; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_68 = pipe10_io_pipe_phv_out_data_68; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_69 = pipe10_io_pipe_phv_out_data_69; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_70 = pipe10_io_pipe_phv_out_data_70; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_71 = pipe10_io_pipe_phv_out_data_71; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_72 = pipe10_io_pipe_phv_out_data_72; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_73 = pipe10_io_pipe_phv_out_data_73; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_74 = pipe10_io_pipe_phv_out_data_74; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_75 = pipe10_io_pipe_phv_out_data_75; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_76 = pipe10_io_pipe_phv_out_data_76; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_77 = pipe10_io_pipe_phv_out_data_77; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_78 = pipe10_io_pipe_phv_out_data_78; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_79 = pipe10_io_pipe_phv_out_data_79; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_80 = pipe10_io_pipe_phv_out_data_80; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_81 = pipe10_io_pipe_phv_out_data_81; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_82 = pipe10_io_pipe_phv_out_data_82; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_83 = pipe10_io_pipe_phv_out_data_83; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_84 = pipe10_io_pipe_phv_out_data_84; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_85 = pipe10_io_pipe_phv_out_data_85; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_86 = pipe10_io_pipe_phv_out_data_86; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_87 = pipe10_io_pipe_phv_out_data_87; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_88 = pipe10_io_pipe_phv_out_data_88; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_89 = pipe10_io_pipe_phv_out_data_89; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_90 = pipe10_io_pipe_phv_out_data_90; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_91 = pipe10_io_pipe_phv_out_data_91; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_92 = pipe10_io_pipe_phv_out_data_92; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_93 = pipe10_io_pipe_phv_out_data_93; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_94 = pipe10_io_pipe_phv_out_data_94; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_95 = pipe10_io_pipe_phv_out_data_95; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_96 = pipe10_io_pipe_phv_out_data_96; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_97 = pipe10_io_pipe_phv_out_data_97; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_98 = pipe10_io_pipe_phv_out_data_98; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_99 = pipe10_io_pipe_phv_out_data_99; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_100 = pipe10_io_pipe_phv_out_data_100; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_101 = pipe10_io_pipe_phv_out_data_101; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_102 = pipe10_io_pipe_phv_out_data_102; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_103 = pipe10_io_pipe_phv_out_data_103; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_104 = pipe10_io_pipe_phv_out_data_104; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_105 = pipe10_io_pipe_phv_out_data_105; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_106 = pipe10_io_pipe_phv_out_data_106; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_107 = pipe10_io_pipe_phv_out_data_107; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_108 = pipe10_io_pipe_phv_out_data_108; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_109 = pipe10_io_pipe_phv_out_data_109; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_110 = pipe10_io_pipe_phv_out_data_110; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_111 = pipe10_io_pipe_phv_out_data_111; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_112 = pipe10_io_pipe_phv_out_data_112; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_113 = pipe10_io_pipe_phv_out_data_113; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_114 = pipe10_io_pipe_phv_out_data_114; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_115 = pipe10_io_pipe_phv_out_data_115; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_116 = pipe10_io_pipe_phv_out_data_116; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_117 = pipe10_io_pipe_phv_out_data_117; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_118 = pipe10_io_pipe_phv_out_data_118; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_119 = pipe10_io_pipe_phv_out_data_119; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_120 = pipe10_io_pipe_phv_out_data_120; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_121 = pipe10_io_pipe_phv_out_data_121; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_122 = pipe10_io_pipe_phv_out_data_122; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_123 = pipe10_io_pipe_phv_out_data_123; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_124 = pipe10_io_pipe_phv_out_data_124; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_125 = pipe10_io_pipe_phv_out_data_125; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_126 = pipe10_io_pipe_phv_out_data_126; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_127 = pipe10_io_pipe_phv_out_data_127; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_128 = pipe10_io_pipe_phv_out_data_128; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_129 = pipe10_io_pipe_phv_out_data_129; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_130 = pipe10_io_pipe_phv_out_data_130; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_131 = pipe10_io_pipe_phv_out_data_131; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_132 = pipe10_io_pipe_phv_out_data_132; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_133 = pipe10_io_pipe_phv_out_data_133; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_134 = pipe10_io_pipe_phv_out_data_134; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_135 = pipe10_io_pipe_phv_out_data_135; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_136 = pipe10_io_pipe_phv_out_data_136; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_137 = pipe10_io_pipe_phv_out_data_137; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_138 = pipe10_io_pipe_phv_out_data_138; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_139 = pipe10_io_pipe_phv_out_data_139; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_140 = pipe10_io_pipe_phv_out_data_140; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_141 = pipe10_io_pipe_phv_out_data_141; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_142 = pipe10_io_pipe_phv_out_data_142; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_143 = pipe10_io_pipe_phv_out_data_143; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_144 = pipe10_io_pipe_phv_out_data_144; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_145 = pipe10_io_pipe_phv_out_data_145; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_146 = pipe10_io_pipe_phv_out_data_146; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_147 = pipe10_io_pipe_phv_out_data_147; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_148 = pipe10_io_pipe_phv_out_data_148; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_149 = pipe10_io_pipe_phv_out_data_149; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_150 = pipe10_io_pipe_phv_out_data_150; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_151 = pipe10_io_pipe_phv_out_data_151; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_152 = pipe10_io_pipe_phv_out_data_152; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_153 = pipe10_io_pipe_phv_out_data_153; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_154 = pipe10_io_pipe_phv_out_data_154; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_155 = pipe10_io_pipe_phv_out_data_155; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_156 = pipe10_io_pipe_phv_out_data_156; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_157 = pipe10_io_pipe_phv_out_data_157; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_158 = pipe10_io_pipe_phv_out_data_158; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_159 = pipe10_io_pipe_phv_out_data_159; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_160 = pipe10_io_pipe_phv_out_data_160; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_161 = pipe10_io_pipe_phv_out_data_161; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_162 = pipe10_io_pipe_phv_out_data_162; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_163 = pipe10_io_pipe_phv_out_data_163; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_164 = pipe10_io_pipe_phv_out_data_164; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_165 = pipe10_io_pipe_phv_out_data_165; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_166 = pipe10_io_pipe_phv_out_data_166; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_167 = pipe10_io_pipe_phv_out_data_167; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_168 = pipe10_io_pipe_phv_out_data_168; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_169 = pipe10_io_pipe_phv_out_data_169; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_170 = pipe10_io_pipe_phv_out_data_170; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_171 = pipe10_io_pipe_phv_out_data_171; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_172 = pipe10_io_pipe_phv_out_data_172; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_173 = pipe10_io_pipe_phv_out_data_173; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_174 = pipe10_io_pipe_phv_out_data_174; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_175 = pipe10_io_pipe_phv_out_data_175; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_176 = pipe10_io_pipe_phv_out_data_176; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_177 = pipe10_io_pipe_phv_out_data_177; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_178 = pipe10_io_pipe_phv_out_data_178; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_179 = pipe10_io_pipe_phv_out_data_179; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_180 = pipe10_io_pipe_phv_out_data_180; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_181 = pipe10_io_pipe_phv_out_data_181; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_182 = pipe10_io_pipe_phv_out_data_182; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_183 = pipe10_io_pipe_phv_out_data_183; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_184 = pipe10_io_pipe_phv_out_data_184; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_185 = pipe10_io_pipe_phv_out_data_185; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_186 = pipe10_io_pipe_phv_out_data_186; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_187 = pipe10_io_pipe_phv_out_data_187; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_188 = pipe10_io_pipe_phv_out_data_188; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_189 = pipe10_io_pipe_phv_out_data_189; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_190 = pipe10_io_pipe_phv_out_data_190; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_191 = pipe10_io_pipe_phv_out_data_191; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_192 = pipe10_io_pipe_phv_out_data_192; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_193 = pipe10_io_pipe_phv_out_data_193; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_194 = pipe10_io_pipe_phv_out_data_194; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_195 = pipe10_io_pipe_phv_out_data_195; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_196 = pipe10_io_pipe_phv_out_data_196; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_197 = pipe10_io_pipe_phv_out_data_197; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_198 = pipe10_io_pipe_phv_out_data_198; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_199 = pipe10_io_pipe_phv_out_data_199; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_200 = pipe10_io_pipe_phv_out_data_200; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_201 = pipe10_io_pipe_phv_out_data_201; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_202 = pipe10_io_pipe_phv_out_data_202; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_203 = pipe10_io_pipe_phv_out_data_203; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_204 = pipe10_io_pipe_phv_out_data_204; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_205 = pipe10_io_pipe_phv_out_data_205; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_206 = pipe10_io_pipe_phv_out_data_206; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_207 = pipe10_io_pipe_phv_out_data_207; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_208 = pipe10_io_pipe_phv_out_data_208; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_209 = pipe10_io_pipe_phv_out_data_209; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_210 = pipe10_io_pipe_phv_out_data_210; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_211 = pipe10_io_pipe_phv_out_data_211; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_212 = pipe10_io_pipe_phv_out_data_212; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_213 = pipe10_io_pipe_phv_out_data_213; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_214 = pipe10_io_pipe_phv_out_data_214; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_215 = pipe10_io_pipe_phv_out_data_215; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_216 = pipe10_io_pipe_phv_out_data_216; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_217 = pipe10_io_pipe_phv_out_data_217; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_218 = pipe10_io_pipe_phv_out_data_218; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_219 = pipe10_io_pipe_phv_out_data_219; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_220 = pipe10_io_pipe_phv_out_data_220; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_221 = pipe10_io_pipe_phv_out_data_221; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_222 = pipe10_io_pipe_phv_out_data_222; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_223 = pipe10_io_pipe_phv_out_data_223; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_224 = pipe10_io_pipe_phv_out_data_224; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_225 = pipe10_io_pipe_phv_out_data_225; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_226 = pipe10_io_pipe_phv_out_data_226; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_227 = pipe10_io_pipe_phv_out_data_227; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_228 = pipe10_io_pipe_phv_out_data_228; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_229 = pipe10_io_pipe_phv_out_data_229; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_230 = pipe10_io_pipe_phv_out_data_230; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_231 = pipe10_io_pipe_phv_out_data_231; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_232 = pipe10_io_pipe_phv_out_data_232; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_233 = pipe10_io_pipe_phv_out_data_233; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_234 = pipe10_io_pipe_phv_out_data_234; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_235 = pipe10_io_pipe_phv_out_data_235; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_236 = pipe10_io_pipe_phv_out_data_236; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_237 = pipe10_io_pipe_phv_out_data_237; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_238 = pipe10_io_pipe_phv_out_data_238; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_239 = pipe10_io_pipe_phv_out_data_239; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_240 = pipe10_io_pipe_phv_out_data_240; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_241 = pipe10_io_pipe_phv_out_data_241; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_242 = pipe10_io_pipe_phv_out_data_242; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_243 = pipe10_io_pipe_phv_out_data_243; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_244 = pipe10_io_pipe_phv_out_data_244; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_245 = pipe10_io_pipe_phv_out_data_245; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_246 = pipe10_io_pipe_phv_out_data_246; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_247 = pipe10_io_pipe_phv_out_data_247; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_248 = pipe10_io_pipe_phv_out_data_248; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_249 = pipe10_io_pipe_phv_out_data_249; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_250 = pipe10_io_pipe_phv_out_data_250; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_251 = pipe10_io_pipe_phv_out_data_251; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_252 = pipe10_io_pipe_phv_out_data_252; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_253 = pipe10_io_pipe_phv_out_data_253; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_254 = pipe10_io_pipe_phv_out_data_254; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_255 = pipe10_io_pipe_phv_out_data_255; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_256 = pipe10_io_pipe_phv_out_data_256; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_257 = pipe10_io_pipe_phv_out_data_257; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_258 = pipe10_io_pipe_phv_out_data_258; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_259 = pipe10_io_pipe_phv_out_data_259; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_260 = pipe10_io_pipe_phv_out_data_260; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_261 = pipe10_io_pipe_phv_out_data_261; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_262 = pipe10_io_pipe_phv_out_data_262; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_263 = pipe10_io_pipe_phv_out_data_263; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_264 = pipe10_io_pipe_phv_out_data_264; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_265 = pipe10_io_pipe_phv_out_data_265; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_266 = pipe10_io_pipe_phv_out_data_266; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_267 = pipe10_io_pipe_phv_out_data_267; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_268 = pipe10_io_pipe_phv_out_data_268; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_269 = pipe10_io_pipe_phv_out_data_269; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_270 = pipe10_io_pipe_phv_out_data_270; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_271 = pipe10_io_pipe_phv_out_data_271; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_272 = pipe10_io_pipe_phv_out_data_272; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_273 = pipe10_io_pipe_phv_out_data_273; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_274 = pipe10_io_pipe_phv_out_data_274; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_275 = pipe10_io_pipe_phv_out_data_275; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_276 = pipe10_io_pipe_phv_out_data_276; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_277 = pipe10_io_pipe_phv_out_data_277; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_278 = pipe10_io_pipe_phv_out_data_278; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_279 = pipe10_io_pipe_phv_out_data_279; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_280 = pipe10_io_pipe_phv_out_data_280; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_281 = pipe10_io_pipe_phv_out_data_281; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_282 = pipe10_io_pipe_phv_out_data_282; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_283 = pipe10_io_pipe_phv_out_data_283; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_284 = pipe10_io_pipe_phv_out_data_284; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_285 = pipe10_io_pipe_phv_out_data_285; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_286 = pipe10_io_pipe_phv_out_data_286; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_287 = pipe10_io_pipe_phv_out_data_287; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_288 = pipe10_io_pipe_phv_out_data_288; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_289 = pipe10_io_pipe_phv_out_data_289; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_290 = pipe10_io_pipe_phv_out_data_290; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_291 = pipe10_io_pipe_phv_out_data_291; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_292 = pipe10_io_pipe_phv_out_data_292; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_293 = pipe10_io_pipe_phv_out_data_293; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_294 = pipe10_io_pipe_phv_out_data_294; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_295 = pipe10_io_pipe_phv_out_data_295; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_296 = pipe10_io_pipe_phv_out_data_296; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_297 = pipe10_io_pipe_phv_out_data_297; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_298 = pipe10_io_pipe_phv_out_data_298; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_299 = pipe10_io_pipe_phv_out_data_299; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_300 = pipe10_io_pipe_phv_out_data_300; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_301 = pipe10_io_pipe_phv_out_data_301; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_302 = pipe10_io_pipe_phv_out_data_302; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_303 = pipe10_io_pipe_phv_out_data_303; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_304 = pipe10_io_pipe_phv_out_data_304; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_305 = pipe10_io_pipe_phv_out_data_305; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_306 = pipe10_io_pipe_phv_out_data_306; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_307 = pipe10_io_pipe_phv_out_data_307; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_308 = pipe10_io_pipe_phv_out_data_308; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_309 = pipe10_io_pipe_phv_out_data_309; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_310 = pipe10_io_pipe_phv_out_data_310; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_311 = pipe10_io_pipe_phv_out_data_311; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_312 = pipe10_io_pipe_phv_out_data_312; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_313 = pipe10_io_pipe_phv_out_data_313; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_314 = pipe10_io_pipe_phv_out_data_314; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_315 = pipe10_io_pipe_phv_out_data_315; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_316 = pipe10_io_pipe_phv_out_data_316; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_317 = pipe10_io_pipe_phv_out_data_317; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_318 = pipe10_io_pipe_phv_out_data_318; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_319 = pipe10_io_pipe_phv_out_data_319; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_320 = pipe10_io_pipe_phv_out_data_320; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_321 = pipe10_io_pipe_phv_out_data_321; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_322 = pipe10_io_pipe_phv_out_data_322; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_323 = pipe10_io_pipe_phv_out_data_323; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_324 = pipe10_io_pipe_phv_out_data_324; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_325 = pipe10_io_pipe_phv_out_data_325; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_326 = pipe10_io_pipe_phv_out_data_326; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_327 = pipe10_io_pipe_phv_out_data_327; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_328 = pipe10_io_pipe_phv_out_data_328; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_329 = pipe10_io_pipe_phv_out_data_329; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_330 = pipe10_io_pipe_phv_out_data_330; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_331 = pipe10_io_pipe_phv_out_data_331; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_332 = pipe10_io_pipe_phv_out_data_332; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_333 = pipe10_io_pipe_phv_out_data_333; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_334 = pipe10_io_pipe_phv_out_data_334; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_335 = pipe10_io_pipe_phv_out_data_335; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_336 = pipe10_io_pipe_phv_out_data_336; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_337 = pipe10_io_pipe_phv_out_data_337; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_338 = pipe10_io_pipe_phv_out_data_338; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_339 = pipe10_io_pipe_phv_out_data_339; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_340 = pipe10_io_pipe_phv_out_data_340; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_341 = pipe10_io_pipe_phv_out_data_341; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_342 = pipe10_io_pipe_phv_out_data_342; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_343 = pipe10_io_pipe_phv_out_data_343; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_344 = pipe10_io_pipe_phv_out_data_344; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_345 = pipe10_io_pipe_phv_out_data_345; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_346 = pipe10_io_pipe_phv_out_data_346; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_347 = pipe10_io_pipe_phv_out_data_347; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_348 = pipe10_io_pipe_phv_out_data_348; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_349 = pipe10_io_pipe_phv_out_data_349; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_350 = pipe10_io_pipe_phv_out_data_350; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_351 = pipe10_io_pipe_phv_out_data_351; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_352 = pipe10_io_pipe_phv_out_data_352; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_353 = pipe10_io_pipe_phv_out_data_353; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_354 = pipe10_io_pipe_phv_out_data_354; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_355 = pipe10_io_pipe_phv_out_data_355; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_356 = pipe10_io_pipe_phv_out_data_356; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_357 = pipe10_io_pipe_phv_out_data_357; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_358 = pipe10_io_pipe_phv_out_data_358; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_359 = pipe10_io_pipe_phv_out_data_359; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_360 = pipe10_io_pipe_phv_out_data_360; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_361 = pipe10_io_pipe_phv_out_data_361; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_362 = pipe10_io_pipe_phv_out_data_362; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_363 = pipe10_io_pipe_phv_out_data_363; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_364 = pipe10_io_pipe_phv_out_data_364; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_365 = pipe10_io_pipe_phv_out_data_365; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_366 = pipe10_io_pipe_phv_out_data_366; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_367 = pipe10_io_pipe_phv_out_data_367; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_368 = pipe10_io_pipe_phv_out_data_368; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_369 = pipe10_io_pipe_phv_out_data_369; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_370 = pipe10_io_pipe_phv_out_data_370; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_371 = pipe10_io_pipe_phv_out_data_371; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_372 = pipe10_io_pipe_phv_out_data_372; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_373 = pipe10_io_pipe_phv_out_data_373; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_374 = pipe10_io_pipe_phv_out_data_374; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_375 = pipe10_io_pipe_phv_out_data_375; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_376 = pipe10_io_pipe_phv_out_data_376; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_377 = pipe10_io_pipe_phv_out_data_377; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_378 = pipe10_io_pipe_phv_out_data_378; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_379 = pipe10_io_pipe_phv_out_data_379; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_380 = pipe10_io_pipe_phv_out_data_380; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_381 = pipe10_io_pipe_phv_out_data_381; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_382 = pipe10_io_pipe_phv_out_data_382; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_383 = pipe10_io_pipe_phv_out_data_383; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_384 = pipe10_io_pipe_phv_out_data_384; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_385 = pipe10_io_pipe_phv_out_data_385; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_386 = pipe10_io_pipe_phv_out_data_386; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_387 = pipe10_io_pipe_phv_out_data_387; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_388 = pipe10_io_pipe_phv_out_data_388; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_389 = pipe10_io_pipe_phv_out_data_389; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_390 = pipe10_io_pipe_phv_out_data_390; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_391 = pipe10_io_pipe_phv_out_data_391; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_392 = pipe10_io_pipe_phv_out_data_392; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_393 = pipe10_io_pipe_phv_out_data_393; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_394 = pipe10_io_pipe_phv_out_data_394; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_395 = pipe10_io_pipe_phv_out_data_395; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_396 = pipe10_io_pipe_phv_out_data_396; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_397 = pipe10_io_pipe_phv_out_data_397; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_398 = pipe10_io_pipe_phv_out_data_398; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_399 = pipe10_io_pipe_phv_out_data_399; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_400 = pipe10_io_pipe_phv_out_data_400; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_401 = pipe10_io_pipe_phv_out_data_401; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_402 = pipe10_io_pipe_phv_out_data_402; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_403 = pipe10_io_pipe_phv_out_data_403; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_404 = pipe10_io_pipe_phv_out_data_404; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_405 = pipe10_io_pipe_phv_out_data_405; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_406 = pipe10_io_pipe_phv_out_data_406; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_407 = pipe10_io_pipe_phv_out_data_407; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_408 = pipe10_io_pipe_phv_out_data_408; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_409 = pipe10_io_pipe_phv_out_data_409; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_410 = pipe10_io_pipe_phv_out_data_410; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_411 = pipe10_io_pipe_phv_out_data_411; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_412 = pipe10_io_pipe_phv_out_data_412; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_413 = pipe10_io_pipe_phv_out_data_413; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_414 = pipe10_io_pipe_phv_out_data_414; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_415 = pipe10_io_pipe_phv_out_data_415; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_416 = pipe10_io_pipe_phv_out_data_416; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_417 = pipe10_io_pipe_phv_out_data_417; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_418 = pipe10_io_pipe_phv_out_data_418; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_419 = pipe10_io_pipe_phv_out_data_419; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_420 = pipe10_io_pipe_phv_out_data_420; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_421 = pipe10_io_pipe_phv_out_data_421; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_422 = pipe10_io_pipe_phv_out_data_422; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_423 = pipe10_io_pipe_phv_out_data_423; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_424 = pipe10_io_pipe_phv_out_data_424; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_425 = pipe10_io_pipe_phv_out_data_425; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_426 = pipe10_io_pipe_phv_out_data_426; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_427 = pipe10_io_pipe_phv_out_data_427; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_428 = pipe10_io_pipe_phv_out_data_428; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_429 = pipe10_io_pipe_phv_out_data_429; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_430 = pipe10_io_pipe_phv_out_data_430; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_431 = pipe10_io_pipe_phv_out_data_431; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_432 = pipe10_io_pipe_phv_out_data_432; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_433 = pipe10_io_pipe_phv_out_data_433; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_434 = pipe10_io_pipe_phv_out_data_434; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_435 = pipe10_io_pipe_phv_out_data_435; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_436 = pipe10_io_pipe_phv_out_data_436; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_437 = pipe10_io_pipe_phv_out_data_437; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_438 = pipe10_io_pipe_phv_out_data_438; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_439 = pipe10_io_pipe_phv_out_data_439; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_440 = pipe10_io_pipe_phv_out_data_440; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_441 = pipe10_io_pipe_phv_out_data_441; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_442 = pipe10_io_pipe_phv_out_data_442; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_443 = pipe10_io_pipe_phv_out_data_443; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_444 = pipe10_io_pipe_phv_out_data_444; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_445 = pipe10_io_pipe_phv_out_data_445; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_446 = pipe10_io_pipe_phv_out_data_446; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_447 = pipe10_io_pipe_phv_out_data_447; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_448 = pipe10_io_pipe_phv_out_data_448; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_449 = pipe10_io_pipe_phv_out_data_449; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_450 = pipe10_io_pipe_phv_out_data_450; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_451 = pipe10_io_pipe_phv_out_data_451; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_452 = pipe10_io_pipe_phv_out_data_452; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_453 = pipe10_io_pipe_phv_out_data_453; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_454 = pipe10_io_pipe_phv_out_data_454; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_455 = pipe10_io_pipe_phv_out_data_455; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_456 = pipe10_io_pipe_phv_out_data_456; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_457 = pipe10_io_pipe_phv_out_data_457; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_458 = pipe10_io_pipe_phv_out_data_458; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_459 = pipe10_io_pipe_phv_out_data_459; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_460 = pipe10_io_pipe_phv_out_data_460; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_461 = pipe10_io_pipe_phv_out_data_461; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_462 = pipe10_io_pipe_phv_out_data_462; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_463 = pipe10_io_pipe_phv_out_data_463; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_464 = pipe10_io_pipe_phv_out_data_464; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_465 = pipe10_io_pipe_phv_out_data_465; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_466 = pipe10_io_pipe_phv_out_data_466; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_467 = pipe10_io_pipe_phv_out_data_467; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_468 = pipe10_io_pipe_phv_out_data_468; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_469 = pipe10_io_pipe_phv_out_data_469; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_470 = pipe10_io_pipe_phv_out_data_470; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_471 = pipe10_io_pipe_phv_out_data_471; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_472 = pipe10_io_pipe_phv_out_data_472; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_473 = pipe10_io_pipe_phv_out_data_473; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_474 = pipe10_io_pipe_phv_out_data_474; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_475 = pipe10_io_pipe_phv_out_data_475; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_476 = pipe10_io_pipe_phv_out_data_476; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_477 = pipe10_io_pipe_phv_out_data_477; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_478 = pipe10_io_pipe_phv_out_data_478; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_479 = pipe10_io_pipe_phv_out_data_479; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_480 = pipe10_io_pipe_phv_out_data_480; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_481 = pipe10_io_pipe_phv_out_data_481; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_482 = pipe10_io_pipe_phv_out_data_482; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_483 = pipe10_io_pipe_phv_out_data_483; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_484 = pipe10_io_pipe_phv_out_data_484; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_485 = pipe10_io_pipe_phv_out_data_485; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_486 = pipe10_io_pipe_phv_out_data_486; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_487 = pipe10_io_pipe_phv_out_data_487; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_488 = pipe10_io_pipe_phv_out_data_488; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_489 = pipe10_io_pipe_phv_out_data_489; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_490 = pipe10_io_pipe_phv_out_data_490; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_491 = pipe10_io_pipe_phv_out_data_491; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_492 = pipe10_io_pipe_phv_out_data_492; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_493 = pipe10_io_pipe_phv_out_data_493; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_494 = pipe10_io_pipe_phv_out_data_494; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_495 = pipe10_io_pipe_phv_out_data_495; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_496 = pipe10_io_pipe_phv_out_data_496; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_497 = pipe10_io_pipe_phv_out_data_497; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_498 = pipe10_io_pipe_phv_out_data_498; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_499 = pipe10_io_pipe_phv_out_data_499; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_500 = pipe10_io_pipe_phv_out_data_500; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_501 = pipe10_io_pipe_phv_out_data_501; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_502 = pipe10_io_pipe_phv_out_data_502; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_503 = pipe10_io_pipe_phv_out_data_503; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_504 = pipe10_io_pipe_phv_out_data_504; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_505 = pipe10_io_pipe_phv_out_data_505; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_506 = pipe10_io_pipe_phv_out_data_506; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_507 = pipe10_io_pipe_phv_out_data_507; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_508 = pipe10_io_pipe_phv_out_data_508; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_509 = pipe10_io_pipe_phv_out_data_509; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_510 = pipe10_io_pipe_phv_out_data_510; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_511 = pipe10_io_pipe_phv_out_data_511; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_0 = pipe10_io_pipe_phv_out_header_0; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_1 = pipe10_io_pipe_phv_out_header_1; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_2 = pipe10_io_pipe_phv_out_header_2; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_3 = pipe10_io_pipe_phv_out_header_3; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_4 = pipe10_io_pipe_phv_out_header_4; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_5 = pipe10_io_pipe_phv_out_header_5; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_6 = pipe10_io_pipe_phv_out_header_6; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_7 = pipe10_io_pipe_phv_out_header_7; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_8 = pipe10_io_pipe_phv_out_header_8; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_9 = pipe10_io_pipe_phv_out_header_9; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_10 = pipe10_io_pipe_phv_out_header_10; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_11 = pipe10_io_pipe_phv_out_header_11; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_12 = pipe10_io_pipe_phv_out_header_12; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_13 = pipe10_io_pipe_phv_out_header_13; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_14 = pipe10_io_pipe_phv_out_header_14; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_15 = pipe10_io_pipe_phv_out_header_15; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_parse_current_state = pipe10_io_pipe_phv_out_parse_current_state; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_parse_current_offset = pipe10_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_parse_transition_field = pipe10_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_next_processor_id = pipe10_io_pipe_phv_out_next_processor_id; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_next_config_id = pipe10_io_pipe_phv_out_next_config_id; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_is_valid_processor = pipe10_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 377:27]
  assign pipe11_io_table_config_0_table_width = table_config_0_table_width; // @[matcher.scala 381:28]
  assign pipe11_io_table_config_0_table_depth = table_config_0_table_depth; // @[matcher.scala 381:28]
  assign pipe11_io_table_config_1_table_width = table_config_1_table_width; // @[matcher.scala 381:28]
  assign pipe11_io_table_config_1_table_depth = table_config_1_table_depth; // @[matcher.scala 381:28]
  assign pipe11_io_key_in = pipe10_io_key_out; // @[matcher.scala 378:27]
  assign pipe11_io_cs_in = pipe10_io_cs_out; // @[matcher.scala 379:27]
  assign pipe11_io_data_in_0 = pipe10_io_data_out_0; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_1 = pipe10_io_data_out_1; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_2 = pipe10_io_data_out_2; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_3 = pipe10_io_data_out_3; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_4 = pipe10_io_data_out_4; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_5 = pipe10_io_data_out_5; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_6 = pipe10_io_data_out_6; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_7 = pipe10_io_data_out_7; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_8 = pipe10_io_data_out_8; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_9 = pipe10_io_data_out_9; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_10 = pipe10_io_data_out_10; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_11 = pipe10_io_data_out_11; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_12 = pipe10_io_data_out_12; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_13 = pipe10_io_data_out_13; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_14 = pipe10_io_data_out_14; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_15 = pipe10_io_data_out_15; // @[matcher.scala 380:27]
  assign pipe12_clock = clock;
  assign pipe12_io_pipe_phv_in_data_0 = pipe11_io_pipe_phv_out_data_0; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_1 = pipe11_io_pipe_phv_out_data_1; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_2 = pipe11_io_pipe_phv_out_data_2; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_3 = pipe11_io_pipe_phv_out_data_3; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_4 = pipe11_io_pipe_phv_out_data_4; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_5 = pipe11_io_pipe_phv_out_data_5; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_6 = pipe11_io_pipe_phv_out_data_6; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_7 = pipe11_io_pipe_phv_out_data_7; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_8 = pipe11_io_pipe_phv_out_data_8; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_9 = pipe11_io_pipe_phv_out_data_9; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_10 = pipe11_io_pipe_phv_out_data_10; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_11 = pipe11_io_pipe_phv_out_data_11; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_12 = pipe11_io_pipe_phv_out_data_12; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_13 = pipe11_io_pipe_phv_out_data_13; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_14 = pipe11_io_pipe_phv_out_data_14; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_15 = pipe11_io_pipe_phv_out_data_15; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_16 = pipe11_io_pipe_phv_out_data_16; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_17 = pipe11_io_pipe_phv_out_data_17; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_18 = pipe11_io_pipe_phv_out_data_18; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_19 = pipe11_io_pipe_phv_out_data_19; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_20 = pipe11_io_pipe_phv_out_data_20; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_21 = pipe11_io_pipe_phv_out_data_21; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_22 = pipe11_io_pipe_phv_out_data_22; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_23 = pipe11_io_pipe_phv_out_data_23; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_24 = pipe11_io_pipe_phv_out_data_24; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_25 = pipe11_io_pipe_phv_out_data_25; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_26 = pipe11_io_pipe_phv_out_data_26; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_27 = pipe11_io_pipe_phv_out_data_27; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_28 = pipe11_io_pipe_phv_out_data_28; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_29 = pipe11_io_pipe_phv_out_data_29; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_30 = pipe11_io_pipe_phv_out_data_30; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_31 = pipe11_io_pipe_phv_out_data_31; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_32 = pipe11_io_pipe_phv_out_data_32; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_33 = pipe11_io_pipe_phv_out_data_33; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_34 = pipe11_io_pipe_phv_out_data_34; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_35 = pipe11_io_pipe_phv_out_data_35; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_36 = pipe11_io_pipe_phv_out_data_36; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_37 = pipe11_io_pipe_phv_out_data_37; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_38 = pipe11_io_pipe_phv_out_data_38; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_39 = pipe11_io_pipe_phv_out_data_39; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_40 = pipe11_io_pipe_phv_out_data_40; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_41 = pipe11_io_pipe_phv_out_data_41; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_42 = pipe11_io_pipe_phv_out_data_42; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_43 = pipe11_io_pipe_phv_out_data_43; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_44 = pipe11_io_pipe_phv_out_data_44; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_45 = pipe11_io_pipe_phv_out_data_45; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_46 = pipe11_io_pipe_phv_out_data_46; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_47 = pipe11_io_pipe_phv_out_data_47; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_48 = pipe11_io_pipe_phv_out_data_48; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_49 = pipe11_io_pipe_phv_out_data_49; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_50 = pipe11_io_pipe_phv_out_data_50; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_51 = pipe11_io_pipe_phv_out_data_51; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_52 = pipe11_io_pipe_phv_out_data_52; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_53 = pipe11_io_pipe_phv_out_data_53; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_54 = pipe11_io_pipe_phv_out_data_54; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_55 = pipe11_io_pipe_phv_out_data_55; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_56 = pipe11_io_pipe_phv_out_data_56; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_57 = pipe11_io_pipe_phv_out_data_57; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_58 = pipe11_io_pipe_phv_out_data_58; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_59 = pipe11_io_pipe_phv_out_data_59; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_60 = pipe11_io_pipe_phv_out_data_60; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_61 = pipe11_io_pipe_phv_out_data_61; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_62 = pipe11_io_pipe_phv_out_data_62; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_63 = pipe11_io_pipe_phv_out_data_63; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_64 = pipe11_io_pipe_phv_out_data_64; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_65 = pipe11_io_pipe_phv_out_data_65; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_66 = pipe11_io_pipe_phv_out_data_66; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_67 = pipe11_io_pipe_phv_out_data_67; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_68 = pipe11_io_pipe_phv_out_data_68; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_69 = pipe11_io_pipe_phv_out_data_69; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_70 = pipe11_io_pipe_phv_out_data_70; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_71 = pipe11_io_pipe_phv_out_data_71; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_72 = pipe11_io_pipe_phv_out_data_72; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_73 = pipe11_io_pipe_phv_out_data_73; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_74 = pipe11_io_pipe_phv_out_data_74; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_75 = pipe11_io_pipe_phv_out_data_75; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_76 = pipe11_io_pipe_phv_out_data_76; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_77 = pipe11_io_pipe_phv_out_data_77; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_78 = pipe11_io_pipe_phv_out_data_78; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_79 = pipe11_io_pipe_phv_out_data_79; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_80 = pipe11_io_pipe_phv_out_data_80; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_81 = pipe11_io_pipe_phv_out_data_81; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_82 = pipe11_io_pipe_phv_out_data_82; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_83 = pipe11_io_pipe_phv_out_data_83; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_84 = pipe11_io_pipe_phv_out_data_84; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_85 = pipe11_io_pipe_phv_out_data_85; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_86 = pipe11_io_pipe_phv_out_data_86; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_87 = pipe11_io_pipe_phv_out_data_87; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_88 = pipe11_io_pipe_phv_out_data_88; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_89 = pipe11_io_pipe_phv_out_data_89; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_90 = pipe11_io_pipe_phv_out_data_90; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_91 = pipe11_io_pipe_phv_out_data_91; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_92 = pipe11_io_pipe_phv_out_data_92; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_93 = pipe11_io_pipe_phv_out_data_93; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_94 = pipe11_io_pipe_phv_out_data_94; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_95 = pipe11_io_pipe_phv_out_data_95; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_96 = pipe11_io_pipe_phv_out_data_96; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_97 = pipe11_io_pipe_phv_out_data_97; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_98 = pipe11_io_pipe_phv_out_data_98; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_99 = pipe11_io_pipe_phv_out_data_99; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_100 = pipe11_io_pipe_phv_out_data_100; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_101 = pipe11_io_pipe_phv_out_data_101; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_102 = pipe11_io_pipe_phv_out_data_102; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_103 = pipe11_io_pipe_phv_out_data_103; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_104 = pipe11_io_pipe_phv_out_data_104; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_105 = pipe11_io_pipe_phv_out_data_105; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_106 = pipe11_io_pipe_phv_out_data_106; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_107 = pipe11_io_pipe_phv_out_data_107; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_108 = pipe11_io_pipe_phv_out_data_108; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_109 = pipe11_io_pipe_phv_out_data_109; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_110 = pipe11_io_pipe_phv_out_data_110; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_111 = pipe11_io_pipe_phv_out_data_111; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_112 = pipe11_io_pipe_phv_out_data_112; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_113 = pipe11_io_pipe_phv_out_data_113; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_114 = pipe11_io_pipe_phv_out_data_114; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_115 = pipe11_io_pipe_phv_out_data_115; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_116 = pipe11_io_pipe_phv_out_data_116; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_117 = pipe11_io_pipe_phv_out_data_117; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_118 = pipe11_io_pipe_phv_out_data_118; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_119 = pipe11_io_pipe_phv_out_data_119; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_120 = pipe11_io_pipe_phv_out_data_120; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_121 = pipe11_io_pipe_phv_out_data_121; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_122 = pipe11_io_pipe_phv_out_data_122; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_123 = pipe11_io_pipe_phv_out_data_123; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_124 = pipe11_io_pipe_phv_out_data_124; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_125 = pipe11_io_pipe_phv_out_data_125; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_126 = pipe11_io_pipe_phv_out_data_126; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_127 = pipe11_io_pipe_phv_out_data_127; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_128 = pipe11_io_pipe_phv_out_data_128; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_129 = pipe11_io_pipe_phv_out_data_129; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_130 = pipe11_io_pipe_phv_out_data_130; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_131 = pipe11_io_pipe_phv_out_data_131; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_132 = pipe11_io_pipe_phv_out_data_132; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_133 = pipe11_io_pipe_phv_out_data_133; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_134 = pipe11_io_pipe_phv_out_data_134; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_135 = pipe11_io_pipe_phv_out_data_135; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_136 = pipe11_io_pipe_phv_out_data_136; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_137 = pipe11_io_pipe_phv_out_data_137; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_138 = pipe11_io_pipe_phv_out_data_138; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_139 = pipe11_io_pipe_phv_out_data_139; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_140 = pipe11_io_pipe_phv_out_data_140; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_141 = pipe11_io_pipe_phv_out_data_141; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_142 = pipe11_io_pipe_phv_out_data_142; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_143 = pipe11_io_pipe_phv_out_data_143; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_144 = pipe11_io_pipe_phv_out_data_144; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_145 = pipe11_io_pipe_phv_out_data_145; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_146 = pipe11_io_pipe_phv_out_data_146; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_147 = pipe11_io_pipe_phv_out_data_147; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_148 = pipe11_io_pipe_phv_out_data_148; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_149 = pipe11_io_pipe_phv_out_data_149; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_150 = pipe11_io_pipe_phv_out_data_150; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_151 = pipe11_io_pipe_phv_out_data_151; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_152 = pipe11_io_pipe_phv_out_data_152; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_153 = pipe11_io_pipe_phv_out_data_153; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_154 = pipe11_io_pipe_phv_out_data_154; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_155 = pipe11_io_pipe_phv_out_data_155; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_156 = pipe11_io_pipe_phv_out_data_156; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_157 = pipe11_io_pipe_phv_out_data_157; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_158 = pipe11_io_pipe_phv_out_data_158; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_159 = pipe11_io_pipe_phv_out_data_159; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_160 = pipe11_io_pipe_phv_out_data_160; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_161 = pipe11_io_pipe_phv_out_data_161; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_162 = pipe11_io_pipe_phv_out_data_162; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_163 = pipe11_io_pipe_phv_out_data_163; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_164 = pipe11_io_pipe_phv_out_data_164; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_165 = pipe11_io_pipe_phv_out_data_165; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_166 = pipe11_io_pipe_phv_out_data_166; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_167 = pipe11_io_pipe_phv_out_data_167; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_168 = pipe11_io_pipe_phv_out_data_168; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_169 = pipe11_io_pipe_phv_out_data_169; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_170 = pipe11_io_pipe_phv_out_data_170; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_171 = pipe11_io_pipe_phv_out_data_171; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_172 = pipe11_io_pipe_phv_out_data_172; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_173 = pipe11_io_pipe_phv_out_data_173; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_174 = pipe11_io_pipe_phv_out_data_174; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_175 = pipe11_io_pipe_phv_out_data_175; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_176 = pipe11_io_pipe_phv_out_data_176; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_177 = pipe11_io_pipe_phv_out_data_177; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_178 = pipe11_io_pipe_phv_out_data_178; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_179 = pipe11_io_pipe_phv_out_data_179; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_180 = pipe11_io_pipe_phv_out_data_180; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_181 = pipe11_io_pipe_phv_out_data_181; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_182 = pipe11_io_pipe_phv_out_data_182; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_183 = pipe11_io_pipe_phv_out_data_183; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_184 = pipe11_io_pipe_phv_out_data_184; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_185 = pipe11_io_pipe_phv_out_data_185; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_186 = pipe11_io_pipe_phv_out_data_186; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_187 = pipe11_io_pipe_phv_out_data_187; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_188 = pipe11_io_pipe_phv_out_data_188; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_189 = pipe11_io_pipe_phv_out_data_189; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_190 = pipe11_io_pipe_phv_out_data_190; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_191 = pipe11_io_pipe_phv_out_data_191; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_192 = pipe11_io_pipe_phv_out_data_192; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_193 = pipe11_io_pipe_phv_out_data_193; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_194 = pipe11_io_pipe_phv_out_data_194; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_195 = pipe11_io_pipe_phv_out_data_195; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_196 = pipe11_io_pipe_phv_out_data_196; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_197 = pipe11_io_pipe_phv_out_data_197; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_198 = pipe11_io_pipe_phv_out_data_198; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_199 = pipe11_io_pipe_phv_out_data_199; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_200 = pipe11_io_pipe_phv_out_data_200; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_201 = pipe11_io_pipe_phv_out_data_201; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_202 = pipe11_io_pipe_phv_out_data_202; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_203 = pipe11_io_pipe_phv_out_data_203; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_204 = pipe11_io_pipe_phv_out_data_204; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_205 = pipe11_io_pipe_phv_out_data_205; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_206 = pipe11_io_pipe_phv_out_data_206; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_207 = pipe11_io_pipe_phv_out_data_207; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_208 = pipe11_io_pipe_phv_out_data_208; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_209 = pipe11_io_pipe_phv_out_data_209; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_210 = pipe11_io_pipe_phv_out_data_210; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_211 = pipe11_io_pipe_phv_out_data_211; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_212 = pipe11_io_pipe_phv_out_data_212; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_213 = pipe11_io_pipe_phv_out_data_213; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_214 = pipe11_io_pipe_phv_out_data_214; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_215 = pipe11_io_pipe_phv_out_data_215; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_216 = pipe11_io_pipe_phv_out_data_216; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_217 = pipe11_io_pipe_phv_out_data_217; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_218 = pipe11_io_pipe_phv_out_data_218; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_219 = pipe11_io_pipe_phv_out_data_219; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_220 = pipe11_io_pipe_phv_out_data_220; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_221 = pipe11_io_pipe_phv_out_data_221; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_222 = pipe11_io_pipe_phv_out_data_222; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_223 = pipe11_io_pipe_phv_out_data_223; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_224 = pipe11_io_pipe_phv_out_data_224; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_225 = pipe11_io_pipe_phv_out_data_225; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_226 = pipe11_io_pipe_phv_out_data_226; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_227 = pipe11_io_pipe_phv_out_data_227; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_228 = pipe11_io_pipe_phv_out_data_228; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_229 = pipe11_io_pipe_phv_out_data_229; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_230 = pipe11_io_pipe_phv_out_data_230; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_231 = pipe11_io_pipe_phv_out_data_231; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_232 = pipe11_io_pipe_phv_out_data_232; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_233 = pipe11_io_pipe_phv_out_data_233; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_234 = pipe11_io_pipe_phv_out_data_234; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_235 = pipe11_io_pipe_phv_out_data_235; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_236 = pipe11_io_pipe_phv_out_data_236; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_237 = pipe11_io_pipe_phv_out_data_237; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_238 = pipe11_io_pipe_phv_out_data_238; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_239 = pipe11_io_pipe_phv_out_data_239; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_240 = pipe11_io_pipe_phv_out_data_240; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_241 = pipe11_io_pipe_phv_out_data_241; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_242 = pipe11_io_pipe_phv_out_data_242; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_243 = pipe11_io_pipe_phv_out_data_243; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_244 = pipe11_io_pipe_phv_out_data_244; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_245 = pipe11_io_pipe_phv_out_data_245; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_246 = pipe11_io_pipe_phv_out_data_246; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_247 = pipe11_io_pipe_phv_out_data_247; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_248 = pipe11_io_pipe_phv_out_data_248; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_249 = pipe11_io_pipe_phv_out_data_249; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_250 = pipe11_io_pipe_phv_out_data_250; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_251 = pipe11_io_pipe_phv_out_data_251; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_252 = pipe11_io_pipe_phv_out_data_252; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_253 = pipe11_io_pipe_phv_out_data_253; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_254 = pipe11_io_pipe_phv_out_data_254; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_255 = pipe11_io_pipe_phv_out_data_255; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_256 = pipe11_io_pipe_phv_out_data_256; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_257 = pipe11_io_pipe_phv_out_data_257; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_258 = pipe11_io_pipe_phv_out_data_258; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_259 = pipe11_io_pipe_phv_out_data_259; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_260 = pipe11_io_pipe_phv_out_data_260; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_261 = pipe11_io_pipe_phv_out_data_261; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_262 = pipe11_io_pipe_phv_out_data_262; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_263 = pipe11_io_pipe_phv_out_data_263; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_264 = pipe11_io_pipe_phv_out_data_264; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_265 = pipe11_io_pipe_phv_out_data_265; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_266 = pipe11_io_pipe_phv_out_data_266; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_267 = pipe11_io_pipe_phv_out_data_267; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_268 = pipe11_io_pipe_phv_out_data_268; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_269 = pipe11_io_pipe_phv_out_data_269; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_270 = pipe11_io_pipe_phv_out_data_270; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_271 = pipe11_io_pipe_phv_out_data_271; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_272 = pipe11_io_pipe_phv_out_data_272; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_273 = pipe11_io_pipe_phv_out_data_273; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_274 = pipe11_io_pipe_phv_out_data_274; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_275 = pipe11_io_pipe_phv_out_data_275; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_276 = pipe11_io_pipe_phv_out_data_276; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_277 = pipe11_io_pipe_phv_out_data_277; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_278 = pipe11_io_pipe_phv_out_data_278; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_279 = pipe11_io_pipe_phv_out_data_279; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_280 = pipe11_io_pipe_phv_out_data_280; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_281 = pipe11_io_pipe_phv_out_data_281; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_282 = pipe11_io_pipe_phv_out_data_282; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_283 = pipe11_io_pipe_phv_out_data_283; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_284 = pipe11_io_pipe_phv_out_data_284; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_285 = pipe11_io_pipe_phv_out_data_285; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_286 = pipe11_io_pipe_phv_out_data_286; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_287 = pipe11_io_pipe_phv_out_data_287; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_288 = pipe11_io_pipe_phv_out_data_288; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_289 = pipe11_io_pipe_phv_out_data_289; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_290 = pipe11_io_pipe_phv_out_data_290; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_291 = pipe11_io_pipe_phv_out_data_291; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_292 = pipe11_io_pipe_phv_out_data_292; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_293 = pipe11_io_pipe_phv_out_data_293; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_294 = pipe11_io_pipe_phv_out_data_294; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_295 = pipe11_io_pipe_phv_out_data_295; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_296 = pipe11_io_pipe_phv_out_data_296; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_297 = pipe11_io_pipe_phv_out_data_297; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_298 = pipe11_io_pipe_phv_out_data_298; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_299 = pipe11_io_pipe_phv_out_data_299; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_300 = pipe11_io_pipe_phv_out_data_300; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_301 = pipe11_io_pipe_phv_out_data_301; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_302 = pipe11_io_pipe_phv_out_data_302; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_303 = pipe11_io_pipe_phv_out_data_303; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_304 = pipe11_io_pipe_phv_out_data_304; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_305 = pipe11_io_pipe_phv_out_data_305; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_306 = pipe11_io_pipe_phv_out_data_306; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_307 = pipe11_io_pipe_phv_out_data_307; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_308 = pipe11_io_pipe_phv_out_data_308; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_309 = pipe11_io_pipe_phv_out_data_309; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_310 = pipe11_io_pipe_phv_out_data_310; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_311 = pipe11_io_pipe_phv_out_data_311; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_312 = pipe11_io_pipe_phv_out_data_312; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_313 = pipe11_io_pipe_phv_out_data_313; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_314 = pipe11_io_pipe_phv_out_data_314; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_315 = pipe11_io_pipe_phv_out_data_315; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_316 = pipe11_io_pipe_phv_out_data_316; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_317 = pipe11_io_pipe_phv_out_data_317; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_318 = pipe11_io_pipe_phv_out_data_318; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_319 = pipe11_io_pipe_phv_out_data_319; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_320 = pipe11_io_pipe_phv_out_data_320; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_321 = pipe11_io_pipe_phv_out_data_321; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_322 = pipe11_io_pipe_phv_out_data_322; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_323 = pipe11_io_pipe_phv_out_data_323; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_324 = pipe11_io_pipe_phv_out_data_324; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_325 = pipe11_io_pipe_phv_out_data_325; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_326 = pipe11_io_pipe_phv_out_data_326; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_327 = pipe11_io_pipe_phv_out_data_327; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_328 = pipe11_io_pipe_phv_out_data_328; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_329 = pipe11_io_pipe_phv_out_data_329; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_330 = pipe11_io_pipe_phv_out_data_330; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_331 = pipe11_io_pipe_phv_out_data_331; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_332 = pipe11_io_pipe_phv_out_data_332; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_333 = pipe11_io_pipe_phv_out_data_333; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_334 = pipe11_io_pipe_phv_out_data_334; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_335 = pipe11_io_pipe_phv_out_data_335; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_336 = pipe11_io_pipe_phv_out_data_336; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_337 = pipe11_io_pipe_phv_out_data_337; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_338 = pipe11_io_pipe_phv_out_data_338; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_339 = pipe11_io_pipe_phv_out_data_339; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_340 = pipe11_io_pipe_phv_out_data_340; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_341 = pipe11_io_pipe_phv_out_data_341; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_342 = pipe11_io_pipe_phv_out_data_342; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_343 = pipe11_io_pipe_phv_out_data_343; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_344 = pipe11_io_pipe_phv_out_data_344; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_345 = pipe11_io_pipe_phv_out_data_345; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_346 = pipe11_io_pipe_phv_out_data_346; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_347 = pipe11_io_pipe_phv_out_data_347; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_348 = pipe11_io_pipe_phv_out_data_348; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_349 = pipe11_io_pipe_phv_out_data_349; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_350 = pipe11_io_pipe_phv_out_data_350; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_351 = pipe11_io_pipe_phv_out_data_351; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_352 = pipe11_io_pipe_phv_out_data_352; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_353 = pipe11_io_pipe_phv_out_data_353; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_354 = pipe11_io_pipe_phv_out_data_354; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_355 = pipe11_io_pipe_phv_out_data_355; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_356 = pipe11_io_pipe_phv_out_data_356; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_357 = pipe11_io_pipe_phv_out_data_357; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_358 = pipe11_io_pipe_phv_out_data_358; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_359 = pipe11_io_pipe_phv_out_data_359; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_360 = pipe11_io_pipe_phv_out_data_360; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_361 = pipe11_io_pipe_phv_out_data_361; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_362 = pipe11_io_pipe_phv_out_data_362; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_363 = pipe11_io_pipe_phv_out_data_363; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_364 = pipe11_io_pipe_phv_out_data_364; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_365 = pipe11_io_pipe_phv_out_data_365; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_366 = pipe11_io_pipe_phv_out_data_366; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_367 = pipe11_io_pipe_phv_out_data_367; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_368 = pipe11_io_pipe_phv_out_data_368; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_369 = pipe11_io_pipe_phv_out_data_369; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_370 = pipe11_io_pipe_phv_out_data_370; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_371 = pipe11_io_pipe_phv_out_data_371; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_372 = pipe11_io_pipe_phv_out_data_372; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_373 = pipe11_io_pipe_phv_out_data_373; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_374 = pipe11_io_pipe_phv_out_data_374; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_375 = pipe11_io_pipe_phv_out_data_375; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_376 = pipe11_io_pipe_phv_out_data_376; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_377 = pipe11_io_pipe_phv_out_data_377; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_378 = pipe11_io_pipe_phv_out_data_378; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_379 = pipe11_io_pipe_phv_out_data_379; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_380 = pipe11_io_pipe_phv_out_data_380; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_381 = pipe11_io_pipe_phv_out_data_381; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_382 = pipe11_io_pipe_phv_out_data_382; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_383 = pipe11_io_pipe_phv_out_data_383; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_384 = pipe11_io_pipe_phv_out_data_384; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_385 = pipe11_io_pipe_phv_out_data_385; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_386 = pipe11_io_pipe_phv_out_data_386; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_387 = pipe11_io_pipe_phv_out_data_387; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_388 = pipe11_io_pipe_phv_out_data_388; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_389 = pipe11_io_pipe_phv_out_data_389; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_390 = pipe11_io_pipe_phv_out_data_390; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_391 = pipe11_io_pipe_phv_out_data_391; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_392 = pipe11_io_pipe_phv_out_data_392; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_393 = pipe11_io_pipe_phv_out_data_393; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_394 = pipe11_io_pipe_phv_out_data_394; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_395 = pipe11_io_pipe_phv_out_data_395; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_396 = pipe11_io_pipe_phv_out_data_396; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_397 = pipe11_io_pipe_phv_out_data_397; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_398 = pipe11_io_pipe_phv_out_data_398; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_399 = pipe11_io_pipe_phv_out_data_399; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_400 = pipe11_io_pipe_phv_out_data_400; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_401 = pipe11_io_pipe_phv_out_data_401; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_402 = pipe11_io_pipe_phv_out_data_402; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_403 = pipe11_io_pipe_phv_out_data_403; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_404 = pipe11_io_pipe_phv_out_data_404; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_405 = pipe11_io_pipe_phv_out_data_405; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_406 = pipe11_io_pipe_phv_out_data_406; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_407 = pipe11_io_pipe_phv_out_data_407; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_408 = pipe11_io_pipe_phv_out_data_408; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_409 = pipe11_io_pipe_phv_out_data_409; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_410 = pipe11_io_pipe_phv_out_data_410; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_411 = pipe11_io_pipe_phv_out_data_411; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_412 = pipe11_io_pipe_phv_out_data_412; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_413 = pipe11_io_pipe_phv_out_data_413; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_414 = pipe11_io_pipe_phv_out_data_414; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_415 = pipe11_io_pipe_phv_out_data_415; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_416 = pipe11_io_pipe_phv_out_data_416; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_417 = pipe11_io_pipe_phv_out_data_417; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_418 = pipe11_io_pipe_phv_out_data_418; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_419 = pipe11_io_pipe_phv_out_data_419; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_420 = pipe11_io_pipe_phv_out_data_420; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_421 = pipe11_io_pipe_phv_out_data_421; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_422 = pipe11_io_pipe_phv_out_data_422; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_423 = pipe11_io_pipe_phv_out_data_423; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_424 = pipe11_io_pipe_phv_out_data_424; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_425 = pipe11_io_pipe_phv_out_data_425; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_426 = pipe11_io_pipe_phv_out_data_426; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_427 = pipe11_io_pipe_phv_out_data_427; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_428 = pipe11_io_pipe_phv_out_data_428; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_429 = pipe11_io_pipe_phv_out_data_429; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_430 = pipe11_io_pipe_phv_out_data_430; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_431 = pipe11_io_pipe_phv_out_data_431; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_432 = pipe11_io_pipe_phv_out_data_432; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_433 = pipe11_io_pipe_phv_out_data_433; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_434 = pipe11_io_pipe_phv_out_data_434; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_435 = pipe11_io_pipe_phv_out_data_435; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_436 = pipe11_io_pipe_phv_out_data_436; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_437 = pipe11_io_pipe_phv_out_data_437; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_438 = pipe11_io_pipe_phv_out_data_438; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_439 = pipe11_io_pipe_phv_out_data_439; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_440 = pipe11_io_pipe_phv_out_data_440; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_441 = pipe11_io_pipe_phv_out_data_441; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_442 = pipe11_io_pipe_phv_out_data_442; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_443 = pipe11_io_pipe_phv_out_data_443; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_444 = pipe11_io_pipe_phv_out_data_444; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_445 = pipe11_io_pipe_phv_out_data_445; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_446 = pipe11_io_pipe_phv_out_data_446; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_447 = pipe11_io_pipe_phv_out_data_447; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_448 = pipe11_io_pipe_phv_out_data_448; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_449 = pipe11_io_pipe_phv_out_data_449; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_450 = pipe11_io_pipe_phv_out_data_450; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_451 = pipe11_io_pipe_phv_out_data_451; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_452 = pipe11_io_pipe_phv_out_data_452; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_453 = pipe11_io_pipe_phv_out_data_453; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_454 = pipe11_io_pipe_phv_out_data_454; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_455 = pipe11_io_pipe_phv_out_data_455; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_456 = pipe11_io_pipe_phv_out_data_456; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_457 = pipe11_io_pipe_phv_out_data_457; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_458 = pipe11_io_pipe_phv_out_data_458; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_459 = pipe11_io_pipe_phv_out_data_459; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_460 = pipe11_io_pipe_phv_out_data_460; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_461 = pipe11_io_pipe_phv_out_data_461; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_462 = pipe11_io_pipe_phv_out_data_462; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_463 = pipe11_io_pipe_phv_out_data_463; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_464 = pipe11_io_pipe_phv_out_data_464; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_465 = pipe11_io_pipe_phv_out_data_465; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_466 = pipe11_io_pipe_phv_out_data_466; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_467 = pipe11_io_pipe_phv_out_data_467; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_468 = pipe11_io_pipe_phv_out_data_468; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_469 = pipe11_io_pipe_phv_out_data_469; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_470 = pipe11_io_pipe_phv_out_data_470; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_471 = pipe11_io_pipe_phv_out_data_471; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_472 = pipe11_io_pipe_phv_out_data_472; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_473 = pipe11_io_pipe_phv_out_data_473; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_474 = pipe11_io_pipe_phv_out_data_474; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_475 = pipe11_io_pipe_phv_out_data_475; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_476 = pipe11_io_pipe_phv_out_data_476; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_477 = pipe11_io_pipe_phv_out_data_477; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_478 = pipe11_io_pipe_phv_out_data_478; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_479 = pipe11_io_pipe_phv_out_data_479; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_480 = pipe11_io_pipe_phv_out_data_480; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_481 = pipe11_io_pipe_phv_out_data_481; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_482 = pipe11_io_pipe_phv_out_data_482; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_483 = pipe11_io_pipe_phv_out_data_483; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_484 = pipe11_io_pipe_phv_out_data_484; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_485 = pipe11_io_pipe_phv_out_data_485; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_486 = pipe11_io_pipe_phv_out_data_486; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_487 = pipe11_io_pipe_phv_out_data_487; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_488 = pipe11_io_pipe_phv_out_data_488; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_489 = pipe11_io_pipe_phv_out_data_489; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_490 = pipe11_io_pipe_phv_out_data_490; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_491 = pipe11_io_pipe_phv_out_data_491; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_492 = pipe11_io_pipe_phv_out_data_492; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_493 = pipe11_io_pipe_phv_out_data_493; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_494 = pipe11_io_pipe_phv_out_data_494; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_495 = pipe11_io_pipe_phv_out_data_495; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_496 = pipe11_io_pipe_phv_out_data_496; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_497 = pipe11_io_pipe_phv_out_data_497; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_498 = pipe11_io_pipe_phv_out_data_498; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_499 = pipe11_io_pipe_phv_out_data_499; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_500 = pipe11_io_pipe_phv_out_data_500; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_501 = pipe11_io_pipe_phv_out_data_501; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_502 = pipe11_io_pipe_phv_out_data_502; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_503 = pipe11_io_pipe_phv_out_data_503; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_504 = pipe11_io_pipe_phv_out_data_504; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_505 = pipe11_io_pipe_phv_out_data_505; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_506 = pipe11_io_pipe_phv_out_data_506; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_507 = pipe11_io_pipe_phv_out_data_507; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_508 = pipe11_io_pipe_phv_out_data_508; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_509 = pipe11_io_pipe_phv_out_data_509; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_510 = pipe11_io_pipe_phv_out_data_510; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_511 = pipe11_io_pipe_phv_out_data_511; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_0 = pipe11_io_pipe_phv_out_header_0; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_1 = pipe11_io_pipe_phv_out_header_1; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_2 = pipe11_io_pipe_phv_out_header_2; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_3 = pipe11_io_pipe_phv_out_header_3; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_4 = pipe11_io_pipe_phv_out_header_4; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_5 = pipe11_io_pipe_phv_out_header_5; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_6 = pipe11_io_pipe_phv_out_header_6; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_7 = pipe11_io_pipe_phv_out_header_7; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_8 = pipe11_io_pipe_phv_out_header_8; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_9 = pipe11_io_pipe_phv_out_header_9; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_10 = pipe11_io_pipe_phv_out_header_10; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_11 = pipe11_io_pipe_phv_out_header_11; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_12 = pipe11_io_pipe_phv_out_header_12; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_13 = pipe11_io_pipe_phv_out_header_13; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_14 = pipe11_io_pipe_phv_out_header_14; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_15 = pipe11_io_pipe_phv_out_header_15; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_parse_current_state = pipe11_io_pipe_phv_out_parse_current_state; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_parse_current_offset = pipe11_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_parse_transition_field = pipe11_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_next_processor_id = pipe11_io_pipe_phv_out_next_processor_id; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_next_config_id = pipe11_io_pipe_phv_out_next_config_id; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_is_valid_processor = pipe11_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 383:27]
  assign pipe12_io_key_config_0_key_length = key_config_0_key_length; // @[matcher.scala 386:27]
  assign pipe12_io_key_config_1_key_length = key_config_1_key_length; // @[matcher.scala 386:27]
  assign pipe12_io_key_in = pipe11_io_key_out; // @[matcher.scala 384:27]
  assign pipe12_io_data_in = pipe11_io_data_out; // @[matcher.scala 385:27]
  always @(posedge clock) begin
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_0_header_id <= io_mod_key_mod_header_id; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_0_internal_offset <= io_mod_key_mod_internal_offset; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_0_key_length <= io_mod_key_mod_key_length; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_1_header_id <= io_mod_key_mod_header_id; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_1_internal_offset <= io_mod_key_mod_internal_offset; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_1_key_length <= io_mod_key_mod_key_length; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_table_width <= io_mod_table_mod_table_width; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_table_depth <= io_mod_table_mod_table_depth; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_table_width <= io_mod_table_mod_table_width; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_table_depth <= io_mod_table_mod_table_depth; // @[matcher.scala 22:40]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  key_config_0_header_id = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  key_config_0_internal_offset = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  key_config_0_key_length = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  key_config_1_header_id = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  key_config_1_internal_offset = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  key_config_1_key_length = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  table_config_0_table_width = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  table_config_0_table_depth = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  table_config_1_table_width = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  table_config_1_table_depth = _RAND_9[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
